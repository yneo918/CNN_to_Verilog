module layer
	#(parameter WIDTH = 8)
	(x, z);
	localparam IN = 400;
	input [WIDTH-1:0] x[0:IN-1];
	output [WIDTH*2+$clog2(82)-1:0] z;
	wire [WIDTH*2-1+0:0] tmp00[0:81];
	wire [WIDTH*2-1+1:0] tmp01[0:40];
	wire [WIDTH*2-1+2:0] tmp02[0:20];
	wire [WIDTH*2-1+3:0] tmp03[0:10];
	wire [WIDTH*2-1+4:0] tmp04[0:5];
	wire [WIDTH*2-1+5:0] tmp05[0:2];
	wire [WIDTH*2-1+6:0] tmp06[0:1];
	wire [WIDTH*2-1+7:0] tmp07[0:0];
	booth__004 #(.WIDTH(WIDTH)) mul00(.x(x[2]), .z(tmp00[0]));
	booth__004 #(.WIDTH(WIDTH)) mul01(.x(x[4]), .z(tmp00[1]));
	booth_0002 #(.WIDTH(WIDTH)) mul02(.x(x[5]), .z(tmp00[2]));
	booth_0004 #(.WIDTH(WIDTH)) mul03(.x(x[10]), .z(tmp00[3]));
	booth__004 #(.WIDTH(WIDTH)) mul04(.x(x[25]), .z(tmp00[4]));
	booth__002 #(.WIDTH(WIDTH)) mul05(.x(x[26]), .z(tmp00[5]));
	booth_0004 #(.WIDTH(WIDTH)) mul06(.x(x[30]), .z(tmp00[6]));
	booth_0004 #(.WIDTH(WIDTH)) mul07(.x(x[32]), .z(tmp00[7]));
	booth__002 #(.WIDTH(WIDTH)) mul08(.x(x[40]), .z(tmp00[8]));
	booth__004 #(.WIDTH(WIDTH)) mul09(.x(x[41]), .z(tmp00[9]));
	booth__002 #(.WIDTH(WIDTH)) mul10(.x(x[46]), .z(tmp00[10]));
	booth__004 #(.WIDTH(WIDTH)) mul11(.x(x[47]), .z(tmp00[11]));
	booth_0002 #(.WIDTH(WIDTH)) mul12(.x(x[55]), .z(tmp00[12]));
	booth__004 #(.WIDTH(WIDTH)) mul13(.x(x[58]), .z(tmp00[13]));
	booth__002 #(.WIDTH(WIDTH)) mul14(.x(x[60]), .z(tmp00[14]));
	booth__004 #(.WIDTH(WIDTH)) mul15(.x(x[66]), .z(tmp00[15]));
	booth__004 #(.WIDTH(WIDTH)) mul16(.x(x[68]), .z(tmp00[16]));
	booth__006 #(.WIDTH(WIDTH)) mul17(.x(x[76]), .z(tmp00[17]));
	booth__004 #(.WIDTH(WIDTH)) mul18(.x(x[79]), .z(tmp00[18]));
	booth__004 #(.WIDTH(WIDTH)) mul19(.x(x[94]), .z(tmp00[19]));
	booth_0004 #(.WIDTH(WIDTH)) mul20(.x(x[110]), .z(tmp00[20]));
	booth__004 #(.WIDTH(WIDTH)) mul21(.x(x[113]), .z(tmp00[21]));
	booth__004 #(.WIDTH(WIDTH)) mul22(.x(x[124]), .z(tmp00[22]));
	booth_0004 #(.WIDTH(WIDTH)) mul23(.x(x[126]), .z(tmp00[23]));
	booth__004 #(.WIDTH(WIDTH)) mul24(.x(x[134]), .z(tmp00[24]));
	booth__004 #(.WIDTH(WIDTH)) mul25(.x(x[142]), .z(tmp00[25]));
	booth__002 #(.WIDTH(WIDTH)) mul26(.x(x[143]), .z(tmp00[26]));
	booth__004 #(.WIDTH(WIDTH)) mul27(.x(x[145]), .z(tmp00[27]));
	booth__002 #(.WIDTH(WIDTH)) mul28(.x(x[146]), .z(tmp00[28]));
	booth__004 #(.WIDTH(WIDTH)) mul29(.x(x[148]), .z(tmp00[29]));
	booth__004 #(.WIDTH(WIDTH)) mul30(.x(x[149]), .z(tmp00[30]));
	booth__004 #(.WIDTH(WIDTH)) mul31(.x(x[151]), .z(tmp00[31]));
	booth__006 #(.WIDTH(WIDTH)) mul32(.x(x[159]), .z(tmp00[32]));
	booth__004 #(.WIDTH(WIDTH)) mul33(.x(x[161]), .z(tmp00[33]));
	booth__004 #(.WIDTH(WIDTH)) mul34(.x(x[173]), .z(tmp00[34]));
	booth__008 #(.WIDTH(WIDTH)) mul35(.x(x[175]), .z(tmp00[35]));
	booth_0002 #(.WIDTH(WIDTH)) mul36(.x(x[177]), .z(tmp00[36]));
	booth__004 #(.WIDTH(WIDTH)) mul37(.x(x[181]), .z(tmp00[37]));
	booth_0004 #(.WIDTH(WIDTH)) mul38(.x(x[185]), .z(tmp00[38]));
	booth__002 #(.WIDTH(WIDTH)) mul39(.x(x[187]), .z(tmp00[39]));
	booth__004 #(.WIDTH(WIDTH)) mul40(.x(x[188]), .z(tmp00[40]));
	booth__004 #(.WIDTH(WIDTH)) mul41(.x(x[191]), .z(tmp00[41]));
	booth_0002 #(.WIDTH(WIDTH)) mul42(.x(x[192]), .z(tmp00[42]));
	booth_0002 #(.WIDTH(WIDTH)) mul43(.x(x[193]), .z(tmp00[43]));
	booth__002 #(.WIDTH(WIDTH)) mul44(.x(x[201]), .z(tmp00[44]));
	booth__004 #(.WIDTH(WIDTH)) mul45(.x(x[203]), .z(tmp00[45]));
	booth__004 #(.WIDTH(WIDTH)) mul46(.x(x[204]), .z(tmp00[46]));
	booth__004 #(.WIDTH(WIDTH)) mul47(.x(x[206]), .z(tmp00[47]));
	booth__004 #(.WIDTH(WIDTH)) mul48(.x(x[208]), .z(tmp00[48]));
	booth__004 #(.WIDTH(WIDTH)) mul49(.x(x[209]), .z(tmp00[49]));
	booth_0004 #(.WIDTH(WIDTH)) mul50(.x(x[211]), .z(tmp00[50]));
	booth__004 #(.WIDTH(WIDTH)) mul51(.x(x[220]), .z(tmp00[51]));
	booth_0004 #(.WIDTH(WIDTH)) mul52(.x(x[225]), .z(tmp00[52]));
	booth_0002 #(.WIDTH(WIDTH)) mul53(.x(x[226]), .z(tmp00[53]));
	booth__002 #(.WIDTH(WIDTH)) mul54(.x(x[242]), .z(tmp00[54]));
	booth__002 #(.WIDTH(WIDTH)) mul55(.x(x[243]), .z(tmp00[55]));
	booth__004 #(.WIDTH(WIDTH)) mul56(.x(x[250]), .z(tmp00[56]));
	booth__002 #(.WIDTH(WIDTH)) mul57(.x(x[252]), .z(tmp00[57]));
	booth__002 #(.WIDTH(WIDTH)) mul58(.x(x[258]), .z(tmp00[58]));
	booth__002 #(.WIDTH(WIDTH)) mul59(.x(x[264]), .z(tmp00[59]));
	booth__004 #(.WIDTH(WIDTH)) mul60(.x(x[266]), .z(tmp00[60]));
	booth__004 #(.WIDTH(WIDTH)) mul61(.x(x[267]), .z(tmp00[61]));
	booth_0004 #(.WIDTH(WIDTH)) mul62(.x(x[271]), .z(tmp00[62]));
	booth_0004 #(.WIDTH(WIDTH)) mul63(.x(x[274]), .z(tmp00[63]));
	booth__002 #(.WIDTH(WIDTH)) mul64(.x(x[290]), .z(tmp00[64]));
	booth_0002 #(.WIDTH(WIDTH)) mul65(.x(x[301]), .z(tmp00[65]));
	booth__004 #(.WIDTH(WIDTH)) mul66(.x(x[306]), .z(tmp00[66]));
	booth_0002 #(.WIDTH(WIDTH)) mul67(.x(x[310]), .z(tmp00[67]));
	booth__004 #(.WIDTH(WIDTH)) mul68(.x(x[312]), .z(tmp00[68]));
	booth_0004 #(.WIDTH(WIDTH)) mul69(.x(x[321]), .z(tmp00[69]));
	booth__004 #(.WIDTH(WIDTH)) mul70(.x(x[329]), .z(tmp00[70]));
	booth__004 #(.WIDTH(WIDTH)) mul71(.x(x[330]), .z(tmp00[71]));
	booth_0002 #(.WIDTH(WIDTH)) mul72(.x(x[332]), .z(tmp00[72]));
	booth_0002 #(.WIDTH(WIDTH)) mul73(.x(x[337]), .z(tmp00[73]));
	booth__004 #(.WIDTH(WIDTH)) mul74(.x(x[356]), .z(tmp00[74]));
	booth_0002 #(.WIDTH(WIDTH)) mul75(.x(x[377]), .z(tmp00[75]));
	booth__002 #(.WIDTH(WIDTH)) mul76(.x(x[378]), .z(tmp00[76]));
	booth__002 #(.WIDTH(WIDTH)) mul77(.x(x[384]), .z(tmp00[77]));
	booth__002 #(.WIDTH(WIDTH)) mul78(.x(x[386]), .z(tmp00[78]));
	booth__004 #(.WIDTH(WIDTH)) mul79(.x(x[387]), .z(tmp00[79]));
	booth__004 #(.WIDTH(WIDTH)) mul80(.x(x[389]), .z(tmp00[80]));
	booth__004 #(.WIDTH(WIDTH)) mul81(.x(x[398]), .z(tmp00[81]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000000(.in0(tmp00[0]), .in1(tmp00[1]), .out(tmp01[0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000001(.in0(tmp00[2]), .in1(tmp00[3]), .out(tmp01[1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000002(.in0(tmp00[4]), .in1(tmp00[5]), .out(tmp01[2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000003(.in0(tmp00[6]), .in1(tmp00[7]), .out(tmp01[3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000004(.in0(tmp00[8]), .in1(tmp00[9]), .out(tmp01[4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000005(.in0(tmp00[10]), .in1(tmp00[11]), .out(tmp01[5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000006(.in0(tmp00[12]), .in1(tmp00[13]), .out(tmp01[6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000007(.in0(tmp00[14]), .in1(tmp00[15]), .out(tmp01[7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000008(.in0(tmp00[16]), .in1(tmp00[17]), .out(tmp01[8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000009(.in0(tmp00[18]), .in1(tmp00[19]), .out(tmp01[9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000010(.in0(tmp00[20]), .in1(tmp00[21]), .out(tmp01[10]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000011(.in0(tmp00[22]), .in1(tmp00[23]), .out(tmp01[11]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000012(.in0(tmp00[24]), .in1(tmp00[25]), .out(tmp01[12]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000013(.in0(tmp00[26]), .in1(tmp00[27]), .out(tmp01[13]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000014(.in0(tmp00[28]), .in1(tmp00[29]), .out(tmp01[14]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000015(.in0(tmp00[30]), .in1(tmp00[31]), .out(tmp01[15]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000016(.in0(tmp00[32]), .in1(tmp00[33]), .out(tmp01[16]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000017(.in0(tmp00[34]), .in1(tmp00[35]), .out(tmp01[17]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000018(.in0(tmp00[36]), .in1(tmp00[37]), .out(tmp01[18]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000019(.in0(tmp00[38]), .in1(tmp00[39]), .out(tmp01[19]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000020(.in0(tmp00[40]), .in1(tmp00[41]), .out(tmp01[20]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000021(.in0(tmp00[42]), .in1(tmp00[43]), .out(tmp01[21]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000022(.in0(tmp00[44]), .in1(tmp00[45]), .out(tmp01[22]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000023(.in0(tmp00[46]), .in1(tmp00[47]), .out(tmp01[23]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000024(.in0(tmp00[48]), .in1(tmp00[49]), .out(tmp01[24]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000025(.in0(tmp00[50]), .in1(tmp00[51]), .out(tmp01[25]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000026(.in0(tmp00[52]), .in1(tmp00[53]), .out(tmp01[26]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000027(.in0(tmp00[54]), .in1(tmp00[55]), .out(tmp01[27]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000028(.in0(tmp00[56]), .in1(tmp00[57]), .out(tmp01[28]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000029(.in0(tmp00[58]), .in1(tmp00[59]), .out(tmp01[29]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000030(.in0(tmp00[60]), .in1(tmp00[61]), .out(tmp01[30]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000031(.in0(tmp00[62]), .in1(tmp00[63]), .out(tmp01[31]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000032(.in0(tmp00[64]), .in1(tmp00[65]), .out(tmp01[32]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000033(.in0(tmp00[66]), .in1(tmp00[67]), .out(tmp01[33]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000034(.in0(tmp00[68]), .in1(tmp00[69]), .out(tmp01[34]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000035(.in0(tmp00[70]), .in1(tmp00[71]), .out(tmp01[35]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000036(.in0(tmp00[72]), .in1(tmp00[73]), .out(tmp01[36]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000037(.in0(tmp00[74]), .in1(tmp00[75]), .out(tmp01[37]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000038(.in0(tmp00[76]), .in1(tmp00[77]), .out(tmp01[38]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000039(.in0(tmp00[78]), .in1(tmp00[79]), .out(tmp01[39]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000040(.in0(tmp00[80]), .in1(tmp00[81]), .out(tmp01[40]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000041(.in0(tmp01[0]), .in1(tmp01[1]), .out(tmp02[0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000042(.in0(tmp01[2]), .in1(tmp01[3]), .out(tmp02[1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000043(.in0(tmp01[4]), .in1(tmp01[5]), .out(tmp02[2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000044(.in0(tmp01[6]), .in1(tmp01[7]), .out(tmp02[3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000045(.in0(tmp01[8]), .in1(tmp01[9]), .out(tmp02[4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000046(.in0(tmp01[10]), .in1(tmp01[11]), .out(tmp02[5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000047(.in0(tmp01[12]), .in1(tmp01[13]), .out(tmp02[6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000048(.in0(tmp01[14]), .in1(tmp01[15]), .out(tmp02[7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000049(.in0(tmp01[16]), .in1(tmp01[17]), .out(tmp02[8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000050(.in0(tmp01[18]), .in1(tmp01[19]), .out(tmp02[9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000051(.in0(tmp01[20]), .in1(tmp01[21]), .out(tmp02[10]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000052(.in0(tmp01[22]), .in1(tmp01[23]), .out(tmp02[11]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000053(.in0(tmp01[24]), .in1(tmp01[25]), .out(tmp02[12]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000054(.in0(tmp01[26]), .in1(tmp01[27]), .out(tmp02[13]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000055(.in0(tmp01[28]), .in1(tmp01[29]), .out(tmp02[14]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000056(.in0(tmp01[30]), .in1(tmp01[31]), .out(tmp02[15]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000057(.in0(tmp01[32]), .in1(tmp01[33]), .out(tmp02[16]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000058(.in0(tmp01[34]), .in1(tmp01[35]), .out(tmp02[17]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000059(.in0(tmp01[36]), .in1(tmp01[37]), .out(tmp02[18]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000060(.in0(tmp01[38]), .in1(tmp01[39]), .out(tmp02[19]));
	assign tmp02[20] = $signed(tmp01[40]);
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000061(.in0(tmp02[0]), .in1(tmp02[1]), .out(tmp03[0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000062(.in0(tmp02[2]), .in1(tmp02[3]), .out(tmp03[1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000063(.in0(tmp02[4]), .in1(tmp02[5]), .out(tmp03[2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000064(.in0(tmp02[6]), .in1(tmp02[7]), .out(tmp03[3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000065(.in0(tmp02[8]), .in1(tmp02[9]), .out(tmp03[4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000066(.in0(tmp02[10]), .in1(tmp02[11]), .out(tmp03[5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000067(.in0(tmp02[12]), .in1(tmp02[13]), .out(tmp03[6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000068(.in0(tmp02[14]), .in1(tmp02[15]), .out(tmp03[7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000069(.in0(tmp02[16]), .in1(tmp02[17]), .out(tmp03[8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000070(.in0(tmp02[18]), .in1(tmp02[19]), .out(tmp03[9]));
	assign tmp03[10] = $signed(tmp02[20]);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000071(.in0(tmp03[0]), .in1(tmp03[1]), .out(tmp04[0]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000072(.in0(tmp03[2]), .in1(tmp03[3]), .out(tmp04[1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000073(.in0(tmp03[4]), .in1(tmp03[5]), .out(tmp04[2]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000074(.in0(tmp03[6]), .in1(tmp03[7]), .out(tmp04[3]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000075(.in0(tmp03[8]), .in1(tmp03[9]), .out(tmp04[4]));
	assign tmp04[5] = $signed(tmp03[10]);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000076(.in0(tmp04[0]), .in1(tmp04[1]), .out(tmp05[0]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000077(.in0(tmp04[2]), .in1(tmp04[3]), .out(tmp05[1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000078(.in0(tmp04[4]), .in1(tmp04[5]), .out(tmp05[2]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000079(.in0(tmp05[0]), .in1(tmp05[1]), .out(tmp06[0]));
	assign tmp06[1] = $signed(tmp05[2]);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000080(.in0(tmp06[0]), .in1(tmp06[1]), .out(tmp07[0]));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU(.a(tmp07[0]), .b(23'h0), .sel(tmp07[0][WIDTH*2+$clog2(IN)-1]), .out(z));
endmodule

