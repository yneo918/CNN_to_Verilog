module fc128_84
	#(parameter WIDTH = 8)
	(x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7, x_8, x_9, x_10, x_11, x_12, x_13, x_14, x_15, x_16, x_17, x_18, x_19, x_20, x_21, x_22, x_23, x_24, x_25, x_26, x_27, x_28, x_29, x_30, x_31, x_32, x_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, x_84, x_85, x_86, x_87, x_88, x_89, x_90, x_91, x_92, x_93, x_94, x_95, x_96, x_97, x_98, x_99, x_100, x_101, x_102, x_103, x_104, x_105, x_106, x_107, x_108, x_109, x_110, x_111, x_112, x_113, x_114, x_115, x_116, x_117, x_118, x_119, x_120, x_121, x_122, x_123, x_124, x_125, x_126, x_127, z_0, z_1, z_2, z_3, z_4, z_5, z_6, z_7, z_8, z_9, z_10, z_11, z_12, z_13, z_14, z_15, z_16, z_17, z_18, z_19, z_20, z_21, z_22, z_23, z_24, z_25, z_26, z_27, z_28, z_29, z_30, z_31, z_32, z_33, z_34, z_35, z_36, z_37, z_38, z_39, z_40, z_41, z_42, z_43, z_44, z_45, z_46, z_47, z_48, z_49, z_50, z_51, z_52, z_53, z_54, z_55, z_56, z_57, z_58, z_59, z_60, z_61, z_62, z_63, z_64, z_65, z_66, z_67, z_68, z_69, z_70, z_71, z_72, z_73, z_74, z_75, z_76, z_77, z_78, z_79, z_80, z_81, z_82, z_83 );
	localparam IN = 128, OUT = 84;
	input [WIDTH-1:0] x_0;
	input [WIDTH-1:0] x_1;
	input [WIDTH-1:0] x_2;
	input [WIDTH-1:0] x_3;
	input [WIDTH-1:0] x_4;
	input [WIDTH-1:0] x_5;
	input [WIDTH-1:0] x_6;
	input [WIDTH-1:0] x_7;
	input [WIDTH-1:0] x_8;
	input [WIDTH-1:0] x_9;
	input [WIDTH-1:0] x_10;
	input [WIDTH-1:0] x_11;
	input [WIDTH-1:0] x_12;
	input [WIDTH-1:0] x_13;
	input [WIDTH-1:0] x_14;
	input [WIDTH-1:0] x_15;
	input [WIDTH-1:0] x_16;
	input [WIDTH-1:0] x_17;
	input [WIDTH-1:0] x_18;
	input [WIDTH-1:0] x_19;
	input [WIDTH-1:0] x_20;
	input [WIDTH-1:0] x_21;
	input [WIDTH-1:0] x_22;
	input [WIDTH-1:0] x_23;
	input [WIDTH-1:0] x_24;
	input [WIDTH-1:0] x_25;
	input [WIDTH-1:0] x_26;
	input [WIDTH-1:0] x_27;
	input [WIDTH-1:0] x_28;
	input [WIDTH-1:0] x_29;
	input [WIDTH-1:0] x_30;
	input [WIDTH-1:0] x_31;
	input [WIDTH-1:0] x_32;
	input [WIDTH-1:0] x_33;
	input [WIDTH-1:0] x_34;
	input [WIDTH-1:0] x_35;
	input [WIDTH-1:0] x_36;
	input [WIDTH-1:0] x_37;
	input [WIDTH-1:0] x_38;
	input [WIDTH-1:0] x_39;
	input [WIDTH-1:0] x_40;
	input [WIDTH-1:0] x_41;
	input [WIDTH-1:0] x_42;
	input [WIDTH-1:0] x_43;
	input [WIDTH-1:0] x_44;
	input [WIDTH-1:0] x_45;
	input [WIDTH-1:0] x_46;
	input [WIDTH-1:0] x_47;
	input [WIDTH-1:0] x_48;
	input [WIDTH-1:0] x_49;
	input [WIDTH-1:0] x_50;
	input [WIDTH-1:0] x_51;
	input [WIDTH-1:0] x_52;
	input [WIDTH-1:0] x_53;
	input [WIDTH-1:0] x_54;
	input [WIDTH-1:0] x_55;
	input [WIDTH-1:0] x_56;
	input [WIDTH-1:0] x_57;
	input [WIDTH-1:0] x_58;
	input [WIDTH-1:0] x_59;
	input [WIDTH-1:0] x_60;
	input [WIDTH-1:0] x_61;
	input [WIDTH-1:0] x_62;
	input [WIDTH-1:0] x_63;
	input [WIDTH-1:0] x_64;
	input [WIDTH-1:0] x_65;
	input [WIDTH-1:0] x_66;
	input [WIDTH-1:0] x_67;
	input [WIDTH-1:0] x_68;
	input [WIDTH-1:0] x_69;
	input [WIDTH-1:0] x_70;
	input [WIDTH-1:0] x_71;
	input [WIDTH-1:0] x_72;
	input [WIDTH-1:0] x_73;
	input [WIDTH-1:0] x_74;
	input [WIDTH-1:0] x_75;
	input [WIDTH-1:0] x_76;
	input [WIDTH-1:0] x_77;
	input [WIDTH-1:0] x_78;
	input [WIDTH-1:0] x_79;
	input [WIDTH-1:0] x_80;
	input [WIDTH-1:0] x_81;
	input [WIDTH-1:0] x_82;
	input [WIDTH-1:0] x_83;
	input [WIDTH-1:0] x_84;
	input [WIDTH-1:0] x_85;
	input [WIDTH-1:0] x_86;
	input [WIDTH-1:0] x_87;
	input [WIDTH-1:0] x_88;
	input [WIDTH-1:0] x_89;
	input [WIDTH-1:0] x_90;
	input [WIDTH-1:0] x_91;
	input [WIDTH-1:0] x_92;
	input [WIDTH-1:0] x_93;
	input [WIDTH-1:0] x_94;
	input [WIDTH-1:0] x_95;
	input [WIDTH-1:0] x_96;
	input [WIDTH-1:0] x_97;
	input [WIDTH-1:0] x_98;
	input [WIDTH-1:0] x_99;
	input [WIDTH-1:0] x_100;
	input [WIDTH-1:0] x_101;
	input [WIDTH-1:0] x_102;
	input [WIDTH-1:0] x_103;
	input [WIDTH-1:0] x_104;
	input [WIDTH-1:0] x_105;
	input [WIDTH-1:0] x_106;
	input [WIDTH-1:0] x_107;
	input [WIDTH-1:0] x_108;
	input [WIDTH-1:0] x_109;
	input [WIDTH-1:0] x_110;
	input [WIDTH-1:0] x_111;
	input [WIDTH-1:0] x_112;
	input [WIDTH-1:0] x_113;
	input [WIDTH-1:0] x_114;
	input [WIDTH-1:0] x_115;
	input [WIDTH-1:0] x_116;
	input [WIDTH-1:0] x_117;
	input [WIDTH-1:0] x_118;
	input [WIDTH-1:0] x_119;
	input [WIDTH-1:0] x_120;
	input [WIDTH-1:0] x_121;
	input [WIDTH-1:0] x_122;
	input [WIDTH-1:0] x_123;
	input [WIDTH-1:0] x_124;
	input [WIDTH-1:0] x_125;
	input [WIDTH-1:0] x_126;
	input [WIDTH-1:0] x_127;
	output [WIDTH-1:0] z_0;
	output [WIDTH-1:0] z_1;
	output [WIDTH-1:0] z_2;
	output [WIDTH-1:0] z_3;
	output [WIDTH-1:0] z_4;
	output [WIDTH-1:0] z_5;
	output [WIDTH-1:0] z_6;
	output [WIDTH-1:0] z_7;
	output [WIDTH-1:0] z_8;
	output [WIDTH-1:0] z_9;
	output [WIDTH-1:0] z_10;
	output [WIDTH-1:0] z_11;
	output [WIDTH-1:0] z_12;
	output [WIDTH-1:0] z_13;
	output [WIDTH-1:0] z_14;
	output [WIDTH-1:0] z_15;
	output [WIDTH-1:0] z_16;
	output [WIDTH-1:0] z_17;
	output [WIDTH-1:0] z_18;
	output [WIDTH-1:0] z_19;
	output [WIDTH-1:0] z_20;
	output [WIDTH-1:0] z_21;
	output [WIDTH-1:0] z_22;
	output [WIDTH-1:0] z_23;
	output [WIDTH-1:0] z_24;
	output [WIDTH-1:0] z_25;
	output [WIDTH-1:0] z_26;
	output [WIDTH-1:0] z_27;
	output [WIDTH-1:0] z_28;
	output [WIDTH-1:0] z_29;
	output [WIDTH-1:0] z_30;
	output [WIDTH-1:0] z_31;
	output [WIDTH-1:0] z_32;
	output [WIDTH-1:0] z_33;
	output [WIDTH-1:0] z_34;
	output [WIDTH-1:0] z_35;
	output [WIDTH-1:0] z_36;
	output [WIDTH-1:0] z_37;
	output [WIDTH-1:0] z_38;
	output [WIDTH-1:0] z_39;
	output [WIDTH-1:0] z_40;
	output [WIDTH-1:0] z_41;
	output [WIDTH-1:0] z_42;
	output [WIDTH-1:0] z_43;
	output [WIDTH-1:0] z_44;
	output [WIDTH-1:0] z_45;
	output [WIDTH-1:0] z_46;
	output [WIDTH-1:0] z_47;
	output [WIDTH-1:0] z_48;
	output [WIDTH-1:0] z_49;
	output [WIDTH-1:0] z_50;
	output [WIDTH-1:0] z_51;
	output [WIDTH-1:0] z_52;
	output [WIDTH-1:0] z_53;
	output [WIDTH-1:0] z_54;
	output [WIDTH-1:0] z_55;
	output [WIDTH-1:0] z_56;
	output [WIDTH-1:0] z_57;
	output [WIDTH-1:0] z_58;
	output [WIDTH-1:0] z_59;
	output [WIDTH-1:0] z_60;
	output [WIDTH-1:0] z_61;
	output [WIDTH-1:0] z_62;
	output [WIDTH-1:0] z_63;
	output [WIDTH-1:0] z_64;
	output [WIDTH-1:0] z_65;
	output [WIDTH-1:0] z_66;
	output [WIDTH-1:0] z_67;
	output [WIDTH-1:0] z_68;
	output [WIDTH-1:0] z_69;
	output [WIDTH-1:0] z_70;
	output [WIDTH-1:0] z_71;
	output [WIDTH-1:0] z_72;
	output [WIDTH-1:0] z_73;
	output [WIDTH-1:0] z_74;
	output [WIDTH-1:0] z_75;
	output [WIDTH-1:0] z_76;
	output [WIDTH-1:0] z_77;
	output [WIDTH-1:0] z_78;
	output [WIDTH-1:0] z_79;
	output [WIDTH-1:0] z_80;
	output [WIDTH-1:0] z_81;
	output [WIDTH-1:0] z_82;
	output [WIDTH-1:0] z_83;
	wire [WIDTH*2-1+0:0] tmp00_0_0;
	wire [WIDTH*2-1+0:0] tmp00_0_1;
	wire [WIDTH*2-1+0:0] tmp00_0_2;
	wire [WIDTH*2-1+0:0] tmp00_0_3;
	wire [WIDTH*2-1+0:0] tmp00_0_4;
	wire [WIDTH*2-1+0:0] tmp00_0_5;
	wire [WIDTH*2-1+0:0] tmp00_0_6;
	wire [WIDTH*2-1+0:0] tmp00_0_7;
	wire [WIDTH*2-1+0:0] tmp00_0_8;
	wire [WIDTH*2-1+0:0] tmp00_0_9;
	wire [WIDTH*2-1+0:0] tmp00_0_10;
	wire [WIDTH*2-1+0:0] tmp00_0_11;
	wire [WIDTH*2-1+0:0] tmp00_0_12;
	wire [WIDTH*2-1+0:0] tmp00_0_13;
	wire [WIDTH*2-1+0:0] tmp00_0_14;
	wire [WIDTH*2-1+0:0] tmp00_0_15;
	wire [WIDTH*2-1+0:0] tmp00_0_16;
	wire [WIDTH*2-1+0:0] tmp00_0_17;
	wire [WIDTH*2-1+0:0] tmp00_0_18;
	wire [WIDTH*2-1+0:0] tmp00_0_19;
	wire [WIDTH*2-1+0:0] tmp00_0_20;
	wire [WIDTH*2-1+0:0] tmp00_0_21;
	wire [WIDTH*2-1+0:0] tmp00_0_22;
	wire [WIDTH*2-1+0:0] tmp00_0_23;
	wire [WIDTH*2-1+0:0] tmp00_0_24;
	wire [WIDTH*2-1+0:0] tmp00_0_25;
	wire [WIDTH*2-1+0:0] tmp00_0_26;
	wire [WIDTH*2-1+0:0] tmp00_0_27;
	wire [WIDTH*2-1+0:0] tmp00_0_28;
	wire [WIDTH*2-1+0:0] tmp00_0_29;
	wire [WIDTH*2-1+0:0] tmp00_0_30;
	wire [WIDTH*2-1+0:0] tmp00_0_31;
	wire [WIDTH*2-1+0:0] tmp00_0_32;
	wire [WIDTH*2-1+0:0] tmp00_0_33;
	wire [WIDTH*2-1+0:0] tmp00_0_34;
	wire [WIDTH*2-1+0:0] tmp00_0_35;
	wire [WIDTH*2-1+0:0] tmp00_0_36;
	wire [WIDTH*2-1+0:0] tmp00_0_37;
	wire [WIDTH*2-1+0:0] tmp00_0_38;
	wire [WIDTH*2-1+0:0] tmp00_0_39;
	wire [WIDTH*2-1+0:0] tmp00_0_40;
	wire [WIDTH*2-1+0:0] tmp00_0_41;
	wire [WIDTH*2-1+0:0] tmp00_0_42;
	wire [WIDTH*2-1+0:0] tmp00_0_43;
	wire [WIDTH*2-1+0:0] tmp00_0_44;
	wire [WIDTH*2-1+0:0] tmp00_0_45;
	wire [WIDTH*2-1+0:0] tmp00_0_46;
	wire [WIDTH*2-1+0:0] tmp00_0_47;
	wire [WIDTH*2-1+0:0] tmp00_0_48;
	wire [WIDTH*2-1+0:0] tmp00_0_49;
	wire [WIDTH*2-1+0:0] tmp00_0_50;
	wire [WIDTH*2-1+0:0] tmp00_0_51;
	wire [WIDTH*2-1+0:0] tmp00_0_52;
	wire [WIDTH*2-1+0:0] tmp00_0_53;
	wire [WIDTH*2-1+0:0] tmp00_0_54;
	wire [WIDTH*2-1+0:0] tmp00_0_55;
	wire [WIDTH*2-1+0:0] tmp00_0_56;
	wire [WIDTH*2-1+0:0] tmp00_0_57;
	wire [WIDTH*2-1+0:0] tmp00_0_58;
	wire [WIDTH*2-1+0:0] tmp00_0_59;
	wire [WIDTH*2-1+0:0] tmp00_0_60;
	wire [WIDTH*2-1+0:0] tmp00_0_61;
	wire [WIDTH*2-1+0:0] tmp00_0_62;
	wire [WIDTH*2-1+0:0] tmp00_0_63;
	wire [WIDTH*2-1+0:0] tmp00_0_64;
	wire [WIDTH*2-1+0:0] tmp00_0_65;
	wire [WIDTH*2-1+0:0] tmp00_0_66;
	wire [WIDTH*2-1+0:0] tmp00_0_67;
	wire [WIDTH*2-1+0:0] tmp00_0_68;
	wire [WIDTH*2-1+0:0] tmp00_0_69;
	wire [WIDTH*2-1+0:0] tmp00_0_70;
	wire [WIDTH*2-1+0:0] tmp00_0_71;
	wire [WIDTH*2-1+0:0] tmp00_0_72;
	wire [WIDTH*2-1+0:0] tmp00_0_73;
	wire [WIDTH*2-1+0:0] tmp00_0_74;
	wire [WIDTH*2-1+0:0] tmp00_0_75;
	wire [WIDTH*2-1+0:0] tmp00_0_76;
	wire [WIDTH*2-1+0:0] tmp00_0_77;
	wire [WIDTH*2-1+0:0] tmp00_0_78;
	wire [WIDTH*2-1+0:0] tmp00_0_79;
	wire [WIDTH*2-1+0:0] tmp00_0_80;
	wire [WIDTH*2-1+0:0] tmp00_0_81;
	wire [WIDTH*2-1+0:0] tmp00_0_82;
	wire [WIDTH*2-1+0:0] tmp00_0_83;
	wire [WIDTH*2-1+0:0] tmp00_1_0;
	wire [WIDTH*2-1+0:0] tmp00_1_1;
	wire [WIDTH*2-1+0:0] tmp00_1_2;
	wire [WIDTH*2-1+0:0] tmp00_1_3;
	wire [WIDTH*2-1+0:0] tmp00_1_4;
	wire [WIDTH*2-1+0:0] tmp00_1_5;
	wire [WIDTH*2-1+0:0] tmp00_1_6;
	wire [WIDTH*2-1+0:0] tmp00_1_7;
	wire [WIDTH*2-1+0:0] tmp00_1_8;
	wire [WIDTH*2-1+0:0] tmp00_1_9;
	wire [WIDTH*2-1+0:0] tmp00_1_10;
	wire [WIDTH*2-1+0:0] tmp00_1_11;
	wire [WIDTH*2-1+0:0] tmp00_1_12;
	wire [WIDTH*2-1+0:0] tmp00_1_13;
	wire [WIDTH*2-1+0:0] tmp00_1_14;
	wire [WIDTH*2-1+0:0] tmp00_1_15;
	wire [WIDTH*2-1+0:0] tmp00_1_16;
	wire [WIDTH*2-1+0:0] tmp00_1_17;
	wire [WIDTH*2-1+0:0] tmp00_1_18;
	wire [WIDTH*2-1+0:0] tmp00_1_19;
	wire [WIDTH*2-1+0:0] tmp00_1_20;
	wire [WIDTH*2-1+0:0] tmp00_1_21;
	wire [WIDTH*2-1+0:0] tmp00_1_22;
	wire [WIDTH*2-1+0:0] tmp00_1_23;
	wire [WIDTH*2-1+0:0] tmp00_1_24;
	wire [WIDTH*2-1+0:0] tmp00_1_25;
	wire [WIDTH*2-1+0:0] tmp00_1_26;
	wire [WIDTH*2-1+0:0] tmp00_1_27;
	wire [WIDTH*2-1+0:0] tmp00_1_28;
	wire [WIDTH*2-1+0:0] tmp00_1_29;
	wire [WIDTH*2-1+0:0] tmp00_1_30;
	wire [WIDTH*2-1+0:0] tmp00_1_31;
	wire [WIDTH*2-1+0:0] tmp00_1_32;
	wire [WIDTH*2-1+0:0] tmp00_1_33;
	wire [WIDTH*2-1+0:0] tmp00_1_34;
	wire [WIDTH*2-1+0:0] tmp00_1_35;
	wire [WIDTH*2-1+0:0] tmp00_1_36;
	wire [WIDTH*2-1+0:0] tmp00_1_37;
	wire [WIDTH*2-1+0:0] tmp00_1_38;
	wire [WIDTH*2-1+0:0] tmp00_1_39;
	wire [WIDTH*2-1+0:0] tmp00_1_40;
	wire [WIDTH*2-1+0:0] tmp00_1_41;
	wire [WIDTH*2-1+0:0] tmp00_1_42;
	wire [WIDTH*2-1+0:0] tmp00_1_43;
	wire [WIDTH*2-1+0:0] tmp00_1_44;
	wire [WIDTH*2-1+0:0] tmp00_1_45;
	wire [WIDTH*2-1+0:0] tmp00_1_46;
	wire [WIDTH*2-1+0:0] tmp00_1_47;
	wire [WIDTH*2-1+0:0] tmp00_1_48;
	wire [WIDTH*2-1+0:0] tmp00_1_49;
	wire [WIDTH*2-1+0:0] tmp00_1_50;
	wire [WIDTH*2-1+0:0] tmp00_1_51;
	wire [WIDTH*2-1+0:0] tmp00_1_52;
	wire [WIDTH*2-1+0:0] tmp00_1_53;
	wire [WIDTH*2-1+0:0] tmp00_1_54;
	wire [WIDTH*2-1+0:0] tmp00_1_55;
	wire [WIDTH*2-1+0:0] tmp00_1_56;
	wire [WIDTH*2-1+0:0] tmp00_1_57;
	wire [WIDTH*2-1+0:0] tmp00_1_58;
	wire [WIDTH*2-1+0:0] tmp00_1_59;
	wire [WIDTH*2-1+0:0] tmp00_1_60;
	wire [WIDTH*2-1+0:0] tmp00_1_61;
	wire [WIDTH*2-1+0:0] tmp00_1_62;
	wire [WIDTH*2-1+0:0] tmp00_1_63;
	wire [WIDTH*2-1+0:0] tmp00_1_64;
	wire [WIDTH*2-1+0:0] tmp00_1_65;
	wire [WIDTH*2-1+0:0] tmp00_1_66;
	wire [WIDTH*2-1+0:0] tmp00_1_67;
	wire [WIDTH*2-1+0:0] tmp00_1_68;
	wire [WIDTH*2-1+0:0] tmp00_1_69;
	wire [WIDTH*2-1+0:0] tmp00_1_70;
	wire [WIDTH*2-1+0:0] tmp00_1_71;
	wire [WIDTH*2-1+0:0] tmp00_1_72;
	wire [WIDTH*2-1+0:0] tmp00_1_73;
	wire [WIDTH*2-1+0:0] tmp00_1_74;
	wire [WIDTH*2-1+0:0] tmp00_1_75;
	wire [WIDTH*2-1+0:0] tmp00_1_76;
	wire [WIDTH*2-1+0:0] tmp00_1_77;
	wire [WIDTH*2-1+0:0] tmp00_1_78;
	wire [WIDTH*2-1+0:0] tmp00_1_79;
	wire [WIDTH*2-1+0:0] tmp00_1_80;
	wire [WIDTH*2-1+0:0] tmp00_1_81;
	wire [WIDTH*2-1+0:0] tmp00_1_82;
	wire [WIDTH*2-1+0:0] tmp00_1_83;
	wire [WIDTH*2-1+0:0] tmp00_2_0;
	wire [WIDTH*2-1+0:0] tmp00_2_1;
	wire [WIDTH*2-1+0:0] tmp00_2_2;
	wire [WIDTH*2-1+0:0] tmp00_2_3;
	wire [WIDTH*2-1+0:0] tmp00_2_4;
	wire [WIDTH*2-1+0:0] tmp00_2_5;
	wire [WIDTH*2-1+0:0] tmp00_2_6;
	wire [WIDTH*2-1+0:0] tmp00_2_7;
	wire [WIDTH*2-1+0:0] tmp00_2_8;
	wire [WIDTH*2-1+0:0] tmp00_2_9;
	wire [WIDTH*2-1+0:0] tmp00_2_10;
	wire [WIDTH*2-1+0:0] tmp00_2_11;
	wire [WIDTH*2-1+0:0] tmp00_2_12;
	wire [WIDTH*2-1+0:0] tmp00_2_13;
	wire [WIDTH*2-1+0:0] tmp00_2_14;
	wire [WIDTH*2-1+0:0] tmp00_2_15;
	wire [WIDTH*2-1+0:0] tmp00_2_16;
	wire [WIDTH*2-1+0:0] tmp00_2_17;
	wire [WIDTH*2-1+0:0] tmp00_2_18;
	wire [WIDTH*2-1+0:0] tmp00_2_19;
	wire [WIDTH*2-1+0:0] tmp00_2_20;
	wire [WIDTH*2-1+0:0] tmp00_2_21;
	wire [WIDTH*2-1+0:0] tmp00_2_22;
	wire [WIDTH*2-1+0:0] tmp00_2_23;
	wire [WIDTH*2-1+0:0] tmp00_2_24;
	wire [WIDTH*2-1+0:0] tmp00_2_25;
	wire [WIDTH*2-1+0:0] tmp00_2_26;
	wire [WIDTH*2-1+0:0] tmp00_2_27;
	wire [WIDTH*2-1+0:0] tmp00_2_28;
	wire [WIDTH*2-1+0:0] tmp00_2_29;
	wire [WIDTH*2-1+0:0] tmp00_2_30;
	wire [WIDTH*2-1+0:0] tmp00_2_31;
	wire [WIDTH*2-1+0:0] tmp00_2_32;
	wire [WIDTH*2-1+0:0] tmp00_2_33;
	wire [WIDTH*2-1+0:0] tmp00_2_34;
	wire [WIDTH*2-1+0:0] tmp00_2_35;
	wire [WIDTH*2-1+0:0] tmp00_2_36;
	wire [WIDTH*2-1+0:0] tmp00_2_37;
	wire [WIDTH*2-1+0:0] tmp00_2_38;
	wire [WIDTH*2-1+0:0] tmp00_2_39;
	wire [WIDTH*2-1+0:0] tmp00_2_40;
	wire [WIDTH*2-1+0:0] tmp00_2_41;
	wire [WIDTH*2-1+0:0] tmp00_2_42;
	wire [WIDTH*2-1+0:0] tmp00_2_43;
	wire [WIDTH*2-1+0:0] tmp00_2_44;
	wire [WIDTH*2-1+0:0] tmp00_2_45;
	wire [WIDTH*2-1+0:0] tmp00_2_46;
	wire [WIDTH*2-1+0:0] tmp00_2_47;
	wire [WIDTH*2-1+0:0] tmp00_2_48;
	wire [WIDTH*2-1+0:0] tmp00_2_49;
	wire [WIDTH*2-1+0:0] tmp00_2_50;
	wire [WIDTH*2-1+0:0] tmp00_2_51;
	wire [WIDTH*2-1+0:0] tmp00_2_52;
	wire [WIDTH*2-1+0:0] tmp00_2_53;
	wire [WIDTH*2-1+0:0] tmp00_2_54;
	wire [WIDTH*2-1+0:0] tmp00_2_55;
	wire [WIDTH*2-1+0:0] tmp00_2_56;
	wire [WIDTH*2-1+0:0] tmp00_2_57;
	wire [WIDTH*2-1+0:0] tmp00_2_58;
	wire [WIDTH*2-1+0:0] tmp00_2_59;
	wire [WIDTH*2-1+0:0] tmp00_2_60;
	wire [WIDTH*2-1+0:0] tmp00_2_61;
	wire [WIDTH*2-1+0:0] tmp00_2_62;
	wire [WIDTH*2-1+0:0] tmp00_2_63;
	wire [WIDTH*2-1+0:0] tmp00_2_64;
	wire [WIDTH*2-1+0:0] tmp00_2_65;
	wire [WIDTH*2-1+0:0] tmp00_2_66;
	wire [WIDTH*2-1+0:0] tmp00_2_67;
	wire [WIDTH*2-1+0:0] tmp00_2_68;
	wire [WIDTH*2-1+0:0] tmp00_2_69;
	wire [WIDTH*2-1+0:0] tmp00_2_70;
	wire [WIDTH*2-1+0:0] tmp00_2_71;
	wire [WIDTH*2-1+0:0] tmp00_2_72;
	wire [WIDTH*2-1+0:0] tmp00_2_73;
	wire [WIDTH*2-1+0:0] tmp00_2_74;
	wire [WIDTH*2-1+0:0] tmp00_2_75;
	wire [WIDTH*2-1+0:0] tmp00_2_76;
	wire [WIDTH*2-1+0:0] tmp00_2_77;
	wire [WIDTH*2-1+0:0] tmp00_2_78;
	wire [WIDTH*2-1+0:0] tmp00_2_79;
	wire [WIDTH*2-1+0:0] tmp00_2_80;
	wire [WIDTH*2-1+0:0] tmp00_2_81;
	wire [WIDTH*2-1+0:0] tmp00_2_82;
	wire [WIDTH*2-1+0:0] tmp00_2_83;
	wire [WIDTH*2-1+0:0] tmp00_3_0;
	wire [WIDTH*2-1+0:0] tmp00_3_1;
	wire [WIDTH*2-1+0:0] tmp00_3_2;
	wire [WIDTH*2-1+0:0] tmp00_3_3;
	wire [WIDTH*2-1+0:0] tmp00_3_4;
	wire [WIDTH*2-1+0:0] tmp00_3_5;
	wire [WIDTH*2-1+0:0] tmp00_3_6;
	wire [WIDTH*2-1+0:0] tmp00_3_7;
	wire [WIDTH*2-1+0:0] tmp00_3_8;
	wire [WIDTH*2-1+0:0] tmp00_3_9;
	wire [WIDTH*2-1+0:0] tmp00_3_10;
	wire [WIDTH*2-1+0:0] tmp00_3_11;
	wire [WIDTH*2-1+0:0] tmp00_3_12;
	wire [WIDTH*2-1+0:0] tmp00_3_13;
	wire [WIDTH*2-1+0:0] tmp00_3_14;
	wire [WIDTH*2-1+0:0] tmp00_3_15;
	wire [WIDTH*2-1+0:0] tmp00_3_16;
	wire [WIDTH*2-1+0:0] tmp00_3_17;
	wire [WIDTH*2-1+0:0] tmp00_3_18;
	wire [WIDTH*2-1+0:0] tmp00_3_19;
	wire [WIDTH*2-1+0:0] tmp00_3_20;
	wire [WIDTH*2-1+0:0] tmp00_3_21;
	wire [WIDTH*2-1+0:0] tmp00_3_22;
	wire [WIDTH*2-1+0:0] tmp00_3_23;
	wire [WIDTH*2-1+0:0] tmp00_3_24;
	wire [WIDTH*2-1+0:0] tmp00_3_25;
	wire [WIDTH*2-1+0:0] tmp00_3_26;
	wire [WIDTH*2-1+0:0] tmp00_3_27;
	wire [WIDTH*2-1+0:0] tmp00_3_28;
	wire [WIDTH*2-1+0:0] tmp00_3_29;
	wire [WIDTH*2-1+0:0] tmp00_3_30;
	wire [WIDTH*2-1+0:0] tmp00_3_31;
	wire [WIDTH*2-1+0:0] tmp00_3_32;
	wire [WIDTH*2-1+0:0] tmp00_3_33;
	wire [WIDTH*2-1+0:0] tmp00_3_34;
	wire [WIDTH*2-1+0:0] tmp00_3_35;
	wire [WIDTH*2-1+0:0] tmp00_3_36;
	wire [WIDTH*2-1+0:0] tmp00_3_37;
	wire [WIDTH*2-1+0:0] tmp00_3_38;
	wire [WIDTH*2-1+0:0] tmp00_3_39;
	wire [WIDTH*2-1+0:0] tmp00_3_40;
	wire [WIDTH*2-1+0:0] tmp00_3_41;
	wire [WIDTH*2-1+0:0] tmp00_3_42;
	wire [WIDTH*2-1+0:0] tmp00_3_43;
	wire [WIDTH*2-1+0:0] tmp00_3_44;
	wire [WIDTH*2-1+0:0] tmp00_3_45;
	wire [WIDTH*2-1+0:0] tmp00_3_46;
	wire [WIDTH*2-1+0:0] tmp00_3_47;
	wire [WIDTH*2-1+0:0] tmp00_3_48;
	wire [WIDTH*2-1+0:0] tmp00_3_49;
	wire [WIDTH*2-1+0:0] tmp00_3_50;
	wire [WIDTH*2-1+0:0] tmp00_3_51;
	wire [WIDTH*2-1+0:0] tmp00_3_52;
	wire [WIDTH*2-1+0:0] tmp00_3_53;
	wire [WIDTH*2-1+0:0] tmp00_3_54;
	wire [WIDTH*2-1+0:0] tmp00_3_55;
	wire [WIDTH*2-1+0:0] tmp00_3_56;
	wire [WIDTH*2-1+0:0] tmp00_3_57;
	wire [WIDTH*2-1+0:0] tmp00_3_58;
	wire [WIDTH*2-1+0:0] tmp00_3_59;
	wire [WIDTH*2-1+0:0] tmp00_3_60;
	wire [WIDTH*2-1+0:0] tmp00_3_61;
	wire [WIDTH*2-1+0:0] tmp00_3_62;
	wire [WIDTH*2-1+0:0] tmp00_3_63;
	wire [WIDTH*2-1+0:0] tmp00_3_64;
	wire [WIDTH*2-1+0:0] tmp00_3_65;
	wire [WIDTH*2-1+0:0] tmp00_3_66;
	wire [WIDTH*2-1+0:0] tmp00_3_67;
	wire [WIDTH*2-1+0:0] tmp00_3_68;
	wire [WIDTH*2-1+0:0] tmp00_3_69;
	wire [WIDTH*2-1+0:0] tmp00_3_70;
	wire [WIDTH*2-1+0:0] tmp00_3_71;
	wire [WIDTH*2-1+0:0] tmp00_3_72;
	wire [WIDTH*2-1+0:0] tmp00_3_73;
	wire [WIDTH*2-1+0:0] tmp00_3_74;
	wire [WIDTH*2-1+0:0] tmp00_3_75;
	wire [WIDTH*2-1+0:0] tmp00_3_76;
	wire [WIDTH*2-1+0:0] tmp00_3_77;
	wire [WIDTH*2-1+0:0] tmp00_3_78;
	wire [WIDTH*2-1+0:0] tmp00_3_79;
	wire [WIDTH*2-1+0:0] tmp00_3_80;
	wire [WIDTH*2-1+0:0] tmp00_3_81;
	wire [WIDTH*2-1+0:0] tmp00_3_82;
	wire [WIDTH*2-1+0:0] tmp00_3_83;
	wire [WIDTH*2-1+0:0] tmp00_4_0;
	wire [WIDTH*2-1+0:0] tmp00_4_1;
	wire [WIDTH*2-1+0:0] tmp00_4_2;
	wire [WIDTH*2-1+0:0] tmp00_4_3;
	wire [WIDTH*2-1+0:0] tmp00_4_4;
	wire [WIDTH*2-1+0:0] tmp00_4_5;
	wire [WIDTH*2-1+0:0] tmp00_4_6;
	wire [WIDTH*2-1+0:0] tmp00_4_7;
	wire [WIDTH*2-1+0:0] tmp00_4_8;
	wire [WIDTH*2-1+0:0] tmp00_4_9;
	wire [WIDTH*2-1+0:0] tmp00_4_10;
	wire [WIDTH*2-1+0:0] tmp00_4_11;
	wire [WIDTH*2-1+0:0] tmp00_4_12;
	wire [WIDTH*2-1+0:0] tmp00_4_13;
	wire [WIDTH*2-1+0:0] tmp00_4_14;
	wire [WIDTH*2-1+0:0] tmp00_4_15;
	wire [WIDTH*2-1+0:0] tmp00_4_16;
	wire [WIDTH*2-1+0:0] tmp00_4_17;
	wire [WIDTH*2-1+0:0] tmp00_4_18;
	wire [WIDTH*2-1+0:0] tmp00_4_19;
	wire [WIDTH*2-1+0:0] tmp00_4_20;
	wire [WIDTH*2-1+0:0] tmp00_4_21;
	wire [WIDTH*2-1+0:0] tmp00_4_22;
	wire [WIDTH*2-1+0:0] tmp00_4_23;
	wire [WIDTH*2-1+0:0] tmp00_4_24;
	wire [WIDTH*2-1+0:0] tmp00_4_25;
	wire [WIDTH*2-1+0:0] tmp00_4_26;
	wire [WIDTH*2-1+0:0] tmp00_4_27;
	wire [WIDTH*2-1+0:0] tmp00_4_28;
	wire [WIDTH*2-1+0:0] tmp00_4_29;
	wire [WIDTH*2-1+0:0] tmp00_4_30;
	wire [WIDTH*2-1+0:0] tmp00_4_31;
	wire [WIDTH*2-1+0:0] tmp00_4_32;
	wire [WIDTH*2-1+0:0] tmp00_4_33;
	wire [WIDTH*2-1+0:0] tmp00_4_34;
	wire [WIDTH*2-1+0:0] tmp00_4_35;
	wire [WIDTH*2-1+0:0] tmp00_4_36;
	wire [WIDTH*2-1+0:0] tmp00_4_37;
	wire [WIDTH*2-1+0:0] tmp00_4_38;
	wire [WIDTH*2-1+0:0] tmp00_4_39;
	wire [WIDTH*2-1+0:0] tmp00_4_40;
	wire [WIDTH*2-1+0:0] tmp00_4_41;
	wire [WIDTH*2-1+0:0] tmp00_4_42;
	wire [WIDTH*2-1+0:0] tmp00_4_43;
	wire [WIDTH*2-1+0:0] tmp00_4_44;
	wire [WIDTH*2-1+0:0] tmp00_4_45;
	wire [WIDTH*2-1+0:0] tmp00_4_46;
	wire [WIDTH*2-1+0:0] tmp00_4_47;
	wire [WIDTH*2-1+0:0] tmp00_4_48;
	wire [WIDTH*2-1+0:0] tmp00_4_49;
	wire [WIDTH*2-1+0:0] tmp00_4_50;
	wire [WIDTH*2-1+0:0] tmp00_4_51;
	wire [WIDTH*2-1+0:0] tmp00_4_52;
	wire [WIDTH*2-1+0:0] tmp00_4_53;
	wire [WIDTH*2-1+0:0] tmp00_4_54;
	wire [WIDTH*2-1+0:0] tmp00_4_55;
	wire [WIDTH*2-1+0:0] tmp00_4_56;
	wire [WIDTH*2-1+0:0] tmp00_4_57;
	wire [WIDTH*2-1+0:0] tmp00_4_58;
	wire [WIDTH*2-1+0:0] tmp00_4_59;
	wire [WIDTH*2-1+0:0] tmp00_4_60;
	wire [WIDTH*2-1+0:0] tmp00_4_61;
	wire [WIDTH*2-1+0:0] tmp00_4_62;
	wire [WIDTH*2-1+0:0] tmp00_4_63;
	wire [WIDTH*2-1+0:0] tmp00_4_64;
	wire [WIDTH*2-1+0:0] tmp00_4_65;
	wire [WIDTH*2-1+0:0] tmp00_4_66;
	wire [WIDTH*2-1+0:0] tmp00_4_67;
	wire [WIDTH*2-1+0:0] tmp00_4_68;
	wire [WIDTH*2-1+0:0] tmp00_4_69;
	wire [WIDTH*2-1+0:0] tmp00_4_70;
	wire [WIDTH*2-1+0:0] tmp00_4_71;
	wire [WIDTH*2-1+0:0] tmp00_4_72;
	wire [WIDTH*2-1+0:0] tmp00_4_73;
	wire [WIDTH*2-1+0:0] tmp00_4_74;
	wire [WIDTH*2-1+0:0] tmp00_4_75;
	wire [WIDTH*2-1+0:0] tmp00_4_76;
	wire [WIDTH*2-1+0:0] tmp00_4_77;
	wire [WIDTH*2-1+0:0] tmp00_4_78;
	wire [WIDTH*2-1+0:0] tmp00_4_79;
	wire [WIDTH*2-1+0:0] tmp00_4_80;
	wire [WIDTH*2-1+0:0] tmp00_4_81;
	wire [WIDTH*2-1+0:0] tmp00_4_82;
	wire [WIDTH*2-1+0:0] tmp00_4_83;
	wire [WIDTH*2-1+0:0] tmp00_5_0;
	wire [WIDTH*2-1+0:0] tmp00_5_1;
	wire [WIDTH*2-1+0:0] tmp00_5_2;
	wire [WIDTH*2-1+0:0] tmp00_5_3;
	wire [WIDTH*2-1+0:0] tmp00_5_4;
	wire [WIDTH*2-1+0:0] tmp00_5_5;
	wire [WIDTH*2-1+0:0] tmp00_5_6;
	wire [WIDTH*2-1+0:0] tmp00_5_7;
	wire [WIDTH*2-1+0:0] tmp00_5_8;
	wire [WIDTH*2-1+0:0] tmp00_5_9;
	wire [WIDTH*2-1+0:0] tmp00_5_10;
	wire [WIDTH*2-1+0:0] tmp00_5_11;
	wire [WIDTH*2-1+0:0] tmp00_5_12;
	wire [WIDTH*2-1+0:0] tmp00_5_13;
	wire [WIDTH*2-1+0:0] tmp00_5_14;
	wire [WIDTH*2-1+0:0] tmp00_5_15;
	wire [WIDTH*2-1+0:0] tmp00_5_16;
	wire [WIDTH*2-1+0:0] tmp00_5_17;
	wire [WIDTH*2-1+0:0] tmp00_5_18;
	wire [WIDTH*2-1+0:0] tmp00_5_19;
	wire [WIDTH*2-1+0:0] tmp00_5_20;
	wire [WIDTH*2-1+0:0] tmp00_5_21;
	wire [WIDTH*2-1+0:0] tmp00_5_22;
	wire [WIDTH*2-1+0:0] tmp00_5_23;
	wire [WIDTH*2-1+0:0] tmp00_5_24;
	wire [WIDTH*2-1+0:0] tmp00_5_25;
	wire [WIDTH*2-1+0:0] tmp00_5_26;
	wire [WIDTH*2-1+0:0] tmp00_5_27;
	wire [WIDTH*2-1+0:0] tmp00_5_28;
	wire [WIDTH*2-1+0:0] tmp00_5_29;
	wire [WIDTH*2-1+0:0] tmp00_5_30;
	wire [WIDTH*2-1+0:0] tmp00_5_31;
	wire [WIDTH*2-1+0:0] tmp00_5_32;
	wire [WIDTH*2-1+0:0] tmp00_5_33;
	wire [WIDTH*2-1+0:0] tmp00_5_34;
	wire [WIDTH*2-1+0:0] tmp00_5_35;
	wire [WIDTH*2-1+0:0] tmp00_5_36;
	wire [WIDTH*2-1+0:0] tmp00_5_37;
	wire [WIDTH*2-1+0:0] tmp00_5_38;
	wire [WIDTH*2-1+0:0] tmp00_5_39;
	wire [WIDTH*2-1+0:0] tmp00_5_40;
	wire [WIDTH*2-1+0:0] tmp00_5_41;
	wire [WIDTH*2-1+0:0] tmp00_5_42;
	wire [WIDTH*2-1+0:0] tmp00_5_43;
	wire [WIDTH*2-1+0:0] tmp00_5_44;
	wire [WIDTH*2-1+0:0] tmp00_5_45;
	wire [WIDTH*2-1+0:0] tmp00_5_46;
	wire [WIDTH*2-1+0:0] tmp00_5_47;
	wire [WIDTH*2-1+0:0] tmp00_5_48;
	wire [WIDTH*2-1+0:0] tmp00_5_49;
	wire [WIDTH*2-1+0:0] tmp00_5_50;
	wire [WIDTH*2-1+0:0] tmp00_5_51;
	wire [WIDTH*2-1+0:0] tmp00_5_52;
	wire [WIDTH*2-1+0:0] tmp00_5_53;
	wire [WIDTH*2-1+0:0] tmp00_5_54;
	wire [WIDTH*2-1+0:0] tmp00_5_55;
	wire [WIDTH*2-1+0:0] tmp00_5_56;
	wire [WIDTH*2-1+0:0] tmp00_5_57;
	wire [WIDTH*2-1+0:0] tmp00_5_58;
	wire [WIDTH*2-1+0:0] tmp00_5_59;
	wire [WIDTH*2-1+0:0] tmp00_5_60;
	wire [WIDTH*2-1+0:0] tmp00_5_61;
	wire [WIDTH*2-1+0:0] tmp00_5_62;
	wire [WIDTH*2-1+0:0] tmp00_5_63;
	wire [WIDTH*2-1+0:0] tmp00_5_64;
	wire [WIDTH*2-1+0:0] tmp00_5_65;
	wire [WIDTH*2-1+0:0] tmp00_5_66;
	wire [WIDTH*2-1+0:0] tmp00_5_67;
	wire [WIDTH*2-1+0:0] tmp00_5_68;
	wire [WIDTH*2-1+0:0] tmp00_5_69;
	wire [WIDTH*2-1+0:0] tmp00_5_70;
	wire [WIDTH*2-1+0:0] tmp00_5_71;
	wire [WIDTH*2-1+0:0] tmp00_5_72;
	wire [WIDTH*2-1+0:0] tmp00_5_73;
	wire [WIDTH*2-1+0:0] tmp00_5_74;
	wire [WIDTH*2-1+0:0] tmp00_5_75;
	wire [WIDTH*2-1+0:0] tmp00_5_76;
	wire [WIDTH*2-1+0:0] tmp00_5_77;
	wire [WIDTH*2-1+0:0] tmp00_5_78;
	wire [WIDTH*2-1+0:0] tmp00_5_79;
	wire [WIDTH*2-1+0:0] tmp00_5_80;
	wire [WIDTH*2-1+0:0] tmp00_5_81;
	wire [WIDTH*2-1+0:0] tmp00_5_82;
	wire [WIDTH*2-1+0:0] tmp00_5_83;
	wire [WIDTH*2-1+0:0] tmp00_6_0;
	wire [WIDTH*2-1+0:0] tmp00_6_1;
	wire [WIDTH*2-1+0:0] tmp00_6_2;
	wire [WIDTH*2-1+0:0] tmp00_6_3;
	wire [WIDTH*2-1+0:0] tmp00_6_4;
	wire [WIDTH*2-1+0:0] tmp00_6_5;
	wire [WIDTH*2-1+0:0] tmp00_6_6;
	wire [WIDTH*2-1+0:0] tmp00_6_7;
	wire [WIDTH*2-1+0:0] tmp00_6_8;
	wire [WIDTH*2-1+0:0] tmp00_6_9;
	wire [WIDTH*2-1+0:0] tmp00_6_10;
	wire [WIDTH*2-1+0:0] tmp00_6_11;
	wire [WIDTH*2-1+0:0] tmp00_6_12;
	wire [WIDTH*2-1+0:0] tmp00_6_13;
	wire [WIDTH*2-1+0:0] tmp00_6_14;
	wire [WIDTH*2-1+0:0] tmp00_6_15;
	wire [WIDTH*2-1+0:0] tmp00_6_16;
	wire [WIDTH*2-1+0:0] tmp00_6_17;
	wire [WIDTH*2-1+0:0] tmp00_6_18;
	wire [WIDTH*2-1+0:0] tmp00_6_19;
	wire [WIDTH*2-1+0:0] tmp00_6_20;
	wire [WIDTH*2-1+0:0] tmp00_6_21;
	wire [WIDTH*2-1+0:0] tmp00_6_22;
	wire [WIDTH*2-1+0:0] tmp00_6_23;
	wire [WIDTH*2-1+0:0] tmp00_6_24;
	wire [WIDTH*2-1+0:0] tmp00_6_25;
	wire [WIDTH*2-1+0:0] tmp00_6_26;
	wire [WIDTH*2-1+0:0] tmp00_6_27;
	wire [WIDTH*2-1+0:0] tmp00_6_28;
	wire [WIDTH*2-1+0:0] tmp00_6_29;
	wire [WIDTH*2-1+0:0] tmp00_6_30;
	wire [WIDTH*2-1+0:0] tmp00_6_31;
	wire [WIDTH*2-1+0:0] tmp00_6_32;
	wire [WIDTH*2-1+0:0] tmp00_6_33;
	wire [WIDTH*2-1+0:0] tmp00_6_34;
	wire [WIDTH*2-1+0:0] tmp00_6_35;
	wire [WIDTH*2-1+0:0] tmp00_6_36;
	wire [WIDTH*2-1+0:0] tmp00_6_37;
	wire [WIDTH*2-1+0:0] tmp00_6_38;
	wire [WIDTH*2-1+0:0] tmp00_6_39;
	wire [WIDTH*2-1+0:0] tmp00_6_40;
	wire [WIDTH*2-1+0:0] tmp00_6_41;
	wire [WIDTH*2-1+0:0] tmp00_6_42;
	wire [WIDTH*2-1+0:0] tmp00_6_43;
	wire [WIDTH*2-1+0:0] tmp00_6_44;
	wire [WIDTH*2-1+0:0] tmp00_6_45;
	wire [WIDTH*2-1+0:0] tmp00_6_46;
	wire [WIDTH*2-1+0:0] tmp00_6_47;
	wire [WIDTH*2-1+0:0] tmp00_6_48;
	wire [WIDTH*2-1+0:0] tmp00_6_49;
	wire [WIDTH*2-1+0:0] tmp00_6_50;
	wire [WIDTH*2-1+0:0] tmp00_6_51;
	wire [WIDTH*2-1+0:0] tmp00_6_52;
	wire [WIDTH*2-1+0:0] tmp00_6_53;
	wire [WIDTH*2-1+0:0] tmp00_6_54;
	wire [WIDTH*2-1+0:0] tmp00_6_55;
	wire [WIDTH*2-1+0:0] tmp00_6_56;
	wire [WIDTH*2-1+0:0] tmp00_6_57;
	wire [WIDTH*2-1+0:0] tmp00_6_58;
	wire [WIDTH*2-1+0:0] tmp00_6_59;
	wire [WIDTH*2-1+0:0] tmp00_6_60;
	wire [WIDTH*2-1+0:0] tmp00_6_61;
	wire [WIDTH*2-1+0:0] tmp00_6_62;
	wire [WIDTH*2-1+0:0] tmp00_6_63;
	wire [WIDTH*2-1+0:0] tmp00_6_64;
	wire [WIDTH*2-1+0:0] tmp00_6_65;
	wire [WIDTH*2-1+0:0] tmp00_6_66;
	wire [WIDTH*2-1+0:0] tmp00_6_67;
	wire [WIDTH*2-1+0:0] tmp00_6_68;
	wire [WIDTH*2-1+0:0] tmp00_6_69;
	wire [WIDTH*2-1+0:0] tmp00_6_70;
	wire [WIDTH*2-1+0:0] tmp00_6_71;
	wire [WIDTH*2-1+0:0] tmp00_6_72;
	wire [WIDTH*2-1+0:0] tmp00_6_73;
	wire [WIDTH*2-1+0:0] tmp00_6_74;
	wire [WIDTH*2-1+0:0] tmp00_6_75;
	wire [WIDTH*2-1+0:0] tmp00_6_76;
	wire [WIDTH*2-1+0:0] tmp00_6_77;
	wire [WIDTH*2-1+0:0] tmp00_6_78;
	wire [WIDTH*2-1+0:0] tmp00_6_79;
	wire [WIDTH*2-1+0:0] tmp00_6_80;
	wire [WIDTH*2-1+0:0] tmp00_6_81;
	wire [WIDTH*2-1+0:0] tmp00_6_82;
	wire [WIDTH*2-1+0:0] tmp00_6_83;
	wire [WIDTH*2-1+0:0] tmp00_7_0;
	wire [WIDTH*2-1+0:0] tmp00_7_1;
	wire [WIDTH*2-1+0:0] tmp00_7_2;
	wire [WIDTH*2-1+0:0] tmp00_7_3;
	wire [WIDTH*2-1+0:0] tmp00_7_4;
	wire [WIDTH*2-1+0:0] tmp00_7_5;
	wire [WIDTH*2-1+0:0] tmp00_7_6;
	wire [WIDTH*2-1+0:0] tmp00_7_7;
	wire [WIDTH*2-1+0:0] tmp00_7_8;
	wire [WIDTH*2-1+0:0] tmp00_7_9;
	wire [WIDTH*2-1+0:0] tmp00_7_10;
	wire [WIDTH*2-1+0:0] tmp00_7_11;
	wire [WIDTH*2-1+0:0] tmp00_7_12;
	wire [WIDTH*2-1+0:0] tmp00_7_13;
	wire [WIDTH*2-1+0:0] tmp00_7_14;
	wire [WIDTH*2-1+0:0] tmp00_7_15;
	wire [WIDTH*2-1+0:0] tmp00_7_16;
	wire [WIDTH*2-1+0:0] tmp00_7_17;
	wire [WIDTH*2-1+0:0] tmp00_7_18;
	wire [WIDTH*2-1+0:0] tmp00_7_19;
	wire [WIDTH*2-1+0:0] tmp00_7_20;
	wire [WIDTH*2-1+0:0] tmp00_7_21;
	wire [WIDTH*2-1+0:0] tmp00_7_22;
	wire [WIDTH*2-1+0:0] tmp00_7_23;
	wire [WIDTH*2-1+0:0] tmp00_7_24;
	wire [WIDTH*2-1+0:0] tmp00_7_25;
	wire [WIDTH*2-1+0:0] tmp00_7_26;
	wire [WIDTH*2-1+0:0] tmp00_7_27;
	wire [WIDTH*2-1+0:0] tmp00_7_28;
	wire [WIDTH*2-1+0:0] tmp00_7_29;
	wire [WIDTH*2-1+0:0] tmp00_7_30;
	wire [WIDTH*2-1+0:0] tmp00_7_31;
	wire [WIDTH*2-1+0:0] tmp00_7_32;
	wire [WIDTH*2-1+0:0] tmp00_7_33;
	wire [WIDTH*2-1+0:0] tmp00_7_34;
	wire [WIDTH*2-1+0:0] tmp00_7_35;
	wire [WIDTH*2-1+0:0] tmp00_7_36;
	wire [WIDTH*2-1+0:0] tmp00_7_37;
	wire [WIDTH*2-1+0:0] tmp00_7_38;
	wire [WIDTH*2-1+0:0] tmp00_7_39;
	wire [WIDTH*2-1+0:0] tmp00_7_40;
	wire [WIDTH*2-1+0:0] tmp00_7_41;
	wire [WIDTH*2-1+0:0] tmp00_7_42;
	wire [WIDTH*2-1+0:0] tmp00_7_43;
	wire [WIDTH*2-1+0:0] tmp00_7_44;
	wire [WIDTH*2-1+0:0] tmp00_7_45;
	wire [WIDTH*2-1+0:0] tmp00_7_46;
	wire [WIDTH*2-1+0:0] tmp00_7_47;
	wire [WIDTH*2-1+0:0] tmp00_7_48;
	wire [WIDTH*2-1+0:0] tmp00_7_49;
	wire [WIDTH*2-1+0:0] tmp00_7_50;
	wire [WIDTH*2-1+0:0] tmp00_7_51;
	wire [WIDTH*2-1+0:0] tmp00_7_52;
	wire [WIDTH*2-1+0:0] tmp00_7_53;
	wire [WIDTH*2-1+0:0] tmp00_7_54;
	wire [WIDTH*2-1+0:0] tmp00_7_55;
	wire [WIDTH*2-1+0:0] tmp00_7_56;
	wire [WIDTH*2-1+0:0] tmp00_7_57;
	wire [WIDTH*2-1+0:0] tmp00_7_58;
	wire [WIDTH*2-1+0:0] tmp00_7_59;
	wire [WIDTH*2-1+0:0] tmp00_7_60;
	wire [WIDTH*2-1+0:0] tmp00_7_61;
	wire [WIDTH*2-1+0:0] tmp00_7_62;
	wire [WIDTH*2-1+0:0] tmp00_7_63;
	wire [WIDTH*2-1+0:0] tmp00_7_64;
	wire [WIDTH*2-1+0:0] tmp00_7_65;
	wire [WIDTH*2-1+0:0] tmp00_7_66;
	wire [WIDTH*2-1+0:0] tmp00_7_67;
	wire [WIDTH*2-1+0:0] tmp00_7_68;
	wire [WIDTH*2-1+0:0] tmp00_7_69;
	wire [WIDTH*2-1+0:0] tmp00_7_70;
	wire [WIDTH*2-1+0:0] tmp00_7_71;
	wire [WIDTH*2-1+0:0] tmp00_7_72;
	wire [WIDTH*2-1+0:0] tmp00_7_73;
	wire [WIDTH*2-1+0:0] tmp00_7_74;
	wire [WIDTH*2-1+0:0] tmp00_7_75;
	wire [WIDTH*2-1+0:0] tmp00_7_76;
	wire [WIDTH*2-1+0:0] tmp00_7_77;
	wire [WIDTH*2-1+0:0] tmp00_7_78;
	wire [WIDTH*2-1+0:0] tmp00_7_79;
	wire [WIDTH*2-1+0:0] tmp00_7_80;
	wire [WIDTH*2-1+0:0] tmp00_7_81;
	wire [WIDTH*2-1+0:0] tmp00_7_82;
	wire [WIDTH*2-1+0:0] tmp00_7_83;
	wire [WIDTH*2-1+0:0] tmp00_8_0;
	wire [WIDTH*2-1+0:0] tmp00_8_1;
	wire [WIDTH*2-1+0:0] tmp00_8_2;
	wire [WIDTH*2-1+0:0] tmp00_8_3;
	wire [WIDTH*2-1+0:0] tmp00_8_4;
	wire [WIDTH*2-1+0:0] tmp00_8_5;
	wire [WIDTH*2-1+0:0] tmp00_8_6;
	wire [WIDTH*2-1+0:0] tmp00_8_7;
	wire [WIDTH*2-1+0:0] tmp00_8_8;
	wire [WIDTH*2-1+0:0] tmp00_8_9;
	wire [WIDTH*2-1+0:0] tmp00_8_10;
	wire [WIDTH*2-1+0:0] tmp00_8_11;
	wire [WIDTH*2-1+0:0] tmp00_8_12;
	wire [WIDTH*2-1+0:0] tmp00_8_13;
	wire [WIDTH*2-1+0:0] tmp00_8_14;
	wire [WIDTH*2-1+0:0] tmp00_8_15;
	wire [WIDTH*2-1+0:0] tmp00_8_16;
	wire [WIDTH*2-1+0:0] tmp00_8_17;
	wire [WIDTH*2-1+0:0] tmp00_8_18;
	wire [WIDTH*2-1+0:0] tmp00_8_19;
	wire [WIDTH*2-1+0:0] tmp00_8_20;
	wire [WIDTH*2-1+0:0] tmp00_8_21;
	wire [WIDTH*2-1+0:0] tmp00_8_22;
	wire [WIDTH*2-1+0:0] tmp00_8_23;
	wire [WIDTH*2-1+0:0] tmp00_8_24;
	wire [WIDTH*2-1+0:0] tmp00_8_25;
	wire [WIDTH*2-1+0:0] tmp00_8_26;
	wire [WIDTH*2-1+0:0] tmp00_8_27;
	wire [WIDTH*2-1+0:0] tmp00_8_28;
	wire [WIDTH*2-1+0:0] tmp00_8_29;
	wire [WIDTH*2-1+0:0] tmp00_8_30;
	wire [WIDTH*2-1+0:0] tmp00_8_31;
	wire [WIDTH*2-1+0:0] tmp00_8_32;
	wire [WIDTH*2-1+0:0] tmp00_8_33;
	wire [WIDTH*2-1+0:0] tmp00_8_34;
	wire [WIDTH*2-1+0:0] tmp00_8_35;
	wire [WIDTH*2-1+0:0] tmp00_8_36;
	wire [WIDTH*2-1+0:0] tmp00_8_37;
	wire [WIDTH*2-1+0:0] tmp00_8_38;
	wire [WIDTH*2-1+0:0] tmp00_8_39;
	wire [WIDTH*2-1+0:0] tmp00_8_40;
	wire [WIDTH*2-1+0:0] tmp00_8_41;
	wire [WIDTH*2-1+0:0] tmp00_8_42;
	wire [WIDTH*2-1+0:0] tmp00_8_43;
	wire [WIDTH*2-1+0:0] tmp00_8_44;
	wire [WIDTH*2-1+0:0] tmp00_8_45;
	wire [WIDTH*2-1+0:0] tmp00_8_46;
	wire [WIDTH*2-1+0:0] tmp00_8_47;
	wire [WIDTH*2-1+0:0] tmp00_8_48;
	wire [WIDTH*2-1+0:0] tmp00_8_49;
	wire [WIDTH*2-1+0:0] tmp00_8_50;
	wire [WIDTH*2-1+0:0] tmp00_8_51;
	wire [WIDTH*2-1+0:0] tmp00_8_52;
	wire [WIDTH*2-1+0:0] tmp00_8_53;
	wire [WIDTH*2-1+0:0] tmp00_8_54;
	wire [WIDTH*2-1+0:0] tmp00_8_55;
	wire [WIDTH*2-1+0:0] tmp00_8_56;
	wire [WIDTH*2-1+0:0] tmp00_8_57;
	wire [WIDTH*2-1+0:0] tmp00_8_58;
	wire [WIDTH*2-1+0:0] tmp00_8_59;
	wire [WIDTH*2-1+0:0] tmp00_8_60;
	wire [WIDTH*2-1+0:0] tmp00_8_61;
	wire [WIDTH*2-1+0:0] tmp00_8_62;
	wire [WIDTH*2-1+0:0] tmp00_8_63;
	wire [WIDTH*2-1+0:0] tmp00_8_64;
	wire [WIDTH*2-1+0:0] tmp00_8_65;
	wire [WIDTH*2-1+0:0] tmp00_8_66;
	wire [WIDTH*2-1+0:0] tmp00_8_67;
	wire [WIDTH*2-1+0:0] tmp00_8_68;
	wire [WIDTH*2-1+0:0] tmp00_8_69;
	wire [WIDTH*2-1+0:0] tmp00_8_70;
	wire [WIDTH*2-1+0:0] tmp00_8_71;
	wire [WIDTH*2-1+0:0] tmp00_8_72;
	wire [WIDTH*2-1+0:0] tmp00_8_73;
	wire [WIDTH*2-1+0:0] tmp00_8_74;
	wire [WIDTH*2-1+0:0] tmp00_8_75;
	wire [WIDTH*2-1+0:0] tmp00_8_76;
	wire [WIDTH*2-1+0:0] tmp00_8_77;
	wire [WIDTH*2-1+0:0] tmp00_8_78;
	wire [WIDTH*2-1+0:0] tmp00_8_79;
	wire [WIDTH*2-1+0:0] tmp00_8_80;
	wire [WIDTH*2-1+0:0] tmp00_8_81;
	wire [WIDTH*2-1+0:0] tmp00_8_82;
	wire [WIDTH*2-1+0:0] tmp00_8_83;
	wire [WIDTH*2-1+0:0] tmp00_9_0;
	wire [WIDTH*2-1+0:0] tmp00_9_1;
	wire [WIDTH*2-1+0:0] tmp00_9_2;
	wire [WIDTH*2-1+0:0] tmp00_9_3;
	wire [WIDTH*2-1+0:0] tmp00_9_4;
	wire [WIDTH*2-1+0:0] tmp00_9_5;
	wire [WIDTH*2-1+0:0] tmp00_9_6;
	wire [WIDTH*2-1+0:0] tmp00_9_7;
	wire [WIDTH*2-1+0:0] tmp00_9_8;
	wire [WIDTH*2-1+0:0] tmp00_9_9;
	wire [WIDTH*2-1+0:0] tmp00_9_10;
	wire [WIDTH*2-1+0:0] tmp00_9_11;
	wire [WIDTH*2-1+0:0] tmp00_9_12;
	wire [WIDTH*2-1+0:0] tmp00_9_13;
	wire [WIDTH*2-1+0:0] tmp00_9_14;
	wire [WIDTH*2-1+0:0] tmp00_9_15;
	wire [WIDTH*2-1+0:0] tmp00_9_16;
	wire [WIDTH*2-1+0:0] tmp00_9_17;
	wire [WIDTH*2-1+0:0] tmp00_9_18;
	wire [WIDTH*2-1+0:0] tmp00_9_19;
	wire [WIDTH*2-1+0:0] tmp00_9_20;
	wire [WIDTH*2-1+0:0] tmp00_9_21;
	wire [WIDTH*2-1+0:0] tmp00_9_22;
	wire [WIDTH*2-1+0:0] tmp00_9_23;
	wire [WIDTH*2-1+0:0] tmp00_9_24;
	wire [WIDTH*2-1+0:0] tmp00_9_25;
	wire [WIDTH*2-1+0:0] tmp00_9_26;
	wire [WIDTH*2-1+0:0] tmp00_9_27;
	wire [WIDTH*2-1+0:0] tmp00_9_28;
	wire [WIDTH*2-1+0:0] tmp00_9_29;
	wire [WIDTH*2-1+0:0] tmp00_9_30;
	wire [WIDTH*2-1+0:0] tmp00_9_31;
	wire [WIDTH*2-1+0:0] tmp00_9_32;
	wire [WIDTH*2-1+0:0] tmp00_9_33;
	wire [WIDTH*2-1+0:0] tmp00_9_34;
	wire [WIDTH*2-1+0:0] tmp00_9_35;
	wire [WIDTH*2-1+0:0] tmp00_9_36;
	wire [WIDTH*2-1+0:0] tmp00_9_37;
	wire [WIDTH*2-1+0:0] tmp00_9_38;
	wire [WIDTH*2-1+0:0] tmp00_9_39;
	wire [WIDTH*2-1+0:0] tmp00_9_40;
	wire [WIDTH*2-1+0:0] tmp00_9_41;
	wire [WIDTH*2-1+0:0] tmp00_9_42;
	wire [WIDTH*2-1+0:0] tmp00_9_43;
	wire [WIDTH*2-1+0:0] tmp00_9_44;
	wire [WIDTH*2-1+0:0] tmp00_9_45;
	wire [WIDTH*2-1+0:0] tmp00_9_46;
	wire [WIDTH*2-1+0:0] tmp00_9_47;
	wire [WIDTH*2-1+0:0] tmp00_9_48;
	wire [WIDTH*2-1+0:0] tmp00_9_49;
	wire [WIDTH*2-1+0:0] tmp00_9_50;
	wire [WIDTH*2-1+0:0] tmp00_9_51;
	wire [WIDTH*2-1+0:0] tmp00_9_52;
	wire [WIDTH*2-1+0:0] tmp00_9_53;
	wire [WIDTH*2-1+0:0] tmp00_9_54;
	wire [WIDTH*2-1+0:0] tmp00_9_55;
	wire [WIDTH*2-1+0:0] tmp00_9_56;
	wire [WIDTH*2-1+0:0] tmp00_9_57;
	wire [WIDTH*2-1+0:0] tmp00_9_58;
	wire [WIDTH*2-1+0:0] tmp00_9_59;
	wire [WIDTH*2-1+0:0] tmp00_9_60;
	wire [WIDTH*2-1+0:0] tmp00_9_61;
	wire [WIDTH*2-1+0:0] tmp00_9_62;
	wire [WIDTH*2-1+0:0] tmp00_9_63;
	wire [WIDTH*2-1+0:0] tmp00_9_64;
	wire [WIDTH*2-1+0:0] tmp00_9_65;
	wire [WIDTH*2-1+0:0] tmp00_9_66;
	wire [WIDTH*2-1+0:0] tmp00_9_67;
	wire [WIDTH*2-1+0:0] tmp00_9_68;
	wire [WIDTH*2-1+0:0] tmp00_9_69;
	wire [WIDTH*2-1+0:0] tmp00_9_70;
	wire [WIDTH*2-1+0:0] tmp00_9_71;
	wire [WIDTH*2-1+0:0] tmp00_9_72;
	wire [WIDTH*2-1+0:0] tmp00_9_73;
	wire [WIDTH*2-1+0:0] tmp00_9_74;
	wire [WIDTH*2-1+0:0] tmp00_9_75;
	wire [WIDTH*2-1+0:0] tmp00_9_76;
	wire [WIDTH*2-1+0:0] tmp00_9_77;
	wire [WIDTH*2-1+0:0] tmp00_9_78;
	wire [WIDTH*2-1+0:0] tmp00_9_79;
	wire [WIDTH*2-1+0:0] tmp00_9_80;
	wire [WIDTH*2-1+0:0] tmp00_9_81;
	wire [WIDTH*2-1+0:0] tmp00_9_82;
	wire [WIDTH*2-1+0:0] tmp00_9_83;
	wire [WIDTH*2-1+0:0] tmp00_10_0;
	wire [WIDTH*2-1+0:0] tmp00_10_1;
	wire [WIDTH*2-1+0:0] tmp00_10_2;
	wire [WIDTH*2-1+0:0] tmp00_10_3;
	wire [WIDTH*2-1+0:0] tmp00_10_4;
	wire [WIDTH*2-1+0:0] tmp00_10_5;
	wire [WIDTH*2-1+0:0] tmp00_10_6;
	wire [WIDTH*2-1+0:0] tmp00_10_7;
	wire [WIDTH*2-1+0:0] tmp00_10_8;
	wire [WIDTH*2-1+0:0] tmp00_10_9;
	wire [WIDTH*2-1+0:0] tmp00_10_10;
	wire [WIDTH*2-1+0:0] tmp00_10_11;
	wire [WIDTH*2-1+0:0] tmp00_10_12;
	wire [WIDTH*2-1+0:0] tmp00_10_13;
	wire [WIDTH*2-1+0:0] tmp00_10_14;
	wire [WIDTH*2-1+0:0] tmp00_10_15;
	wire [WIDTH*2-1+0:0] tmp00_10_16;
	wire [WIDTH*2-1+0:0] tmp00_10_17;
	wire [WIDTH*2-1+0:0] tmp00_10_18;
	wire [WIDTH*2-1+0:0] tmp00_10_19;
	wire [WIDTH*2-1+0:0] tmp00_10_20;
	wire [WIDTH*2-1+0:0] tmp00_10_21;
	wire [WIDTH*2-1+0:0] tmp00_10_22;
	wire [WIDTH*2-1+0:0] tmp00_10_23;
	wire [WIDTH*2-1+0:0] tmp00_10_24;
	wire [WIDTH*2-1+0:0] tmp00_10_25;
	wire [WIDTH*2-1+0:0] tmp00_10_26;
	wire [WIDTH*2-1+0:0] tmp00_10_27;
	wire [WIDTH*2-1+0:0] tmp00_10_28;
	wire [WIDTH*2-1+0:0] tmp00_10_29;
	wire [WIDTH*2-1+0:0] tmp00_10_30;
	wire [WIDTH*2-1+0:0] tmp00_10_31;
	wire [WIDTH*2-1+0:0] tmp00_10_32;
	wire [WIDTH*2-1+0:0] tmp00_10_33;
	wire [WIDTH*2-1+0:0] tmp00_10_34;
	wire [WIDTH*2-1+0:0] tmp00_10_35;
	wire [WIDTH*2-1+0:0] tmp00_10_36;
	wire [WIDTH*2-1+0:0] tmp00_10_37;
	wire [WIDTH*2-1+0:0] tmp00_10_38;
	wire [WIDTH*2-1+0:0] tmp00_10_39;
	wire [WIDTH*2-1+0:0] tmp00_10_40;
	wire [WIDTH*2-1+0:0] tmp00_10_41;
	wire [WIDTH*2-1+0:0] tmp00_10_42;
	wire [WIDTH*2-1+0:0] tmp00_10_43;
	wire [WIDTH*2-1+0:0] tmp00_10_44;
	wire [WIDTH*2-1+0:0] tmp00_10_45;
	wire [WIDTH*2-1+0:0] tmp00_10_46;
	wire [WIDTH*2-1+0:0] tmp00_10_47;
	wire [WIDTH*2-1+0:0] tmp00_10_48;
	wire [WIDTH*2-1+0:0] tmp00_10_49;
	wire [WIDTH*2-1+0:0] tmp00_10_50;
	wire [WIDTH*2-1+0:0] tmp00_10_51;
	wire [WIDTH*2-1+0:0] tmp00_10_52;
	wire [WIDTH*2-1+0:0] tmp00_10_53;
	wire [WIDTH*2-1+0:0] tmp00_10_54;
	wire [WIDTH*2-1+0:0] tmp00_10_55;
	wire [WIDTH*2-1+0:0] tmp00_10_56;
	wire [WIDTH*2-1+0:0] tmp00_10_57;
	wire [WIDTH*2-1+0:0] tmp00_10_58;
	wire [WIDTH*2-1+0:0] tmp00_10_59;
	wire [WIDTH*2-1+0:0] tmp00_10_60;
	wire [WIDTH*2-1+0:0] tmp00_10_61;
	wire [WIDTH*2-1+0:0] tmp00_10_62;
	wire [WIDTH*2-1+0:0] tmp00_10_63;
	wire [WIDTH*2-1+0:0] tmp00_10_64;
	wire [WIDTH*2-1+0:0] tmp00_10_65;
	wire [WIDTH*2-1+0:0] tmp00_10_66;
	wire [WIDTH*2-1+0:0] tmp00_10_67;
	wire [WIDTH*2-1+0:0] tmp00_10_68;
	wire [WIDTH*2-1+0:0] tmp00_10_69;
	wire [WIDTH*2-1+0:0] tmp00_10_70;
	wire [WIDTH*2-1+0:0] tmp00_10_71;
	wire [WIDTH*2-1+0:0] tmp00_10_72;
	wire [WIDTH*2-1+0:0] tmp00_10_73;
	wire [WIDTH*2-1+0:0] tmp00_10_74;
	wire [WIDTH*2-1+0:0] tmp00_10_75;
	wire [WIDTH*2-1+0:0] tmp00_10_76;
	wire [WIDTH*2-1+0:0] tmp00_10_77;
	wire [WIDTH*2-1+0:0] tmp00_10_78;
	wire [WIDTH*2-1+0:0] tmp00_10_79;
	wire [WIDTH*2-1+0:0] tmp00_10_80;
	wire [WIDTH*2-1+0:0] tmp00_10_81;
	wire [WIDTH*2-1+0:0] tmp00_10_82;
	wire [WIDTH*2-1+0:0] tmp00_10_83;
	wire [WIDTH*2-1+0:0] tmp00_11_0;
	wire [WIDTH*2-1+0:0] tmp00_11_1;
	wire [WIDTH*2-1+0:0] tmp00_11_2;
	wire [WIDTH*2-1+0:0] tmp00_11_3;
	wire [WIDTH*2-1+0:0] tmp00_11_4;
	wire [WIDTH*2-1+0:0] tmp00_11_5;
	wire [WIDTH*2-1+0:0] tmp00_11_6;
	wire [WIDTH*2-1+0:0] tmp00_11_7;
	wire [WIDTH*2-1+0:0] tmp00_11_8;
	wire [WIDTH*2-1+0:0] tmp00_11_9;
	wire [WIDTH*2-1+0:0] tmp00_11_10;
	wire [WIDTH*2-1+0:0] tmp00_11_11;
	wire [WIDTH*2-1+0:0] tmp00_11_12;
	wire [WIDTH*2-1+0:0] tmp00_11_13;
	wire [WIDTH*2-1+0:0] tmp00_11_14;
	wire [WIDTH*2-1+0:0] tmp00_11_15;
	wire [WIDTH*2-1+0:0] tmp00_11_16;
	wire [WIDTH*2-1+0:0] tmp00_11_17;
	wire [WIDTH*2-1+0:0] tmp00_11_18;
	wire [WIDTH*2-1+0:0] tmp00_11_19;
	wire [WIDTH*2-1+0:0] tmp00_11_20;
	wire [WIDTH*2-1+0:0] tmp00_11_21;
	wire [WIDTH*2-1+0:0] tmp00_11_22;
	wire [WIDTH*2-1+0:0] tmp00_11_23;
	wire [WIDTH*2-1+0:0] tmp00_11_24;
	wire [WIDTH*2-1+0:0] tmp00_11_25;
	wire [WIDTH*2-1+0:0] tmp00_11_26;
	wire [WIDTH*2-1+0:0] tmp00_11_27;
	wire [WIDTH*2-1+0:0] tmp00_11_28;
	wire [WIDTH*2-1+0:0] tmp00_11_29;
	wire [WIDTH*2-1+0:0] tmp00_11_30;
	wire [WIDTH*2-1+0:0] tmp00_11_31;
	wire [WIDTH*2-1+0:0] tmp00_11_32;
	wire [WIDTH*2-1+0:0] tmp00_11_33;
	wire [WIDTH*2-1+0:0] tmp00_11_34;
	wire [WIDTH*2-1+0:0] tmp00_11_35;
	wire [WIDTH*2-1+0:0] tmp00_11_36;
	wire [WIDTH*2-1+0:0] tmp00_11_37;
	wire [WIDTH*2-1+0:0] tmp00_11_38;
	wire [WIDTH*2-1+0:0] tmp00_11_39;
	wire [WIDTH*2-1+0:0] tmp00_11_40;
	wire [WIDTH*2-1+0:0] tmp00_11_41;
	wire [WIDTH*2-1+0:0] tmp00_11_42;
	wire [WIDTH*2-1+0:0] tmp00_11_43;
	wire [WIDTH*2-1+0:0] tmp00_11_44;
	wire [WIDTH*2-1+0:0] tmp00_11_45;
	wire [WIDTH*2-1+0:0] tmp00_11_46;
	wire [WIDTH*2-1+0:0] tmp00_11_47;
	wire [WIDTH*2-1+0:0] tmp00_11_48;
	wire [WIDTH*2-1+0:0] tmp00_11_49;
	wire [WIDTH*2-1+0:0] tmp00_11_50;
	wire [WIDTH*2-1+0:0] tmp00_11_51;
	wire [WIDTH*2-1+0:0] tmp00_11_52;
	wire [WIDTH*2-1+0:0] tmp00_11_53;
	wire [WIDTH*2-1+0:0] tmp00_11_54;
	wire [WIDTH*2-1+0:0] tmp00_11_55;
	wire [WIDTH*2-1+0:0] tmp00_11_56;
	wire [WIDTH*2-1+0:0] tmp00_11_57;
	wire [WIDTH*2-1+0:0] tmp00_11_58;
	wire [WIDTH*2-1+0:0] tmp00_11_59;
	wire [WIDTH*2-1+0:0] tmp00_11_60;
	wire [WIDTH*2-1+0:0] tmp00_11_61;
	wire [WIDTH*2-1+0:0] tmp00_11_62;
	wire [WIDTH*2-1+0:0] tmp00_11_63;
	wire [WIDTH*2-1+0:0] tmp00_11_64;
	wire [WIDTH*2-1+0:0] tmp00_11_65;
	wire [WIDTH*2-1+0:0] tmp00_11_66;
	wire [WIDTH*2-1+0:0] tmp00_11_67;
	wire [WIDTH*2-1+0:0] tmp00_11_68;
	wire [WIDTH*2-1+0:0] tmp00_11_69;
	wire [WIDTH*2-1+0:0] tmp00_11_70;
	wire [WIDTH*2-1+0:0] tmp00_11_71;
	wire [WIDTH*2-1+0:0] tmp00_11_72;
	wire [WIDTH*2-1+0:0] tmp00_11_73;
	wire [WIDTH*2-1+0:0] tmp00_11_74;
	wire [WIDTH*2-1+0:0] tmp00_11_75;
	wire [WIDTH*2-1+0:0] tmp00_11_76;
	wire [WIDTH*2-1+0:0] tmp00_11_77;
	wire [WIDTH*2-1+0:0] tmp00_11_78;
	wire [WIDTH*2-1+0:0] tmp00_11_79;
	wire [WIDTH*2-1+0:0] tmp00_11_80;
	wire [WIDTH*2-1+0:0] tmp00_11_81;
	wire [WIDTH*2-1+0:0] tmp00_11_82;
	wire [WIDTH*2-1+0:0] tmp00_11_83;
	wire [WIDTH*2-1+0:0] tmp00_12_0;
	wire [WIDTH*2-1+0:0] tmp00_12_1;
	wire [WIDTH*2-1+0:0] tmp00_12_2;
	wire [WIDTH*2-1+0:0] tmp00_12_3;
	wire [WIDTH*2-1+0:0] tmp00_12_4;
	wire [WIDTH*2-1+0:0] tmp00_12_5;
	wire [WIDTH*2-1+0:0] tmp00_12_6;
	wire [WIDTH*2-1+0:0] tmp00_12_7;
	wire [WIDTH*2-1+0:0] tmp00_12_8;
	wire [WIDTH*2-1+0:0] tmp00_12_9;
	wire [WIDTH*2-1+0:0] tmp00_12_10;
	wire [WIDTH*2-1+0:0] tmp00_12_11;
	wire [WIDTH*2-1+0:0] tmp00_12_12;
	wire [WIDTH*2-1+0:0] tmp00_12_13;
	wire [WIDTH*2-1+0:0] tmp00_12_14;
	wire [WIDTH*2-1+0:0] tmp00_12_15;
	wire [WIDTH*2-1+0:0] tmp00_12_16;
	wire [WIDTH*2-1+0:0] tmp00_12_17;
	wire [WIDTH*2-1+0:0] tmp00_12_18;
	wire [WIDTH*2-1+0:0] tmp00_12_19;
	wire [WIDTH*2-1+0:0] tmp00_12_20;
	wire [WIDTH*2-1+0:0] tmp00_12_21;
	wire [WIDTH*2-1+0:0] tmp00_12_22;
	wire [WIDTH*2-1+0:0] tmp00_12_23;
	wire [WIDTH*2-1+0:0] tmp00_12_24;
	wire [WIDTH*2-1+0:0] tmp00_12_25;
	wire [WIDTH*2-1+0:0] tmp00_12_26;
	wire [WIDTH*2-1+0:0] tmp00_12_27;
	wire [WIDTH*2-1+0:0] tmp00_12_28;
	wire [WIDTH*2-1+0:0] tmp00_12_29;
	wire [WIDTH*2-1+0:0] tmp00_12_30;
	wire [WIDTH*2-1+0:0] tmp00_12_31;
	wire [WIDTH*2-1+0:0] tmp00_12_32;
	wire [WIDTH*2-1+0:0] tmp00_12_33;
	wire [WIDTH*2-1+0:0] tmp00_12_34;
	wire [WIDTH*2-1+0:0] tmp00_12_35;
	wire [WIDTH*2-1+0:0] tmp00_12_36;
	wire [WIDTH*2-1+0:0] tmp00_12_37;
	wire [WIDTH*2-1+0:0] tmp00_12_38;
	wire [WIDTH*2-1+0:0] tmp00_12_39;
	wire [WIDTH*2-1+0:0] tmp00_12_40;
	wire [WIDTH*2-1+0:0] tmp00_12_41;
	wire [WIDTH*2-1+0:0] tmp00_12_42;
	wire [WIDTH*2-1+0:0] tmp00_12_43;
	wire [WIDTH*2-1+0:0] tmp00_12_44;
	wire [WIDTH*2-1+0:0] tmp00_12_45;
	wire [WIDTH*2-1+0:0] tmp00_12_46;
	wire [WIDTH*2-1+0:0] tmp00_12_47;
	wire [WIDTH*2-1+0:0] tmp00_12_48;
	wire [WIDTH*2-1+0:0] tmp00_12_49;
	wire [WIDTH*2-1+0:0] tmp00_12_50;
	wire [WIDTH*2-1+0:0] tmp00_12_51;
	wire [WIDTH*2-1+0:0] tmp00_12_52;
	wire [WIDTH*2-1+0:0] tmp00_12_53;
	wire [WIDTH*2-1+0:0] tmp00_12_54;
	wire [WIDTH*2-1+0:0] tmp00_12_55;
	wire [WIDTH*2-1+0:0] tmp00_12_56;
	wire [WIDTH*2-1+0:0] tmp00_12_57;
	wire [WIDTH*2-1+0:0] tmp00_12_58;
	wire [WIDTH*2-1+0:0] tmp00_12_59;
	wire [WIDTH*2-1+0:0] tmp00_12_60;
	wire [WIDTH*2-1+0:0] tmp00_12_61;
	wire [WIDTH*2-1+0:0] tmp00_12_62;
	wire [WIDTH*2-1+0:0] tmp00_12_63;
	wire [WIDTH*2-1+0:0] tmp00_12_64;
	wire [WIDTH*2-1+0:0] tmp00_12_65;
	wire [WIDTH*2-1+0:0] tmp00_12_66;
	wire [WIDTH*2-1+0:0] tmp00_12_67;
	wire [WIDTH*2-1+0:0] tmp00_12_68;
	wire [WIDTH*2-1+0:0] tmp00_12_69;
	wire [WIDTH*2-1+0:0] tmp00_12_70;
	wire [WIDTH*2-1+0:0] tmp00_12_71;
	wire [WIDTH*2-1+0:0] tmp00_12_72;
	wire [WIDTH*2-1+0:0] tmp00_12_73;
	wire [WIDTH*2-1+0:0] tmp00_12_74;
	wire [WIDTH*2-1+0:0] tmp00_12_75;
	wire [WIDTH*2-1+0:0] tmp00_12_76;
	wire [WIDTH*2-1+0:0] tmp00_12_77;
	wire [WIDTH*2-1+0:0] tmp00_12_78;
	wire [WIDTH*2-1+0:0] tmp00_12_79;
	wire [WIDTH*2-1+0:0] tmp00_12_80;
	wire [WIDTH*2-1+0:0] tmp00_12_81;
	wire [WIDTH*2-1+0:0] tmp00_12_82;
	wire [WIDTH*2-1+0:0] tmp00_12_83;
	wire [WIDTH*2-1+0:0] tmp00_13_0;
	wire [WIDTH*2-1+0:0] tmp00_13_1;
	wire [WIDTH*2-1+0:0] tmp00_13_2;
	wire [WIDTH*2-1+0:0] tmp00_13_3;
	wire [WIDTH*2-1+0:0] tmp00_13_4;
	wire [WIDTH*2-1+0:0] tmp00_13_5;
	wire [WIDTH*2-1+0:0] tmp00_13_6;
	wire [WIDTH*2-1+0:0] tmp00_13_7;
	wire [WIDTH*2-1+0:0] tmp00_13_8;
	wire [WIDTH*2-1+0:0] tmp00_13_9;
	wire [WIDTH*2-1+0:0] tmp00_13_10;
	wire [WIDTH*2-1+0:0] tmp00_13_11;
	wire [WIDTH*2-1+0:0] tmp00_13_12;
	wire [WIDTH*2-1+0:0] tmp00_13_13;
	wire [WIDTH*2-1+0:0] tmp00_13_14;
	wire [WIDTH*2-1+0:0] tmp00_13_15;
	wire [WIDTH*2-1+0:0] tmp00_13_16;
	wire [WIDTH*2-1+0:0] tmp00_13_17;
	wire [WIDTH*2-1+0:0] tmp00_13_18;
	wire [WIDTH*2-1+0:0] tmp00_13_19;
	wire [WIDTH*2-1+0:0] tmp00_13_20;
	wire [WIDTH*2-1+0:0] tmp00_13_21;
	wire [WIDTH*2-1+0:0] tmp00_13_22;
	wire [WIDTH*2-1+0:0] tmp00_13_23;
	wire [WIDTH*2-1+0:0] tmp00_13_24;
	wire [WIDTH*2-1+0:0] tmp00_13_25;
	wire [WIDTH*2-1+0:0] tmp00_13_26;
	wire [WIDTH*2-1+0:0] tmp00_13_27;
	wire [WIDTH*2-1+0:0] tmp00_13_28;
	wire [WIDTH*2-1+0:0] tmp00_13_29;
	wire [WIDTH*2-1+0:0] tmp00_13_30;
	wire [WIDTH*2-1+0:0] tmp00_13_31;
	wire [WIDTH*2-1+0:0] tmp00_13_32;
	wire [WIDTH*2-1+0:0] tmp00_13_33;
	wire [WIDTH*2-1+0:0] tmp00_13_34;
	wire [WIDTH*2-1+0:0] tmp00_13_35;
	wire [WIDTH*2-1+0:0] tmp00_13_36;
	wire [WIDTH*2-1+0:0] tmp00_13_37;
	wire [WIDTH*2-1+0:0] tmp00_13_38;
	wire [WIDTH*2-1+0:0] tmp00_13_39;
	wire [WIDTH*2-1+0:0] tmp00_13_40;
	wire [WIDTH*2-1+0:0] tmp00_13_41;
	wire [WIDTH*2-1+0:0] tmp00_13_42;
	wire [WIDTH*2-1+0:0] tmp00_13_43;
	wire [WIDTH*2-1+0:0] tmp00_13_44;
	wire [WIDTH*2-1+0:0] tmp00_13_45;
	wire [WIDTH*2-1+0:0] tmp00_13_46;
	wire [WIDTH*2-1+0:0] tmp00_13_47;
	wire [WIDTH*2-1+0:0] tmp00_13_48;
	wire [WIDTH*2-1+0:0] tmp00_13_49;
	wire [WIDTH*2-1+0:0] tmp00_13_50;
	wire [WIDTH*2-1+0:0] tmp00_13_51;
	wire [WIDTH*2-1+0:0] tmp00_13_52;
	wire [WIDTH*2-1+0:0] tmp00_13_53;
	wire [WIDTH*2-1+0:0] tmp00_13_54;
	wire [WIDTH*2-1+0:0] tmp00_13_55;
	wire [WIDTH*2-1+0:0] tmp00_13_56;
	wire [WIDTH*2-1+0:0] tmp00_13_57;
	wire [WIDTH*2-1+0:0] tmp00_13_58;
	wire [WIDTH*2-1+0:0] tmp00_13_59;
	wire [WIDTH*2-1+0:0] tmp00_13_60;
	wire [WIDTH*2-1+0:0] tmp00_13_61;
	wire [WIDTH*2-1+0:0] tmp00_13_62;
	wire [WIDTH*2-1+0:0] tmp00_13_63;
	wire [WIDTH*2-1+0:0] tmp00_13_64;
	wire [WIDTH*2-1+0:0] tmp00_13_65;
	wire [WIDTH*2-1+0:0] tmp00_13_66;
	wire [WIDTH*2-1+0:0] tmp00_13_67;
	wire [WIDTH*2-1+0:0] tmp00_13_68;
	wire [WIDTH*2-1+0:0] tmp00_13_69;
	wire [WIDTH*2-1+0:0] tmp00_13_70;
	wire [WIDTH*2-1+0:0] tmp00_13_71;
	wire [WIDTH*2-1+0:0] tmp00_13_72;
	wire [WIDTH*2-1+0:0] tmp00_13_73;
	wire [WIDTH*2-1+0:0] tmp00_13_74;
	wire [WIDTH*2-1+0:0] tmp00_13_75;
	wire [WIDTH*2-1+0:0] tmp00_13_76;
	wire [WIDTH*2-1+0:0] tmp00_13_77;
	wire [WIDTH*2-1+0:0] tmp00_13_78;
	wire [WIDTH*2-1+0:0] tmp00_13_79;
	wire [WIDTH*2-1+0:0] tmp00_13_80;
	wire [WIDTH*2-1+0:0] tmp00_13_81;
	wire [WIDTH*2-1+0:0] tmp00_13_82;
	wire [WIDTH*2-1+0:0] tmp00_13_83;
	wire [WIDTH*2-1+0:0] tmp00_14_0;
	wire [WIDTH*2-1+0:0] tmp00_14_1;
	wire [WIDTH*2-1+0:0] tmp00_14_2;
	wire [WIDTH*2-1+0:0] tmp00_14_3;
	wire [WIDTH*2-1+0:0] tmp00_14_4;
	wire [WIDTH*2-1+0:0] tmp00_14_5;
	wire [WIDTH*2-1+0:0] tmp00_14_6;
	wire [WIDTH*2-1+0:0] tmp00_14_7;
	wire [WIDTH*2-1+0:0] tmp00_14_8;
	wire [WIDTH*2-1+0:0] tmp00_14_9;
	wire [WIDTH*2-1+0:0] tmp00_14_10;
	wire [WIDTH*2-1+0:0] tmp00_14_11;
	wire [WIDTH*2-1+0:0] tmp00_14_12;
	wire [WIDTH*2-1+0:0] tmp00_14_13;
	wire [WIDTH*2-1+0:0] tmp00_14_14;
	wire [WIDTH*2-1+0:0] tmp00_14_15;
	wire [WIDTH*2-1+0:0] tmp00_14_16;
	wire [WIDTH*2-1+0:0] tmp00_14_17;
	wire [WIDTH*2-1+0:0] tmp00_14_18;
	wire [WIDTH*2-1+0:0] tmp00_14_19;
	wire [WIDTH*2-1+0:0] tmp00_14_20;
	wire [WIDTH*2-1+0:0] tmp00_14_21;
	wire [WIDTH*2-1+0:0] tmp00_14_22;
	wire [WIDTH*2-1+0:0] tmp00_14_23;
	wire [WIDTH*2-1+0:0] tmp00_14_24;
	wire [WIDTH*2-1+0:0] tmp00_14_25;
	wire [WIDTH*2-1+0:0] tmp00_14_26;
	wire [WIDTH*2-1+0:0] tmp00_14_27;
	wire [WIDTH*2-1+0:0] tmp00_14_28;
	wire [WIDTH*2-1+0:0] tmp00_14_29;
	wire [WIDTH*2-1+0:0] tmp00_14_30;
	wire [WIDTH*2-1+0:0] tmp00_14_31;
	wire [WIDTH*2-1+0:0] tmp00_14_32;
	wire [WIDTH*2-1+0:0] tmp00_14_33;
	wire [WIDTH*2-1+0:0] tmp00_14_34;
	wire [WIDTH*2-1+0:0] tmp00_14_35;
	wire [WIDTH*2-1+0:0] tmp00_14_36;
	wire [WIDTH*2-1+0:0] tmp00_14_37;
	wire [WIDTH*2-1+0:0] tmp00_14_38;
	wire [WIDTH*2-1+0:0] tmp00_14_39;
	wire [WIDTH*2-1+0:0] tmp00_14_40;
	wire [WIDTH*2-1+0:0] tmp00_14_41;
	wire [WIDTH*2-1+0:0] tmp00_14_42;
	wire [WIDTH*2-1+0:0] tmp00_14_43;
	wire [WIDTH*2-1+0:0] tmp00_14_44;
	wire [WIDTH*2-1+0:0] tmp00_14_45;
	wire [WIDTH*2-1+0:0] tmp00_14_46;
	wire [WIDTH*2-1+0:0] tmp00_14_47;
	wire [WIDTH*2-1+0:0] tmp00_14_48;
	wire [WIDTH*2-1+0:0] tmp00_14_49;
	wire [WIDTH*2-1+0:0] tmp00_14_50;
	wire [WIDTH*2-1+0:0] tmp00_14_51;
	wire [WIDTH*2-1+0:0] tmp00_14_52;
	wire [WIDTH*2-1+0:0] tmp00_14_53;
	wire [WIDTH*2-1+0:0] tmp00_14_54;
	wire [WIDTH*2-1+0:0] tmp00_14_55;
	wire [WIDTH*2-1+0:0] tmp00_14_56;
	wire [WIDTH*2-1+0:0] tmp00_14_57;
	wire [WIDTH*2-1+0:0] tmp00_14_58;
	wire [WIDTH*2-1+0:0] tmp00_14_59;
	wire [WIDTH*2-1+0:0] tmp00_14_60;
	wire [WIDTH*2-1+0:0] tmp00_14_61;
	wire [WIDTH*2-1+0:0] tmp00_14_62;
	wire [WIDTH*2-1+0:0] tmp00_14_63;
	wire [WIDTH*2-1+0:0] tmp00_14_64;
	wire [WIDTH*2-1+0:0] tmp00_14_65;
	wire [WIDTH*2-1+0:0] tmp00_14_66;
	wire [WIDTH*2-1+0:0] tmp00_14_67;
	wire [WIDTH*2-1+0:0] tmp00_14_68;
	wire [WIDTH*2-1+0:0] tmp00_14_69;
	wire [WIDTH*2-1+0:0] tmp00_14_70;
	wire [WIDTH*2-1+0:0] tmp00_14_71;
	wire [WIDTH*2-1+0:0] tmp00_14_72;
	wire [WIDTH*2-1+0:0] tmp00_14_73;
	wire [WIDTH*2-1+0:0] tmp00_14_74;
	wire [WIDTH*2-1+0:0] tmp00_14_75;
	wire [WIDTH*2-1+0:0] tmp00_14_76;
	wire [WIDTH*2-1+0:0] tmp00_14_77;
	wire [WIDTH*2-1+0:0] tmp00_14_78;
	wire [WIDTH*2-1+0:0] tmp00_14_79;
	wire [WIDTH*2-1+0:0] tmp00_14_80;
	wire [WIDTH*2-1+0:0] tmp00_14_81;
	wire [WIDTH*2-1+0:0] tmp00_14_82;
	wire [WIDTH*2-1+0:0] tmp00_14_83;
	wire [WIDTH*2-1+0:0] tmp00_15_0;
	wire [WIDTH*2-1+0:0] tmp00_15_1;
	wire [WIDTH*2-1+0:0] tmp00_15_2;
	wire [WIDTH*2-1+0:0] tmp00_15_3;
	wire [WIDTH*2-1+0:0] tmp00_15_4;
	wire [WIDTH*2-1+0:0] tmp00_15_5;
	wire [WIDTH*2-1+0:0] tmp00_15_6;
	wire [WIDTH*2-1+0:0] tmp00_15_7;
	wire [WIDTH*2-1+0:0] tmp00_15_8;
	wire [WIDTH*2-1+0:0] tmp00_15_9;
	wire [WIDTH*2-1+0:0] tmp00_15_10;
	wire [WIDTH*2-1+0:0] tmp00_15_11;
	wire [WIDTH*2-1+0:0] tmp00_15_12;
	wire [WIDTH*2-1+0:0] tmp00_15_13;
	wire [WIDTH*2-1+0:0] tmp00_15_14;
	wire [WIDTH*2-1+0:0] tmp00_15_15;
	wire [WIDTH*2-1+0:0] tmp00_15_16;
	wire [WIDTH*2-1+0:0] tmp00_15_17;
	wire [WIDTH*2-1+0:0] tmp00_15_18;
	wire [WIDTH*2-1+0:0] tmp00_15_19;
	wire [WIDTH*2-1+0:0] tmp00_15_20;
	wire [WIDTH*2-1+0:0] tmp00_15_21;
	wire [WIDTH*2-1+0:0] tmp00_15_22;
	wire [WIDTH*2-1+0:0] tmp00_15_23;
	wire [WIDTH*2-1+0:0] tmp00_15_24;
	wire [WIDTH*2-1+0:0] tmp00_15_25;
	wire [WIDTH*2-1+0:0] tmp00_15_26;
	wire [WIDTH*2-1+0:0] tmp00_15_27;
	wire [WIDTH*2-1+0:0] tmp00_15_28;
	wire [WIDTH*2-1+0:0] tmp00_15_29;
	wire [WIDTH*2-1+0:0] tmp00_15_30;
	wire [WIDTH*2-1+0:0] tmp00_15_31;
	wire [WIDTH*2-1+0:0] tmp00_15_32;
	wire [WIDTH*2-1+0:0] tmp00_15_33;
	wire [WIDTH*2-1+0:0] tmp00_15_34;
	wire [WIDTH*2-1+0:0] tmp00_15_35;
	wire [WIDTH*2-1+0:0] tmp00_15_36;
	wire [WIDTH*2-1+0:0] tmp00_15_37;
	wire [WIDTH*2-1+0:0] tmp00_15_38;
	wire [WIDTH*2-1+0:0] tmp00_15_39;
	wire [WIDTH*2-1+0:0] tmp00_15_40;
	wire [WIDTH*2-1+0:0] tmp00_15_41;
	wire [WIDTH*2-1+0:0] tmp00_15_42;
	wire [WIDTH*2-1+0:0] tmp00_15_43;
	wire [WIDTH*2-1+0:0] tmp00_15_44;
	wire [WIDTH*2-1+0:0] tmp00_15_45;
	wire [WIDTH*2-1+0:0] tmp00_15_46;
	wire [WIDTH*2-1+0:0] tmp00_15_47;
	wire [WIDTH*2-1+0:0] tmp00_15_48;
	wire [WIDTH*2-1+0:0] tmp00_15_49;
	wire [WIDTH*2-1+0:0] tmp00_15_50;
	wire [WIDTH*2-1+0:0] tmp00_15_51;
	wire [WIDTH*2-1+0:0] tmp00_15_52;
	wire [WIDTH*2-1+0:0] tmp00_15_53;
	wire [WIDTH*2-1+0:0] tmp00_15_54;
	wire [WIDTH*2-1+0:0] tmp00_15_55;
	wire [WIDTH*2-1+0:0] tmp00_15_56;
	wire [WIDTH*2-1+0:0] tmp00_15_57;
	wire [WIDTH*2-1+0:0] tmp00_15_58;
	wire [WIDTH*2-1+0:0] tmp00_15_59;
	wire [WIDTH*2-1+0:0] tmp00_15_60;
	wire [WIDTH*2-1+0:0] tmp00_15_61;
	wire [WIDTH*2-1+0:0] tmp00_15_62;
	wire [WIDTH*2-1+0:0] tmp00_15_63;
	wire [WIDTH*2-1+0:0] tmp00_15_64;
	wire [WIDTH*2-1+0:0] tmp00_15_65;
	wire [WIDTH*2-1+0:0] tmp00_15_66;
	wire [WIDTH*2-1+0:0] tmp00_15_67;
	wire [WIDTH*2-1+0:0] tmp00_15_68;
	wire [WIDTH*2-1+0:0] tmp00_15_69;
	wire [WIDTH*2-1+0:0] tmp00_15_70;
	wire [WIDTH*2-1+0:0] tmp00_15_71;
	wire [WIDTH*2-1+0:0] tmp00_15_72;
	wire [WIDTH*2-1+0:0] tmp00_15_73;
	wire [WIDTH*2-1+0:0] tmp00_15_74;
	wire [WIDTH*2-1+0:0] tmp00_15_75;
	wire [WIDTH*2-1+0:0] tmp00_15_76;
	wire [WIDTH*2-1+0:0] tmp00_15_77;
	wire [WIDTH*2-1+0:0] tmp00_15_78;
	wire [WIDTH*2-1+0:0] tmp00_15_79;
	wire [WIDTH*2-1+0:0] tmp00_15_80;
	wire [WIDTH*2-1+0:0] tmp00_15_81;
	wire [WIDTH*2-1+0:0] tmp00_15_82;
	wire [WIDTH*2-1+0:0] tmp00_15_83;
	wire [WIDTH*2-1+0:0] tmp00_16_0;
	wire [WIDTH*2-1+0:0] tmp00_16_1;
	wire [WIDTH*2-1+0:0] tmp00_16_2;
	wire [WIDTH*2-1+0:0] tmp00_16_3;
	wire [WIDTH*2-1+0:0] tmp00_16_4;
	wire [WIDTH*2-1+0:0] tmp00_16_5;
	wire [WIDTH*2-1+0:0] tmp00_16_6;
	wire [WIDTH*2-1+0:0] tmp00_16_7;
	wire [WIDTH*2-1+0:0] tmp00_16_8;
	wire [WIDTH*2-1+0:0] tmp00_16_9;
	wire [WIDTH*2-1+0:0] tmp00_16_10;
	wire [WIDTH*2-1+0:0] tmp00_16_11;
	wire [WIDTH*2-1+0:0] tmp00_16_12;
	wire [WIDTH*2-1+0:0] tmp00_16_13;
	wire [WIDTH*2-1+0:0] tmp00_16_14;
	wire [WIDTH*2-1+0:0] tmp00_16_15;
	wire [WIDTH*2-1+0:0] tmp00_16_16;
	wire [WIDTH*2-1+0:0] tmp00_16_17;
	wire [WIDTH*2-1+0:0] tmp00_16_18;
	wire [WIDTH*2-1+0:0] tmp00_16_19;
	wire [WIDTH*2-1+0:0] tmp00_16_20;
	wire [WIDTH*2-1+0:0] tmp00_16_21;
	wire [WIDTH*2-1+0:0] tmp00_16_22;
	wire [WIDTH*2-1+0:0] tmp00_16_23;
	wire [WIDTH*2-1+0:0] tmp00_16_24;
	wire [WIDTH*2-1+0:0] tmp00_16_25;
	wire [WIDTH*2-1+0:0] tmp00_16_26;
	wire [WIDTH*2-1+0:0] tmp00_16_27;
	wire [WIDTH*2-1+0:0] tmp00_16_28;
	wire [WIDTH*2-1+0:0] tmp00_16_29;
	wire [WIDTH*2-1+0:0] tmp00_16_30;
	wire [WIDTH*2-1+0:0] tmp00_16_31;
	wire [WIDTH*2-1+0:0] tmp00_16_32;
	wire [WIDTH*2-1+0:0] tmp00_16_33;
	wire [WIDTH*2-1+0:0] tmp00_16_34;
	wire [WIDTH*2-1+0:0] tmp00_16_35;
	wire [WIDTH*2-1+0:0] tmp00_16_36;
	wire [WIDTH*2-1+0:0] tmp00_16_37;
	wire [WIDTH*2-1+0:0] tmp00_16_38;
	wire [WIDTH*2-1+0:0] tmp00_16_39;
	wire [WIDTH*2-1+0:0] tmp00_16_40;
	wire [WIDTH*2-1+0:0] tmp00_16_41;
	wire [WIDTH*2-1+0:0] tmp00_16_42;
	wire [WIDTH*2-1+0:0] tmp00_16_43;
	wire [WIDTH*2-1+0:0] tmp00_16_44;
	wire [WIDTH*2-1+0:0] tmp00_16_45;
	wire [WIDTH*2-1+0:0] tmp00_16_46;
	wire [WIDTH*2-1+0:0] tmp00_16_47;
	wire [WIDTH*2-1+0:0] tmp00_16_48;
	wire [WIDTH*2-1+0:0] tmp00_16_49;
	wire [WIDTH*2-1+0:0] tmp00_16_50;
	wire [WIDTH*2-1+0:0] tmp00_16_51;
	wire [WIDTH*2-1+0:0] tmp00_16_52;
	wire [WIDTH*2-1+0:0] tmp00_16_53;
	wire [WIDTH*2-1+0:0] tmp00_16_54;
	wire [WIDTH*2-1+0:0] tmp00_16_55;
	wire [WIDTH*2-1+0:0] tmp00_16_56;
	wire [WIDTH*2-1+0:0] tmp00_16_57;
	wire [WIDTH*2-1+0:0] tmp00_16_58;
	wire [WIDTH*2-1+0:0] tmp00_16_59;
	wire [WIDTH*2-1+0:0] tmp00_16_60;
	wire [WIDTH*2-1+0:0] tmp00_16_61;
	wire [WIDTH*2-1+0:0] tmp00_16_62;
	wire [WIDTH*2-1+0:0] tmp00_16_63;
	wire [WIDTH*2-1+0:0] tmp00_16_64;
	wire [WIDTH*2-1+0:0] tmp00_16_65;
	wire [WIDTH*2-1+0:0] tmp00_16_66;
	wire [WIDTH*2-1+0:0] tmp00_16_67;
	wire [WIDTH*2-1+0:0] tmp00_16_68;
	wire [WIDTH*2-1+0:0] tmp00_16_69;
	wire [WIDTH*2-1+0:0] tmp00_16_70;
	wire [WIDTH*2-1+0:0] tmp00_16_71;
	wire [WIDTH*2-1+0:0] tmp00_16_72;
	wire [WIDTH*2-1+0:0] tmp00_16_73;
	wire [WIDTH*2-1+0:0] tmp00_16_74;
	wire [WIDTH*2-1+0:0] tmp00_16_75;
	wire [WIDTH*2-1+0:0] tmp00_16_76;
	wire [WIDTH*2-1+0:0] tmp00_16_77;
	wire [WIDTH*2-1+0:0] tmp00_16_78;
	wire [WIDTH*2-1+0:0] tmp00_16_79;
	wire [WIDTH*2-1+0:0] tmp00_16_80;
	wire [WIDTH*2-1+0:0] tmp00_16_81;
	wire [WIDTH*2-1+0:0] tmp00_16_82;
	wire [WIDTH*2-1+0:0] tmp00_16_83;
	wire [WIDTH*2-1+0:0] tmp00_17_0;
	wire [WIDTH*2-1+0:0] tmp00_17_1;
	wire [WIDTH*2-1+0:0] tmp00_17_2;
	wire [WIDTH*2-1+0:0] tmp00_17_3;
	wire [WIDTH*2-1+0:0] tmp00_17_4;
	wire [WIDTH*2-1+0:0] tmp00_17_5;
	wire [WIDTH*2-1+0:0] tmp00_17_6;
	wire [WIDTH*2-1+0:0] tmp00_17_7;
	wire [WIDTH*2-1+0:0] tmp00_17_8;
	wire [WIDTH*2-1+0:0] tmp00_17_9;
	wire [WIDTH*2-1+0:0] tmp00_17_10;
	wire [WIDTH*2-1+0:0] tmp00_17_11;
	wire [WIDTH*2-1+0:0] tmp00_17_12;
	wire [WIDTH*2-1+0:0] tmp00_17_13;
	wire [WIDTH*2-1+0:0] tmp00_17_14;
	wire [WIDTH*2-1+0:0] tmp00_17_15;
	wire [WIDTH*2-1+0:0] tmp00_17_16;
	wire [WIDTH*2-1+0:0] tmp00_17_17;
	wire [WIDTH*2-1+0:0] tmp00_17_18;
	wire [WIDTH*2-1+0:0] tmp00_17_19;
	wire [WIDTH*2-1+0:0] tmp00_17_20;
	wire [WIDTH*2-1+0:0] tmp00_17_21;
	wire [WIDTH*2-1+0:0] tmp00_17_22;
	wire [WIDTH*2-1+0:0] tmp00_17_23;
	wire [WIDTH*2-1+0:0] tmp00_17_24;
	wire [WIDTH*2-1+0:0] tmp00_17_25;
	wire [WIDTH*2-1+0:0] tmp00_17_26;
	wire [WIDTH*2-1+0:0] tmp00_17_27;
	wire [WIDTH*2-1+0:0] tmp00_17_28;
	wire [WIDTH*2-1+0:0] tmp00_17_29;
	wire [WIDTH*2-1+0:0] tmp00_17_30;
	wire [WIDTH*2-1+0:0] tmp00_17_31;
	wire [WIDTH*2-1+0:0] tmp00_17_32;
	wire [WIDTH*2-1+0:0] tmp00_17_33;
	wire [WIDTH*2-1+0:0] tmp00_17_34;
	wire [WIDTH*2-1+0:0] tmp00_17_35;
	wire [WIDTH*2-1+0:0] tmp00_17_36;
	wire [WIDTH*2-1+0:0] tmp00_17_37;
	wire [WIDTH*2-1+0:0] tmp00_17_38;
	wire [WIDTH*2-1+0:0] tmp00_17_39;
	wire [WIDTH*2-1+0:0] tmp00_17_40;
	wire [WIDTH*2-1+0:0] tmp00_17_41;
	wire [WIDTH*2-1+0:0] tmp00_17_42;
	wire [WIDTH*2-1+0:0] tmp00_17_43;
	wire [WIDTH*2-1+0:0] tmp00_17_44;
	wire [WIDTH*2-1+0:0] tmp00_17_45;
	wire [WIDTH*2-1+0:0] tmp00_17_46;
	wire [WIDTH*2-1+0:0] tmp00_17_47;
	wire [WIDTH*2-1+0:0] tmp00_17_48;
	wire [WIDTH*2-1+0:0] tmp00_17_49;
	wire [WIDTH*2-1+0:0] tmp00_17_50;
	wire [WIDTH*2-1+0:0] tmp00_17_51;
	wire [WIDTH*2-1+0:0] tmp00_17_52;
	wire [WIDTH*2-1+0:0] tmp00_17_53;
	wire [WIDTH*2-1+0:0] tmp00_17_54;
	wire [WIDTH*2-1+0:0] tmp00_17_55;
	wire [WIDTH*2-1+0:0] tmp00_17_56;
	wire [WIDTH*2-1+0:0] tmp00_17_57;
	wire [WIDTH*2-1+0:0] tmp00_17_58;
	wire [WIDTH*2-1+0:0] tmp00_17_59;
	wire [WIDTH*2-1+0:0] tmp00_17_60;
	wire [WIDTH*2-1+0:0] tmp00_17_61;
	wire [WIDTH*2-1+0:0] tmp00_17_62;
	wire [WIDTH*2-1+0:0] tmp00_17_63;
	wire [WIDTH*2-1+0:0] tmp00_17_64;
	wire [WIDTH*2-1+0:0] tmp00_17_65;
	wire [WIDTH*2-1+0:0] tmp00_17_66;
	wire [WIDTH*2-1+0:0] tmp00_17_67;
	wire [WIDTH*2-1+0:0] tmp00_17_68;
	wire [WIDTH*2-1+0:0] tmp00_17_69;
	wire [WIDTH*2-1+0:0] tmp00_17_70;
	wire [WIDTH*2-1+0:0] tmp00_17_71;
	wire [WIDTH*2-1+0:0] tmp00_17_72;
	wire [WIDTH*2-1+0:0] tmp00_17_73;
	wire [WIDTH*2-1+0:0] tmp00_17_74;
	wire [WIDTH*2-1+0:0] tmp00_17_75;
	wire [WIDTH*2-1+0:0] tmp00_17_76;
	wire [WIDTH*2-1+0:0] tmp00_17_77;
	wire [WIDTH*2-1+0:0] tmp00_17_78;
	wire [WIDTH*2-1+0:0] tmp00_17_79;
	wire [WIDTH*2-1+0:0] tmp00_17_80;
	wire [WIDTH*2-1+0:0] tmp00_17_81;
	wire [WIDTH*2-1+0:0] tmp00_17_82;
	wire [WIDTH*2-1+0:0] tmp00_17_83;
	wire [WIDTH*2-1+0:0] tmp00_18_0;
	wire [WIDTH*2-1+0:0] tmp00_18_1;
	wire [WIDTH*2-1+0:0] tmp00_18_2;
	wire [WIDTH*2-1+0:0] tmp00_18_3;
	wire [WIDTH*2-1+0:0] tmp00_18_4;
	wire [WIDTH*2-1+0:0] tmp00_18_5;
	wire [WIDTH*2-1+0:0] tmp00_18_6;
	wire [WIDTH*2-1+0:0] tmp00_18_7;
	wire [WIDTH*2-1+0:0] tmp00_18_8;
	wire [WIDTH*2-1+0:0] tmp00_18_9;
	wire [WIDTH*2-1+0:0] tmp00_18_10;
	wire [WIDTH*2-1+0:0] tmp00_18_11;
	wire [WIDTH*2-1+0:0] tmp00_18_12;
	wire [WIDTH*2-1+0:0] tmp00_18_13;
	wire [WIDTH*2-1+0:0] tmp00_18_14;
	wire [WIDTH*2-1+0:0] tmp00_18_15;
	wire [WIDTH*2-1+0:0] tmp00_18_16;
	wire [WIDTH*2-1+0:0] tmp00_18_17;
	wire [WIDTH*2-1+0:0] tmp00_18_18;
	wire [WIDTH*2-1+0:0] tmp00_18_19;
	wire [WIDTH*2-1+0:0] tmp00_18_20;
	wire [WIDTH*2-1+0:0] tmp00_18_21;
	wire [WIDTH*2-1+0:0] tmp00_18_22;
	wire [WIDTH*2-1+0:0] tmp00_18_23;
	wire [WIDTH*2-1+0:0] tmp00_18_24;
	wire [WIDTH*2-1+0:0] tmp00_18_25;
	wire [WIDTH*2-1+0:0] tmp00_18_26;
	wire [WIDTH*2-1+0:0] tmp00_18_27;
	wire [WIDTH*2-1+0:0] tmp00_18_28;
	wire [WIDTH*2-1+0:0] tmp00_18_29;
	wire [WIDTH*2-1+0:0] tmp00_18_30;
	wire [WIDTH*2-1+0:0] tmp00_18_31;
	wire [WIDTH*2-1+0:0] tmp00_18_32;
	wire [WIDTH*2-1+0:0] tmp00_18_33;
	wire [WIDTH*2-1+0:0] tmp00_18_34;
	wire [WIDTH*2-1+0:0] tmp00_18_35;
	wire [WIDTH*2-1+0:0] tmp00_18_36;
	wire [WIDTH*2-1+0:0] tmp00_18_37;
	wire [WIDTH*2-1+0:0] tmp00_18_38;
	wire [WIDTH*2-1+0:0] tmp00_18_39;
	wire [WIDTH*2-1+0:0] tmp00_18_40;
	wire [WIDTH*2-1+0:0] tmp00_18_41;
	wire [WIDTH*2-1+0:0] tmp00_18_42;
	wire [WIDTH*2-1+0:0] tmp00_18_43;
	wire [WIDTH*2-1+0:0] tmp00_18_44;
	wire [WIDTH*2-1+0:0] tmp00_18_45;
	wire [WIDTH*2-1+0:0] tmp00_18_46;
	wire [WIDTH*2-1+0:0] tmp00_18_47;
	wire [WIDTH*2-1+0:0] tmp00_18_48;
	wire [WIDTH*2-1+0:0] tmp00_18_49;
	wire [WIDTH*2-1+0:0] tmp00_18_50;
	wire [WIDTH*2-1+0:0] tmp00_18_51;
	wire [WIDTH*2-1+0:0] tmp00_18_52;
	wire [WIDTH*2-1+0:0] tmp00_18_53;
	wire [WIDTH*2-1+0:0] tmp00_18_54;
	wire [WIDTH*2-1+0:0] tmp00_18_55;
	wire [WIDTH*2-1+0:0] tmp00_18_56;
	wire [WIDTH*2-1+0:0] tmp00_18_57;
	wire [WIDTH*2-1+0:0] tmp00_18_58;
	wire [WIDTH*2-1+0:0] tmp00_18_59;
	wire [WIDTH*2-1+0:0] tmp00_18_60;
	wire [WIDTH*2-1+0:0] tmp00_18_61;
	wire [WIDTH*2-1+0:0] tmp00_18_62;
	wire [WIDTH*2-1+0:0] tmp00_18_63;
	wire [WIDTH*2-1+0:0] tmp00_18_64;
	wire [WIDTH*2-1+0:0] tmp00_18_65;
	wire [WIDTH*2-1+0:0] tmp00_18_66;
	wire [WIDTH*2-1+0:0] tmp00_18_67;
	wire [WIDTH*2-1+0:0] tmp00_18_68;
	wire [WIDTH*2-1+0:0] tmp00_18_69;
	wire [WIDTH*2-1+0:0] tmp00_18_70;
	wire [WIDTH*2-1+0:0] tmp00_18_71;
	wire [WIDTH*2-1+0:0] tmp00_18_72;
	wire [WIDTH*2-1+0:0] tmp00_18_73;
	wire [WIDTH*2-1+0:0] tmp00_18_74;
	wire [WIDTH*2-1+0:0] tmp00_18_75;
	wire [WIDTH*2-1+0:0] tmp00_18_76;
	wire [WIDTH*2-1+0:0] tmp00_18_77;
	wire [WIDTH*2-1+0:0] tmp00_18_78;
	wire [WIDTH*2-1+0:0] tmp00_18_79;
	wire [WIDTH*2-1+0:0] tmp00_18_80;
	wire [WIDTH*2-1+0:0] tmp00_18_81;
	wire [WIDTH*2-1+0:0] tmp00_18_82;
	wire [WIDTH*2-1+0:0] tmp00_18_83;
	wire [WIDTH*2-1+0:0] tmp00_19_0;
	wire [WIDTH*2-1+0:0] tmp00_19_1;
	wire [WIDTH*2-1+0:0] tmp00_19_2;
	wire [WIDTH*2-1+0:0] tmp00_19_3;
	wire [WIDTH*2-1+0:0] tmp00_19_4;
	wire [WIDTH*2-1+0:0] tmp00_19_5;
	wire [WIDTH*2-1+0:0] tmp00_19_6;
	wire [WIDTH*2-1+0:0] tmp00_19_7;
	wire [WIDTH*2-1+0:0] tmp00_19_8;
	wire [WIDTH*2-1+0:0] tmp00_19_9;
	wire [WIDTH*2-1+0:0] tmp00_19_10;
	wire [WIDTH*2-1+0:0] tmp00_19_11;
	wire [WIDTH*2-1+0:0] tmp00_19_12;
	wire [WIDTH*2-1+0:0] tmp00_19_13;
	wire [WIDTH*2-1+0:0] tmp00_19_14;
	wire [WIDTH*2-1+0:0] tmp00_19_15;
	wire [WIDTH*2-1+0:0] tmp00_19_16;
	wire [WIDTH*2-1+0:0] tmp00_19_17;
	wire [WIDTH*2-1+0:0] tmp00_19_18;
	wire [WIDTH*2-1+0:0] tmp00_19_19;
	wire [WIDTH*2-1+0:0] tmp00_19_20;
	wire [WIDTH*2-1+0:0] tmp00_19_21;
	wire [WIDTH*2-1+0:0] tmp00_19_22;
	wire [WIDTH*2-1+0:0] tmp00_19_23;
	wire [WIDTH*2-1+0:0] tmp00_19_24;
	wire [WIDTH*2-1+0:0] tmp00_19_25;
	wire [WIDTH*2-1+0:0] tmp00_19_26;
	wire [WIDTH*2-1+0:0] tmp00_19_27;
	wire [WIDTH*2-1+0:0] tmp00_19_28;
	wire [WIDTH*2-1+0:0] tmp00_19_29;
	wire [WIDTH*2-1+0:0] tmp00_19_30;
	wire [WIDTH*2-1+0:0] tmp00_19_31;
	wire [WIDTH*2-1+0:0] tmp00_19_32;
	wire [WIDTH*2-1+0:0] tmp00_19_33;
	wire [WIDTH*2-1+0:0] tmp00_19_34;
	wire [WIDTH*2-1+0:0] tmp00_19_35;
	wire [WIDTH*2-1+0:0] tmp00_19_36;
	wire [WIDTH*2-1+0:0] tmp00_19_37;
	wire [WIDTH*2-1+0:0] tmp00_19_38;
	wire [WIDTH*2-1+0:0] tmp00_19_39;
	wire [WIDTH*2-1+0:0] tmp00_19_40;
	wire [WIDTH*2-1+0:0] tmp00_19_41;
	wire [WIDTH*2-1+0:0] tmp00_19_42;
	wire [WIDTH*2-1+0:0] tmp00_19_43;
	wire [WIDTH*2-1+0:0] tmp00_19_44;
	wire [WIDTH*2-1+0:0] tmp00_19_45;
	wire [WIDTH*2-1+0:0] tmp00_19_46;
	wire [WIDTH*2-1+0:0] tmp00_19_47;
	wire [WIDTH*2-1+0:0] tmp00_19_48;
	wire [WIDTH*2-1+0:0] tmp00_19_49;
	wire [WIDTH*2-1+0:0] tmp00_19_50;
	wire [WIDTH*2-1+0:0] tmp00_19_51;
	wire [WIDTH*2-1+0:0] tmp00_19_52;
	wire [WIDTH*2-1+0:0] tmp00_19_53;
	wire [WIDTH*2-1+0:0] tmp00_19_54;
	wire [WIDTH*2-1+0:0] tmp00_19_55;
	wire [WIDTH*2-1+0:0] tmp00_19_56;
	wire [WIDTH*2-1+0:0] tmp00_19_57;
	wire [WIDTH*2-1+0:0] tmp00_19_58;
	wire [WIDTH*2-1+0:0] tmp00_19_59;
	wire [WIDTH*2-1+0:0] tmp00_19_60;
	wire [WIDTH*2-1+0:0] tmp00_19_61;
	wire [WIDTH*2-1+0:0] tmp00_19_62;
	wire [WIDTH*2-1+0:0] tmp00_19_63;
	wire [WIDTH*2-1+0:0] tmp00_19_64;
	wire [WIDTH*2-1+0:0] tmp00_19_65;
	wire [WIDTH*2-1+0:0] tmp00_19_66;
	wire [WIDTH*2-1+0:0] tmp00_19_67;
	wire [WIDTH*2-1+0:0] tmp00_19_68;
	wire [WIDTH*2-1+0:0] tmp00_19_69;
	wire [WIDTH*2-1+0:0] tmp00_19_70;
	wire [WIDTH*2-1+0:0] tmp00_19_71;
	wire [WIDTH*2-1+0:0] tmp00_19_72;
	wire [WIDTH*2-1+0:0] tmp00_19_73;
	wire [WIDTH*2-1+0:0] tmp00_19_74;
	wire [WIDTH*2-1+0:0] tmp00_19_75;
	wire [WIDTH*2-1+0:0] tmp00_19_76;
	wire [WIDTH*2-1+0:0] tmp00_19_77;
	wire [WIDTH*2-1+0:0] tmp00_19_78;
	wire [WIDTH*2-1+0:0] tmp00_19_79;
	wire [WIDTH*2-1+0:0] tmp00_19_80;
	wire [WIDTH*2-1+0:0] tmp00_19_81;
	wire [WIDTH*2-1+0:0] tmp00_19_82;
	wire [WIDTH*2-1+0:0] tmp00_19_83;
	wire [WIDTH*2-1+0:0] tmp00_20_0;
	wire [WIDTH*2-1+0:0] tmp00_20_1;
	wire [WIDTH*2-1+0:0] tmp00_20_2;
	wire [WIDTH*2-1+0:0] tmp00_20_3;
	wire [WIDTH*2-1+0:0] tmp00_20_4;
	wire [WIDTH*2-1+0:0] tmp00_20_5;
	wire [WIDTH*2-1+0:0] tmp00_20_6;
	wire [WIDTH*2-1+0:0] tmp00_20_7;
	wire [WIDTH*2-1+0:0] tmp00_20_8;
	wire [WIDTH*2-1+0:0] tmp00_20_9;
	wire [WIDTH*2-1+0:0] tmp00_20_10;
	wire [WIDTH*2-1+0:0] tmp00_20_11;
	wire [WIDTH*2-1+0:0] tmp00_20_12;
	wire [WIDTH*2-1+0:0] tmp00_20_13;
	wire [WIDTH*2-1+0:0] tmp00_20_14;
	wire [WIDTH*2-1+0:0] tmp00_20_15;
	wire [WIDTH*2-1+0:0] tmp00_20_16;
	wire [WIDTH*2-1+0:0] tmp00_20_17;
	wire [WIDTH*2-1+0:0] tmp00_20_18;
	wire [WIDTH*2-1+0:0] tmp00_20_19;
	wire [WIDTH*2-1+0:0] tmp00_20_20;
	wire [WIDTH*2-1+0:0] tmp00_20_21;
	wire [WIDTH*2-1+0:0] tmp00_20_22;
	wire [WIDTH*2-1+0:0] tmp00_20_23;
	wire [WIDTH*2-1+0:0] tmp00_20_24;
	wire [WIDTH*2-1+0:0] tmp00_20_25;
	wire [WIDTH*2-1+0:0] tmp00_20_26;
	wire [WIDTH*2-1+0:0] tmp00_20_27;
	wire [WIDTH*2-1+0:0] tmp00_20_28;
	wire [WIDTH*2-1+0:0] tmp00_20_29;
	wire [WIDTH*2-1+0:0] tmp00_20_30;
	wire [WIDTH*2-1+0:0] tmp00_20_31;
	wire [WIDTH*2-1+0:0] tmp00_20_32;
	wire [WIDTH*2-1+0:0] tmp00_20_33;
	wire [WIDTH*2-1+0:0] tmp00_20_34;
	wire [WIDTH*2-1+0:0] tmp00_20_35;
	wire [WIDTH*2-1+0:0] tmp00_20_36;
	wire [WIDTH*2-1+0:0] tmp00_20_37;
	wire [WIDTH*2-1+0:0] tmp00_20_38;
	wire [WIDTH*2-1+0:0] tmp00_20_39;
	wire [WIDTH*2-1+0:0] tmp00_20_40;
	wire [WIDTH*2-1+0:0] tmp00_20_41;
	wire [WIDTH*2-1+0:0] tmp00_20_42;
	wire [WIDTH*2-1+0:0] tmp00_20_43;
	wire [WIDTH*2-1+0:0] tmp00_20_44;
	wire [WIDTH*2-1+0:0] tmp00_20_45;
	wire [WIDTH*2-1+0:0] tmp00_20_46;
	wire [WIDTH*2-1+0:0] tmp00_20_47;
	wire [WIDTH*2-1+0:0] tmp00_20_48;
	wire [WIDTH*2-1+0:0] tmp00_20_49;
	wire [WIDTH*2-1+0:0] tmp00_20_50;
	wire [WIDTH*2-1+0:0] tmp00_20_51;
	wire [WIDTH*2-1+0:0] tmp00_20_52;
	wire [WIDTH*2-1+0:0] tmp00_20_53;
	wire [WIDTH*2-1+0:0] tmp00_20_54;
	wire [WIDTH*2-1+0:0] tmp00_20_55;
	wire [WIDTH*2-1+0:0] tmp00_20_56;
	wire [WIDTH*2-1+0:0] tmp00_20_57;
	wire [WIDTH*2-1+0:0] tmp00_20_58;
	wire [WIDTH*2-1+0:0] tmp00_20_59;
	wire [WIDTH*2-1+0:0] tmp00_20_60;
	wire [WIDTH*2-1+0:0] tmp00_20_61;
	wire [WIDTH*2-1+0:0] tmp00_20_62;
	wire [WIDTH*2-1+0:0] tmp00_20_63;
	wire [WIDTH*2-1+0:0] tmp00_20_64;
	wire [WIDTH*2-1+0:0] tmp00_20_65;
	wire [WIDTH*2-1+0:0] tmp00_20_66;
	wire [WIDTH*2-1+0:0] tmp00_20_67;
	wire [WIDTH*2-1+0:0] tmp00_20_68;
	wire [WIDTH*2-1+0:0] tmp00_20_69;
	wire [WIDTH*2-1+0:0] tmp00_20_70;
	wire [WIDTH*2-1+0:0] tmp00_20_71;
	wire [WIDTH*2-1+0:0] tmp00_20_72;
	wire [WIDTH*2-1+0:0] tmp00_20_73;
	wire [WIDTH*2-1+0:0] tmp00_20_74;
	wire [WIDTH*2-1+0:0] tmp00_20_75;
	wire [WIDTH*2-1+0:0] tmp00_20_76;
	wire [WIDTH*2-1+0:0] tmp00_20_77;
	wire [WIDTH*2-1+0:0] tmp00_20_78;
	wire [WIDTH*2-1+0:0] tmp00_20_79;
	wire [WIDTH*2-1+0:0] tmp00_20_80;
	wire [WIDTH*2-1+0:0] tmp00_20_81;
	wire [WIDTH*2-1+0:0] tmp00_20_82;
	wire [WIDTH*2-1+0:0] tmp00_20_83;
	wire [WIDTH*2-1+0:0] tmp00_21_0;
	wire [WIDTH*2-1+0:0] tmp00_21_1;
	wire [WIDTH*2-1+0:0] tmp00_21_2;
	wire [WIDTH*2-1+0:0] tmp00_21_3;
	wire [WIDTH*2-1+0:0] tmp00_21_4;
	wire [WIDTH*2-1+0:0] tmp00_21_5;
	wire [WIDTH*2-1+0:0] tmp00_21_6;
	wire [WIDTH*2-1+0:0] tmp00_21_7;
	wire [WIDTH*2-1+0:0] tmp00_21_8;
	wire [WIDTH*2-1+0:0] tmp00_21_9;
	wire [WIDTH*2-1+0:0] tmp00_21_10;
	wire [WIDTH*2-1+0:0] tmp00_21_11;
	wire [WIDTH*2-1+0:0] tmp00_21_12;
	wire [WIDTH*2-1+0:0] tmp00_21_13;
	wire [WIDTH*2-1+0:0] tmp00_21_14;
	wire [WIDTH*2-1+0:0] tmp00_21_15;
	wire [WIDTH*2-1+0:0] tmp00_21_16;
	wire [WIDTH*2-1+0:0] tmp00_21_17;
	wire [WIDTH*2-1+0:0] tmp00_21_18;
	wire [WIDTH*2-1+0:0] tmp00_21_19;
	wire [WIDTH*2-1+0:0] tmp00_21_20;
	wire [WIDTH*2-1+0:0] tmp00_21_21;
	wire [WIDTH*2-1+0:0] tmp00_21_22;
	wire [WIDTH*2-1+0:0] tmp00_21_23;
	wire [WIDTH*2-1+0:0] tmp00_21_24;
	wire [WIDTH*2-1+0:0] tmp00_21_25;
	wire [WIDTH*2-1+0:0] tmp00_21_26;
	wire [WIDTH*2-1+0:0] tmp00_21_27;
	wire [WIDTH*2-1+0:0] tmp00_21_28;
	wire [WIDTH*2-1+0:0] tmp00_21_29;
	wire [WIDTH*2-1+0:0] tmp00_21_30;
	wire [WIDTH*2-1+0:0] tmp00_21_31;
	wire [WIDTH*2-1+0:0] tmp00_21_32;
	wire [WIDTH*2-1+0:0] tmp00_21_33;
	wire [WIDTH*2-1+0:0] tmp00_21_34;
	wire [WIDTH*2-1+0:0] tmp00_21_35;
	wire [WIDTH*2-1+0:0] tmp00_21_36;
	wire [WIDTH*2-1+0:0] tmp00_21_37;
	wire [WIDTH*2-1+0:0] tmp00_21_38;
	wire [WIDTH*2-1+0:0] tmp00_21_39;
	wire [WIDTH*2-1+0:0] tmp00_21_40;
	wire [WIDTH*2-1+0:0] tmp00_21_41;
	wire [WIDTH*2-1+0:0] tmp00_21_42;
	wire [WIDTH*2-1+0:0] tmp00_21_43;
	wire [WIDTH*2-1+0:0] tmp00_21_44;
	wire [WIDTH*2-1+0:0] tmp00_21_45;
	wire [WIDTH*2-1+0:0] tmp00_21_46;
	wire [WIDTH*2-1+0:0] tmp00_21_47;
	wire [WIDTH*2-1+0:0] tmp00_21_48;
	wire [WIDTH*2-1+0:0] tmp00_21_49;
	wire [WIDTH*2-1+0:0] tmp00_21_50;
	wire [WIDTH*2-1+0:0] tmp00_21_51;
	wire [WIDTH*2-1+0:0] tmp00_21_52;
	wire [WIDTH*2-1+0:0] tmp00_21_53;
	wire [WIDTH*2-1+0:0] tmp00_21_54;
	wire [WIDTH*2-1+0:0] tmp00_21_55;
	wire [WIDTH*2-1+0:0] tmp00_21_56;
	wire [WIDTH*2-1+0:0] tmp00_21_57;
	wire [WIDTH*2-1+0:0] tmp00_21_58;
	wire [WIDTH*2-1+0:0] tmp00_21_59;
	wire [WIDTH*2-1+0:0] tmp00_21_60;
	wire [WIDTH*2-1+0:0] tmp00_21_61;
	wire [WIDTH*2-1+0:0] tmp00_21_62;
	wire [WIDTH*2-1+0:0] tmp00_21_63;
	wire [WIDTH*2-1+0:0] tmp00_21_64;
	wire [WIDTH*2-1+0:0] tmp00_21_65;
	wire [WIDTH*2-1+0:0] tmp00_21_66;
	wire [WIDTH*2-1+0:0] tmp00_21_67;
	wire [WIDTH*2-1+0:0] tmp00_21_68;
	wire [WIDTH*2-1+0:0] tmp00_21_69;
	wire [WIDTH*2-1+0:0] tmp00_21_70;
	wire [WIDTH*2-1+0:0] tmp00_21_71;
	wire [WIDTH*2-1+0:0] tmp00_21_72;
	wire [WIDTH*2-1+0:0] tmp00_21_73;
	wire [WIDTH*2-1+0:0] tmp00_21_74;
	wire [WIDTH*2-1+0:0] tmp00_21_75;
	wire [WIDTH*2-1+0:0] tmp00_21_76;
	wire [WIDTH*2-1+0:0] tmp00_21_77;
	wire [WIDTH*2-1+0:0] tmp00_21_78;
	wire [WIDTH*2-1+0:0] tmp00_21_79;
	wire [WIDTH*2-1+0:0] tmp00_21_80;
	wire [WIDTH*2-1+0:0] tmp00_21_81;
	wire [WIDTH*2-1+0:0] tmp00_21_82;
	wire [WIDTH*2-1+0:0] tmp00_21_83;
	wire [WIDTH*2-1+0:0] tmp00_22_0;
	wire [WIDTH*2-1+0:0] tmp00_22_1;
	wire [WIDTH*2-1+0:0] tmp00_22_2;
	wire [WIDTH*2-1+0:0] tmp00_22_3;
	wire [WIDTH*2-1+0:0] tmp00_22_4;
	wire [WIDTH*2-1+0:0] tmp00_22_5;
	wire [WIDTH*2-1+0:0] tmp00_22_6;
	wire [WIDTH*2-1+0:0] tmp00_22_7;
	wire [WIDTH*2-1+0:0] tmp00_22_8;
	wire [WIDTH*2-1+0:0] tmp00_22_9;
	wire [WIDTH*2-1+0:0] tmp00_22_10;
	wire [WIDTH*2-1+0:0] tmp00_22_11;
	wire [WIDTH*2-1+0:0] tmp00_22_12;
	wire [WIDTH*2-1+0:0] tmp00_22_13;
	wire [WIDTH*2-1+0:0] tmp00_22_14;
	wire [WIDTH*2-1+0:0] tmp00_22_15;
	wire [WIDTH*2-1+0:0] tmp00_22_16;
	wire [WIDTH*2-1+0:0] tmp00_22_17;
	wire [WIDTH*2-1+0:0] tmp00_22_18;
	wire [WIDTH*2-1+0:0] tmp00_22_19;
	wire [WIDTH*2-1+0:0] tmp00_22_20;
	wire [WIDTH*2-1+0:0] tmp00_22_21;
	wire [WIDTH*2-1+0:0] tmp00_22_22;
	wire [WIDTH*2-1+0:0] tmp00_22_23;
	wire [WIDTH*2-1+0:0] tmp00_22_24;
	wire [WIDTH*2-1+0:0] tmp00_22_25;
	wire [WIDTH*2-1+0:0] tmp00_22_26;
	wire [WIDTH*2-1+0:0] tmp00_22_27;
	wire [WIDTH*2-1+0:0] tmp00_22_28;
	wire [WIDTH*2-1+0:0] tmp00_22_29;
	wire [WIDTH*2-1+0:0] tmp00_22_30;
	wire [WIDTH*2-1+0:0] tmp00_22_31;
	wire [WIDTH*2-1+0:0] tmp00_22_32;
	wire [WIDTH*2-1+0:0] tmp00_22_33;
	wire [WIDTH*2-1+0:0] tmp00_22_34;
	wire [WIDTH*2-1+0:0] tmp00_22_35;
	wire [WIDTH*2-1+0:0] tmp00_22_36;
	wire [WIDTH*2-1+0:0] tmp00_22_37;
	wire [WIDTH*2-1+0:0] tmp00_22_38;
	wire [WIDTH*2-1+0:0] tmp00_22_39;
	wire [WIDTH*2-1+0:0] tmp00_22_40;
	wire [WIDTH*2-1+0:0] tmp00_22_41;
	wire [WIDTH*2-1+0:0] tmp00_22_42;
	wire [WIDTH*2-1+0:0] tmp00_22_43;
	wire [WIDTH*2-1+0:0] tmp00_22_44;
	wire [WIDTH*2-1+0:0] tmp00_22_45;
	wire [WIDTH*2-1+0:0] tmp00_22_46;
	wire [WIDTH*2-1+0:0] tmp00_22_47;
	wire [WIDTH*2-1+0:0] tmp00_22_48;
	wire [WIDTH*2-1+0:0] tmp00_22_49;
	wire [WIDTH*2-1+0:0] tmp00_22_50;
	wire [WIDTH*2-1+0:0] tmp00_22_51;
	wire [WIDTH*2-1+0:0] tmp00_22_52;
	wire [WIDTH*2-1+0:0] tmp00_22_53;
	wire [WIDTH*2-1+0:0] tmp00_22_54;
	wire [WIDTH*2-1+0:0] tmp00_22_55;
	wire [WIDTH*2-1+0:0] tmp00_22_56;
	wire [WIDTH*2-1+0:0] tmp00_22_57;
	wire [WIDTH*2-1+0:0] tmp00_22_58;
	wire [WIDTH*2-1+0:0] tmp00_22_59;
	wire [WIDTH*2-1+0:0] tmp00_22_60;
	wire [WIDTH*2-1+0:0] tmp00_22_61;
	wire [WIDTH*2-1+0:0] tmp00_22_62;
	wire [WIDTH*2-1+0:0] tmp00_22_63;
	wire [WIDTH*2-1+0:0] tmp00_22_64;
	wire [WIDTH*2-1+0:0] tmp00_22_65;
	wire [WIDTH*2-1+0:0] tmp00_22_66;
	wire [WIDTH*2-1+0:0] tmp00_22_67;
	wire [WIDTH*2-1+0:0] tmp00_22_68;
	wire [WIDTH*2-1+0:0] tmp00_22_69;
	wire [WIDTH*2-1+0:0] tmp00_22_70;
	wire [WIDTH*2-1+0:0] tmp00_22_71;
	wire [WIDTH*2-1+0:0] tmp00_22_72;
	wire [WIDTH*2-1+0:0] tmp00_22_73;
	wire [WIDTH*2-1+0:0] tmp00_22_74;
	wire [WIDTH*2-1+0:0] tmp00_22_75;
	wire [WIDTH*2-1+0:0] tmp00_22_76;
	wire [WIDTH*2-1+0:0] tmp00_22_77;
	wire [WIDTH*2-1+0:0] tmp00_22_78;
	wire [WIDTH*2-1+0:0] tmp00_22_79;
	wire [WIDTH*2-1+0:0] tmp00_22_80;
	wire [WIDTH*2-1+0:0] tmp00_22_81;
	wire [WIDTH*2-1+0:0] tmp00_22_82;
	wire [WIDTH*2-1+0:0] tmp00_22_83;
	wire [WIDTH*2-1+0:0] tmp00_23_0;
	wire [WIDTH*2-1+0:0] tmp00_23_1;
	wire [WIDTH*2-1+0:0] tmp00_23_2;
	wire [WIDTH*2-1+0:0] tmp00_23_3;
	wire [WIDTH*2-1+0:0] tmp00_23_4;
	wire [WIDTH*2-1+0:0] tmp00_23_5;
	wire [WIDTH*2-1+0:0] tmp00_23_6;
	wire [WIDTH*2-1+0:0] tmp00_23_7;
	wire [WIDTH*2-1+0:0] tmp00_23_8;
	wire [WIDTH*2-1+0:0] tmp00_23_9;
	wire [WIDTH*2-1+0:0] tmp00_23_10;
	wire [WIDTH*2-1+0:0] tmp00_23_11;
	wire [WIDTH*2-1+0:0] tmp00_23_12;
	wire [WIDTH*2-1+0:0] tmp00_23_13;
	wire [WIDTH*2-1+0:0] tmp00_23_14;
	wire [WIDTH*2-1+0:0] tmp00_23_15;
	wire [WIDTH*2-1+0:0] tmp00_23_16;
	wire [WIDTH*2-1+0:0] tmp00_23_17;
	wire [WIDTH*2-1+0:0] tmp00_23_18;
	wire [WIDTH*2-1+0:0] tmp00_23_19;
	wire [WIDTH*2-1+0:0] tmp00_23_20;
	wire [WIDTH*2-1+0:0] tmp00_23_21;
	wire [WIDTH*2-1+0:0] tmp00_23_22;
	wire [WIDTH*2-1+0:0] tmp00_23_23;
	wire [WIDTH*2-1+0:0] tmp00_23_24;
	wire [WIDTH*2-1+0:0] tmp00_23_25;
	wire [WIDTH*2-1+0:0] tmp00_23_26;
	wire [WIDTH*2-1+0:0] tmp00_23_27;
	wire [WIDTH*2-1+0:0] tmp00_23_28;
	wire [WIDTH*2-1+0:0] tmp00_23_29;
	wire [WIDTH*2-1+0:0] tmp00_23_30;
	wire [WIDTH*2-1+0:0] tmp00_23_31;
	wire [WIDTH*2-1+0:0] tmp00_23_32;
	wire [WIDTH*2-1+0:0] tmp00_23_33;
	wire [WIDTH*2-1+0:0] tmp00_23_34;
	wire [WIDTH*2-1+0:0] tmp00_23_35;
	wire [WIDTH*2-1+0:0] tmp00_23_36;
	wire [WIDTH*2-1+0:0] tmp00_23_37;
	wire [WIDTH*2-1+0:0] tmp00_23_38;
	wire [WIDTH*2-1+0:0] tmp00_23_39;
	wire [WIDTH*2-1+0:0] tmp00_23_40;
	wire [WIDTH*2-1+0:0] tmp00_23_41;
	wire [WIDTH*2-1+0:0] tmp00_23_42;
	wire [WIDTH*2-1+0:0] tmp00_23_43;
	wire [WIDTH*2-1+0:0] tmp00_23_44;
	wire [WIDTH*2-1+0:0] tmp00_23_45;
	wire [WIDTH*2-1+0:0] tmp00_23_46;
	wire [WIDTH*2-1+0:0] tmp00_23_47;
	wire [WIDTH*2-1+0:0] tmp00_23_48;
	wire [WIDTH*2-1+0:0] tmp00_23_49;
	wire [WIDTH*2-1+0:0] tmp00_23_50;
	wire [WIDTH*2-1+0:0] tmp00_23_51;
	wire [WIDTH*2-1+0:0] tmp00_23_52;
	wire [WIDTH*2-1+0:0] tmp00_23_53;
	wire [WIDTH*2-1+0:0] tmp00_23_54;
	wire [WIDTH*2-1+0:0] tmp00_23_55;
	wire [WIDTH*2-1+0:0] tmp00_23_56;
	wire [WIDTH*2-1+0:0] tmp00_23_57;
	wire [WIDTH*2-1+0:0] tmp00_23_58;
	wire [WIDTH*2-1+0:0] tmp00_23_59;
	wire [WIDTH*2-1+0:0] tmp00_23_60;
	wire [WIDTH*2-1+0:0] tmp00_23_61;
	wire [WIDTH*2-1+0:0] tmp00_23_62;
	wire [WIDTH*2-1+0:0] tmp00_23_63;
	wire [WIDTH*2-1+0:0] tmp00_23_64;
	wire [WIDTH*2-1+0:0] tmp00_23_65;
	wire [WIDTH*2-1+0:0] tmp00_23_66;
	wire [WIDTH*2-1+0:0] tmp00_23_67;
	wire [WIDTH*2-1+0:0] tmp00_23_68;
	wire [WIDTH*2-1+0:0] tmp00_23_69;
	wire [WIDTH*2-1+0:0] tmp00_23_70;
	wire [WIDTH*2-1+0:0] tmp00_23_71;
	wire [WIDTH*2-1+0:0] tmp00_23_72;
	wire [WIDTH*2-1+0:0] tmp00_23_73;
	wire [WIDTH*2-1+0:0] tmp00_23_74;
	wire [WIDTH*2-1+0:0] tmp00_23_75;
	wire [WIDTH*2-1+0:0] tmp00_23_76;
	wire [WIDTH*2-1+0:0] tmp00_23_77;
	wire [WIDTH*2-1+0:0] tmp00_23_78;
	wire [WIDTH*2-1+0:0] tmp00_23_79;
	wire [WIDTH*2-1+0:0] tmp00_23_80;
	wire [WIDTH*2-1+0:0] tmp00_23_81;
	wire [WIDTH*2-1+0:0] tmp00_23_82;
	wire [WIDTH*2-1+0:0] tmp00_23_83;
	wire [WIDTH*2-1+0:0] tmp00_24_0;
	wire [WIDTH*2-1+0:0] tmp00_24_1;
	wire [WIDTH*2-1+0:0] tmp00_24_2;
	wire [WIDTH*2-1+0:0] tmp00_24_3;
	wire [WIDTH*2-1+0:0] tmp00_24_4;
	wire [WIDTH*2-1+0:0] tmp00_24_5;
	wire [WIDTH*2-1+0:0] tmp00_24_6;
	wire [WIDTH*2-1+0:0] tmp00_24_7;
	wire [WIDTH*2-1+0:0] tmp00_24_8;
	wire [WIDTH*2-1+0:0] tmp00_24_9;
	wire [WIDTH*2-1+0:0] tmp00_24_10;
	wire [WIDTH*2-1+0:0] tmp00_24_11;
	wire [WIDTH*2-1+0:0] tmp00_24_12;
	wire [WIDTH*2-1+0:0] tmp00_24_13;
	wire [WIDTH*2-1+0:0] tmp00_24_14;
	wire [WIDTH*2-1+0:0] tmp00_24_15;
	wire [WIDTH*2-1+0:0] tmp00_24_16;
	wire [WIDTH*2-1+0:0] tmp00_24_17;
	wire [WIDTH*2-1+0:0] tmp00_24_18;
	wire [WIDTH*2-1+0:0] tmp00_24_19;
	wire [WIDTH*2-1+0:0] tmp00_24_20;
	wire [WIDTH*2-1+0:0] tmp00_24_21;
	wire [WIDTH*2-1+0:0] tmp00_24_22;
	wire [WIDTH*2-1+0:0] tmp00_24_23;
	wire [WIDTH*2-1+0:0] tmp00_24_24;
	wire [WIDTH*2-1+0:0] tmp00_24_25;
	wire [WIDTH*2-1+0:0] tmp00_24_26;
	wire [WIDTH*2-1+0:0] tmp00_24_27;
	wire [WIDTH*2-1+0:0] tmp00_24_28;
	wire [WIDTH*2-1+0:0] tmp00_24_29;
	wire [WIDTH*2-1+0:0] tmp00_24_30;
	wire [WIDTH*2-1+0:0] tmp00_24_31;
	wire [WIDTH*2-1+0:0] tmp00_24_32;
	wire [WIDTH*2-1+0:0] tmp00_24_33;
	wire [WIDTH*2-1+0:0] tmp00_24_34;
	wire [WIDTH*2-1+0:0] tmp00_24_35;
	wire [WIDTH*2-1+0:0] tmp00_24_36;
	wire [WIDTH*2-1+0:0] tmp00_24_37;
	wire [WIDTH*2-1+0:0] tmp00_24_38;
	wire [WIDTH*2-1+0:0] tmp00_24_39;
	wire [WIDTH*2-1+0:0] tmp00_24_40;
	wire [WIDTH*2-1+0:0] tmp00_24_41;
	wire [WIDTH*2-1+0:0] tmp00_24_42;
	wire [WIDTH*2-1+0:0] tmp00_24_43;
	wire [WIDTH*2-1+0:0] tmp00_24_44;
	wire [WIDTH*2-1+0:0] tmp00_24_45;
	wire [WIDTH*2-1+0:0] tmp00_24_46;
	wire [WIDTH*2-1+0:0] tmp00_24_47;
	wire [WIDTH*2-1+0:0] tmp00_24_48;
	wire [WIDTH*2-1+0:0] tmp00_24_49;
	wire [WIDTH*2-1+0:0] tmp00_24_50;
	wire [WIDTH*2-1+0:0] tmp00_24_51;
	wire [WIDTH*2-1+0:0] tmp00_24_52;
	wire [WIDTH*2-1+0:0] tmp00_24_53;
	wire [WIDTH*2-1+0:0] tmp00_24_54;
	wire [WIDTH*2-1+0:0] tmp00_24_55;
	wire [WIDTH*2-1+0:0] tmp00_24_56;
	wire [WIDTH*2-1+0:0] tmp00_24_57;
	wire [WIDTH*2-1+0:0] tmp00_24_58;
	wire [WIDTH*2-1+0:0] tmp00_24_59;
	wire [WIDTH*2-1+0:0] tmp00_24_60;
	wire [WIDTH*2-1+0:0] tmp00_24_61;
	wire [WIDTH*2-1+0:0] tmp00_24_62;
	wire [WIDTH*2-1+0:0] tmp00_24_63;
	wire [WIDTH*2-1+0:0] tmp00_24_64;
	wire [WIDTH*2-1+0:0] tmp00_24_65;
	wire [WIDTH*2-1+0:0] tmp00_24_66;
	wire [WIDTH*2-1+0:0] tmp00_24_67;
	wire [WIDTH*2-1+0:0] tmp00_24_68;
	wire [WIDTH*2-1+0:0] tmp00_24_69;
	wire [WIDTH*2-1+0:0] tmp00_24_70;
	wire [WIDTH*2-1+0:0] tmp00_24_71;
	wire [WIDTH*2-1+0:0] tmp00_24_72;
	wire [WIDTH*2-1+0:0] tmp00_24_73;
	wire [WIDTH*2-1+0:0] tmp00_24_74;
	wire [WIDTH*2-1+0:0] tmp00_24_75;
	wire [WIDTH*2-1+0:0] tmp00_24_76;
	wire [WIDTH*2-1+0:0] tmp00_24_77;
	wire [WIDTH*2-1+0:0] tmp00_24_78;
	wire [WIDTH*2-1+0:0] tmp00_24_79;
	wire [WIDTH*2-1+0:0] tmp00_24_80;
	wire [WIDTH*2-1+0:0] tmp00_24_81;
	wire [WIDTH*2-1+0:0] tmp00_24_82;
	wire [WIDTH*2-1+0:0] tmp00_24_83;
	wire [WIDTH*2-1+0:0] tmp00_25_0;
	wire [WIDTH*2-1+0:0] tmp00_25_1;
	wire [WIDTH*2-1+0:0] tmp00_25_2;
	wire [WIDTH*2-1+0:0] tmp00_25_3;
	wire [WIDTH*2-1+0:0] tmp00_25_4;
	wire [WIDTH*2-1+0:0] tmp00_25_5;
	wire [WIDTH*2-1+0:0] tmp00_25_6;
	wire [WIDTH*2-1+0:0] tmp00_25_7;
	wire [WIDTH*2-1+0:0] tmp00_25_8;
	wire [WIDTH*2-1+0:0] tmp00_25_9;
	wire [WIDTH*2-1+0:0] tmp00_25_10;
	wire [WIDTH*2-1+0:0] tmp00_25_11;
	wire [WIDTH*2-1+0:0] tmp00_25_12;
	wire [WIDTH*2-1+0:0] tmp00_25_13;
	wire [WIDTH*2-1+0:0] tmp00_25_14;
	wire [WIDTH*2-1+0:0] tmp00_25_15;
	wire [WIDTH*2-1+0:0] tmp00_25_16;
	wire [WIDTH*2-1+0:0] tmp00_25_17;
	wire [WIDTH*2-1+0:0] tmp00_25_18;
	wire [WIDTH*2-1+0:0] tmp00_25_19;
	wire [WIDTH*2-1+0:0] tmp00_25_20;
	wire [WIDTH*2-1+0:0] tmp00_25_21;
	wire [WIDTH*2-1+0:0] tmp00_25_22;
	wire [WIDTH*2-1+0:0] tmp00_25_23;
	wire [WIDTH*2-1+0:0] tmp00_25_24;
	wire [WIDTH*2-1+0:0] tmp00_25_25;
	wire [WIDTH*2-1+0:0] tmp00_25_26;
	wire [WIDTH*2-1+0:0] tmp00_25_27;
	wire [WIDTH*2-1+0:0] tmp00_25_28;
	wire [WIDTH*2-1+0:0] tmp00_25_29;
	wire [WIDTH*2-1+0:0] tmp00_25_30;
	wire [WIDTH*2-1+0:0] tmp00_25_31;
	wire [WIDTH*2-1+0:0] tmp00_25_32;
	wire [WIDTH*2-1+0:0] tmp00_25_33;
	wire [WIDTH*2-1+0:0] tmp00_25_34;
	wire [WIDTH*2-1+0:0] tmp00_25_35;
	wire [WIDTH*2-1+0:0] tmp00_25_36;
	wire [WIDTH*2-1+0:0] tmp00_25_37;
	wire [WIDTH*2-1+0:0] tmp00_25_38;
	wire [WIDTH*2-1+0:0] tmp00_25_39;
	wire [WIDTH*2-1+0:0] tmp00_25_40;
	wire [WIDTH*2-1+0:0] tmp00_25_41;
	wire [WIDTH*2-1+0:0] tmp00_25_42;
	wire [WIDTH*2-1+0:0] tmp00_25_43;
	wire [WIDTH*2-1+0:0] tmp00_25_44;
	wire [WIDTH*2-1+0:0] tmp00_25_45;
	wire [WIDTH*2-1+0:0] tmp00_25_46;
	wire [WIDTH*2-1+0:0] tmp00_25_47;
	wire [WIDTH*2-1+0:0] tmp00_25_48;
	wire [WIDTH*2-1+0:0] tmp00_25_49;
	wire [WIDTH*2-1+0:0] tmp00_25_50;
	wire [WIDTH*2-1+0:0] tmp00_25_51;
	wire [WIDTH*2-1+0:0] tmp00_25_52;
	wire [WIDTH*2-1+0:0] tmp00_25_53;
	wire [WIDTH*2-1+0:0] tmp00_25_54;
	wire [WIDTH*2-1+0:0] tmp00_25_55;
	wire [WIDTH*2-1+0:0] tmp00_25_56;
	wire [WIDTH*2-1+0:0] tmp00_25_57;
	wire [WIDTH*2-1+0:0] tmp00_25_58;
	wire [WIDTH*2-1+0:0] tmp00_25_59;
	wire [WIDTH*2-1+0:0] tmp00_25_60;
	wire [WIDTH*2-1+0:0] tmp00_25_61;
	wire [WIDTH*2-1+0:0] tmp00_25_62;
	wire [WIDTH*2-1+0:0] tmp00_25_63;
	wire [WIDTH*2-1+0:0] tmp00_25_64;
	wire [WIDTH*2-1+0:0] tmp00_25_65;
	wire [WIDTH*2-1+0:0] tmp00_25_66;
	wire [WIDTH*2-1+0:0] tmp00_25_67;
	wire [WIDTH*2-1+0:0] tmp00_25_68;
	wire [WIDTH*2-1+0:0] tmp00_25_69;
	wire [WIDTH*2-1+0:0] tmp00_25_70;
	wire [WIDTH*2-1+0:0] tmp00_25_71;
	wire [WIDTH*2-1+0:0] tmp00_25_72;
	wire [WIDTH*2-1+0:0] tmp00_25_73;
	wire [WIDTH*2-1+0:0] tmp00_25_74;
	wire [WIDTH*2-1+0:0] tmp00_25_75;
	wire [WIDTH*2-1+0:0] tmp00_25_76;
	wire [WIDTH*2-1+0:0] tmp00_25_77;
	wire [WIDTH*2-1+0:0] tmp00_25_78;
	wire [WIDTH*2-1+0:0] tmp00_25_79;
	wire [WIDTH*2-1+0:0] tmp00_25_80;
	wire [WIDTH*2-1+0:0] tmp00_25_81;
	wire [WIDTH*2-1+0:0] tmp00_25_82;
	wire [WIDTH*2-1+0:0] tmp00_25_83;
	wire [WIDTH*2-1+0:0] tmp00_26_0;
	wire [WIDTH*2-1+0:0] tmp00_26_1;
	wire [WIDTH*2-1+0:0] tmp00_26_2;
	wire [WIDTH*2-1+0:0] tmp00_26_3;
	wire [WIDTH*2-1+0:0] tmp00_26_4;
	wire [WIDTH*2-1+0:0] tmp00_26_5;
	wire [WIDTH*2-1+0:0] tmp00_26_6;
	wire [WIDTH*2-1+0:0] tmp00_26_7;
	wire [WIDTH*2-1+0:0] tmp00_26_8;
	wire [WIDTH*2-1+0:0] tmp00_26_9;
	wire [WIDTH*2-1+0:0] tmp00_26_10;
	wire [WIDTH*2-1+0:0] tmp00_26_11;
	wire [WIDTH*2-1+0:0] tmp00_26_12;
	wire [WIDTH*2-1+0:0] tmp00_26_13;
	wire [WIDTH*2-1+0:0] tmp00_26_14;
	wire [WIDTH*2-1+0:0] tmp00_26_15;
	wire [WIDTH*2-1+0:0] tmp00_26_16;
	wire [WIDTH*2-1+0:0] tmp00_26_17;
	wire [WIDTH*2-1+0:0] tmp00_26_18;
	wire [WIDTH*2-1+0:0] tmp00_26_19;
	wire [WIDTH*2-1+0:0] tmp00_26_20;
	wire [WIDTH*2-1+0:0] tmp00_26_21;
	wire [WIDTH*2-1+0:0] tmp00_26_22;
	wire [WIDTH*2-1+0:0] tmp00_26_23;
	wire [WIDTH*2-1+0:0] tmp00_26_24;
	wire [WIDTH*2-1+0:0] tmp00_26_25;
	wire [WIDTH*2-1+0:0] tmp00_26_26;
	wire [WIDTH*2-1+0:0] tmp00_26_27;
	wire [WIDTH*2-1+0:0] tmp00_26_28;
	wire [WIDTH*2-1+0:0] tmp00_26_29;
	wire [WIDTH*2-1+0:0] tmp00_26_30;
	wire [WIDTH*2-1+0:0] tmp00_26_31;
	wire [WIDTH*2-1+0:0] tmp00_26_32;
	wire [WIDTH*2-1+0:0] tmp00_26_33;
	wire [WIDTH*2-1+0:0] tmp00_26_34;
	wire [WIDTH*2-1+0:0] tmp00_26_35;
	wire [WIDTH*2-1+0:0] tmp00_26_36;
	wire [WIDTH*2-1+0:0] tmp00_26_37;
	wire [WIDTH*2-1+0:0] tmp00_26_38;
	wire [WIDTH*2-1+0:0] tmp00_26_39;
	wire [WIDTH*2-1+0:0] tmp00_26_40;
	wire [WIDTH*2-1+0:0] tmp00_26_41;
	wire [WIDTH*2-1+0:0] tmp00_26_42;
	wire [WIDTH*2-1+0:0] tmp00_26_43;
	wire [WIDTH*2-1+0:0] tmp00_26_44;
	wire [WIDTH*2-1+0:0] tmp00_26_45;
	wire [WIDTH*2-1+0:0] tmp00_26_46;
	wire [WIDTH*2-1+0:0] tmp00_26_47;
	wire [WIDTH*2-1+0:0] tmp00_26_48;
	wire [WIDTH*2-1+0:0] tmp00_26_49;
	wire [WIDTH*2-1+0:0] tmp00_26_50;
	wire [WIDTH*2-1+0:0] tmp00_26_51;
	wire [WIDTH*2-1+0:0] tmp00_26_52;
	wire [WIDTH*2-1+0:0] tmp00_26_53;
	wire [WIDTH*2-1+0:0] tmp00_26_54;
	wire [WIDTH*2-1+0:0] tmp00_26_55;
	wire [WIDTH*2-1+0:0] tmp00_26_56;
	wire [WIDTH*2-1+0:0] tmp00_26_57;
	wire [WIDTH*2-1+0:0] tmp00_26_58;
	wire [WIDTH*2-1+0:0] tmp00_26_59;
	wire [WIDTH*2-1+0:0] tmp00_26_60;
	wire [WIDTH*2-1+0:0] tmp00_26_61;
	wire [WIDTH*2-1+0:0] tmp00_26_62;
	wire [WIDTH*2-1+0:0] tmp00_26_63;
	wire [WIDTH*2-1+0:0] tmp00_26_64;
	wire [WIDTH*2-1+0:0] tmp00_26_65;
	wire [WIDTH*2-1+0:0] tmp00_26_66;
	wire [WIDTH*2-1+0:0] tmp00_26_67;
	wire [WIDTH*2-1+0:0] tmp00_26_68;
	wire [WIDTH*2-1+0:0] tmp00_26_69;
	wire [WIDTH*2-1+0:0] tmp00_26_70;
	wire [WIDTH*2-1+0:0] tmp00_26_71;
	wire [WIDTH*2-1+0:0] tmp00_26_72;
	wire [WIDTH*2-1+0:0] tmp00_26_73;
	wire [WIDTH*2-1+0:0] tmp00_26_74;
	wire [WIDTH*2-1+0:0] tmp00_26_75;
	wire [WIDTH*2-1+0:0] tmp00_26_76;
	wire [WIDTH*2-1+0:0] tmp00_26_77;
	wire [WIDTH*2-1+0:0] tmp00_26_78;
	wire [WIDTH*2-1+0:0] tmp00_26_79;
	wire [WIDTH*2-1+0:0] tmp00_26_80;
	wire [WIDTH*2-1+0:0] tmp00_26_81;
	wire [WIDTH*2-1+0:0] tmp00_26_82;
	wire [WIDTH*2-1+0:0] tmp00_26_83;
	wire [WIDTH*2-1+0:0] tmp00_27_0;
	wire [WIDTH*2-1+0:0] tmp00_27_1;
	wire [WIDTH*2-1+0:0] tmp00_27_2;
	wire [WIDTH*2-1+0:0] tmp00_27_3;
	wire [WIDTH*2-1+0:0] tmp00_27_4;
	wire [WIDTH*2-1+0:0] tmp00_27_5;
	wire [WIDTH*2-1+0:0] tmp00_27_6;
	wire [WIDTH*2-1+0:0] tmp00_27_7;
	wire [WIDTH*2-1+0:0] tmp00_27_8;
	wire [WIDTH*2-1+0:0] tmp00_27_9;
	wire [WIDTH*2-1+0:0] tmp00_27_10;
	wire [WIDTH*2-1+0:0] tmp00_27_11;
	wire [WIDTH*2-1+0:0] tmp00_27_12;
	wire [WIDTH*2-1+0:0] tmp00_27_13;
	wire [WIDTH*2-1+0:0] tmp00_27_14;
	wire [WIDTH*2-1+0:0] tmp00_27_15;
	wire [WIDTH*2-1+0:0] tmp00_27_16;
	wire [WIDTH*2-1+0:0] tmp00_27_17;
	wire [WIDTH*2-1+0:0] tmp00_27_18;
	wire [WIDTH*2-1+0:0] tmp00_27_19;
	wire [WIDTH*2-1+0:0] tmp00_27_20;
	wire [WIDTH*2-1+0:0] tmp00_27_21;
	wire [WIDTH*2-1+0:0] tmp00_27_22;
	wire [WIDTH*2-1+0:0] tmp00_27_23;
	wire [WIDTH*2-1+0:0] tmp00_27_24;
	wire [WIDTH*2-1+0:0] tmp00_27_25;
	wire [WIDTH*2-1+0:0] tmp00_27_26;
	wire [WIDTH*2-1+0:0] tmp00_27_27;
	wire [WIDTH*2-1+0:0] tmp00_27_28;
	wire [WIDTH*2-1+0:0] tmp00_27_29;
	wire [WIDTH*2-1+0:0] tmp00_27_30;
	wire [WIDTH*2-1+0:0] tmp00_27_31;
	wire [WIDTH*2-1+0:0] tmp00_27_32;
	wire [WIDTH*2-1+0:0] tmp00_27_33;
	wire [WIDTH*2-1+0:0] tmp00_27_34;
	wire [WIDTH*2-1+0:0] tmp00_27_35;
	wire [WIDTH*2-1+0:0] tmp00_27_36;
	wire [WIDTH*2-1+0:0] tmp00_27_37;
	wire [WIDTH*2-1+0:0] tmp00_27_38;
	wire [WIDTH*2-1+0:0] tmp00_27_39;
	wire [WIDTH*2-1+0:0] tmp00_27_40;
	wire [WIDTH*2-1+0:0] tmp00_27_41;
	wire [WIDTH*2-1+0:0] tmp00_27_42;
	wire [WIDTH*2-1+0:0] tmp00_27_43;
	wire [WIDTH*2-1+0:0] tmp00_27_44;
	wire [WIDTH*2-1+0:0] tmp00_27_45;
	wire [WIDTH*2-1+0:0] tmp00_27_46;
	wire [WIDTH*2-1+0:0] tmp00_27_47;
	wire [WIDTH*2-1+0:0] tmp00_27_48;
	wire [WIDTH*2-1+0:0] tmp00_27_49;
	wire [WIDTH*2-1+0:0] tmp00_27_50;
	wire [WIDTH*2-1+0:0] tmp00_27_51;
	wire [WIDTH*2-1+0:0] tmp00_27_52;
	wire [WIDTH*2-1+0:0] tmp00_27_53;
	wire [WIDTH*2-1+0:0] tmp00_27_54;
	wire [WIDTH*2-1+0:0] tmp00_27_55;
	wire [WIDTH*2-1+0:0] tmp00_27_56;
	wire [WIDTH*2-1+0:0] tmp00_27_57;
	wire [WIDTH*2-1+0:0] tmp00_27_58;
	wire [WIDTH*2-1+0:0] tmp00_27_59;
	wire [WIDTH*2-1+0:0] tmp00_27_60;
	wire [WIDTH*2-1+0:0] tmp00_27_61;
	wire [WIDTH*2-1+0:0] tmp00_27_62;
	wire [WIDTH*2-1+0:0] tmp00_27_63;
	wire [WIDTH*2-1+0:0] tmp00_27_64;
	wire [WIDTH*2-1+0:0] tmp00_27_65;
	wire [WIDTH*2-1+0:0] tmp00_27_66;
	wire [WIDTH*2-1+0:0] tmp00_27_67;
	wire [WIDTH*2-1+0:0] tmp00_27_68;
	wire [WIDTH*2-1+0:0] tmp00_27_69;
	wire [WIDTH*2-1+0:0] tmp00_27_70;
	wire [WIDTH*2-1+0:0] tmp00_27_71;
	wire [WIDTH*2-1+0:0] tmp00_27_72;
	wire [WIDTH*2-1+0:0] tmp00_27_73;
	wire [WIDTH*2-1+0:0] tmp00_27_74;
	wire [WIDTH*2-1+0:0] tmp00_27_75;
	wire [WIDTH*2-1+0:0] tmp00_27_76;
	wire [WIDTH*2-1+0:0] tmp00_27_77;
	wire [WIDTH*2-1+0:0] tmp00_27_78;
	wire [WIDTH*2-1+0:0] tmp00_27_79;
	wire [WIDTH*2-1+0:0] tmp00_27_80;
	wire [WIDTH*2-1+0:0] tmp00_27_81;
	wire [WIDTH*2-1+0:0] tmp00_27_82;
	wire [WIDTH*2-1+0:0] tmp00_27_83;
	wire [WIDTH*2-1+0:0] tmp00_28_0;
	wire [WIDTH*2-1+0:0] tmp00_28_1;
	wire [WIDTH*2-1+0:0] tmp00_28_2;
	wire [WIDTH*2-1+0:0] tmp00_28_3;
	wire [WIDTH*2-1+0:0] tmp00_28_4;
	wire [WIDTH*2-1+0:0] tmp00_28_5;
	wire [WIDTH*2-1+0:0] tmp00_28_6;
	wire [WIDTH*2-1+0:0] tmp00_28_7;
	wire [WIDTH*2-1+0:0] tmp00_28_8;
	wire [WIDTH*2-1+0:0] tmp00_28_9;
	wire [WIDTH*2-1+0:0] tmp00_28_10;
	wire [WIDTH*2-1+0:0] tmp00_28_11;
	wire [WIDTH*2-1+0:0] tmp00_28_12;
	wire [WIDTH*2-1+0:0] tmp00_28_13;
	wire [WIDTH*2-1+0:0] tmp00_28_14;
	wire [WIDTH*2-1+0:0] tmp00_28_15;
	wire [WIDTH*2-1+0:0] tmp00_28_16;
	wire [WIDTH*2-1+0:0] tmp00_28_17;
	wire [WIDTH*2-1+0:0] tmp00_28_18;
	wire [WIDTH*2-1+0:0] tmp00_28_19;
	wire [WIDTH*2-1+0:0] tmp00_28_20;
	wire [WIDTH*2-1+0:0] tmp00_28_21;
	wire [WIDTH*2-1+0:0] tmp00_28_22;
	wire [WIDTH*2-1+0:0] tmp00_28_23;
	wire [WIDTH*2-1+0:0] tmp00_28_24;
	wire [WIDTH*2-1+0:0] tmp00_28_25;
	wire [WIDTH*2-1+0:0] tmp00_28_26;
	wire [WIDTH*2-1+0:0] tmp00_28_27;
	wire [WIDTH*2-1+0:0] tmp00_28_28;
	wire [WIDTH*2-1+0:0] tmp00_28_29;
	wire [WIDTH*2-1+0:0] tmp00_28_30;
	wire [WIDTH*2-1+0:0] tmp00_28_31;
	wire [WIDTH*2-1+0:0] tmp00_28_32;
	wire [WIDTH*2-1+0:0] tmp00_28_33;
	wire [WIDTH*2-1+0:0] tmp00_28_34;
	wire [WIDTH*2-1+0:0] tmp00_28_35;
	wire [WIDTH*2-1+0:0] tmp00_28_36;
	wire [WIDTH*2-1+0:0] tmp00_28_37;
	wire [WIDTH*2-1+0:0] tmp00_28_38;
	wire [WIDTH*2-1+0:0] tmp00_28_39;
	wire [WIDTH*2-1+0:0] tmp00_28_40;
	wire [WIDTH*2-1+0:0] tmp00_28_41;
	wire [WIDTH*2-1+0:0] tmp00_28_42;
	wire [WIDTH*2-1+0:0] tmp00_28_43;
	wire [WIDTH*2-1+0:0] tmp00_28_44;
	wire [WIDTH*2-1+0:0] tmp00_28_45;
	wire [WIDTH*2-1+0:0] tmp00_28_46;
	wire [WIDTH*2-1+0:0] tmp00_28_47;
	wire [WIDTH*2-1+0:0] tmp00_28_48;
	wire [WIDTH*2-1+0:0] tmp00_28_49;
	wire [WIDTH*2-1+0:0] tmp00_28_50;
	wire [WIDTH*2-1+0:0] tmp00_28_51;
	wire [WIDTH*2-1+0:0] tmp00_28_52;
	wire [WIDTH*2-1+0:0] tmp00_28_53;
	wire [WIDTH*2-1+0:0] tmp00_28_54;
	wire [WIDTH*2-1+0:0] tmp00_28_55;
	wire [WIDTH*2-1+0:0] tmp00_28_56;
	wire [WIDTH*2-1+0:0] tmp00_28_57;
	wire [WIDTH*2-1+0:0] tmp00_28_58;
	wire [WIDTH*2-1+0:0] tmp00_28_59;
	wire [WIDTH*2-1+0:0] tmp00_28_60;
	wire [WIDTH*2-1+0:0] tmp00_28_61;
	wire [WIDTH*2-1+0:0] tmp00_28_62;
	wire [WIDTH*2-1+0:0] tmp00_28_63;
	wire [WIDTH*2-1+0:0] tmp00_28_64;
	wire [WIDTH*2-1+0:0] tmp00_28_65;
	wire [WIDTH*2-1+0:0] tmp00_28_66;
	wire [WIDTH*2-1+0:0] tmp00_28_67;
	wire [WIDTH*2-1+0:0] tmp00_28_68;
	wire [WIDTH*2-1+0:0] tmp00_28_69;
	wire [WIDTH*2-1+0:0] tmp00_28_70;
	wire [WIDTH*2-1+0:0] tmp00_28_71;
	wire [WIDTH*2-1+0:0] tmp00_28_72;
	wire [WIDTH*2-1+0:0] tmp00_28_73;
	wire [WIDTH*2-1+0:0] tmp00_28_74;
	wire [WIDTH*2-1+0:0] tmp00_28_75;
	wire [WIDTH*2-1+0:0] tmp00_28_76;
	wire [WIDTH*2-1+0:0] tmp00_28_77;
	wire [WIDTH*2-1+0:0] tmp00_28_78;
	wire [WIDTH*2-1+0:0] tmp00_28_79;
	wire [WIDTH*2-1+0:0] tmp00_28_80;
	wire [WIDTH*2-1+0:0] tmp00_28_81;
	wire [WIDTH*2-1+0:0] tmp00_28_82;
	wire [WIDTH*2-1+0:0] tmp00_28_83;
	wire [WIDTH*2-1+0:0] tmp00_29_0;
	wire [WIDTH*2-1+0:0] tmp00_29_1;
	wire [WIDTH*2-1+0:0] tmp00_29_2;
	wire [WIDTH*2-1+0:0] tmp00_29_3;
	wire [WIDTH*2-1+0:0] tmp00_29_4;
	wire [WIDTH*2-1+0:0] tmp00_29_5;
	wire [WIDTH*2-1+0:0] tmp00_29_6;
	wire [WIDTH*2-1+0:0] tmp00_29_7;
	wire [WIDTH*2-1+0:0] tmp00_29_8;
	wire [WIDTH*2-1+0:0] tmp00_29_9;
	wire [WIDTH*2-1+0:0] tmp00_29_10;
	wire [WIDTH*2-1+0:0] tmp00_29_11;
	wire [WIDTH*2-1+0:0] tmp00_29_12;
	wire [WIDTH*2-1+0:0] tmp00_29_13;
	wire [WIDTH*2-1+0:0] tmp00_29_14;
	wire [WIDTH*2-1+0:0] tmp00_29_15;
	wire [WIDTH*2-1+0:0] tmp00_29_16;
	wire [WIDTH*2-1+0:0] tmp00_29_17;
	wire [WIDTH*2-1+0:0] tmp00_29_18;
	wire [WIDTH*2-1+0:0] tmp00_29_19;
	wire [WIDTH*2-1+0:0] tmp00_29_20;
	wire [WIDTH*2-1+0:0] tmp00_29_21;
	wire [WIDTH*2-1+0:0] tmp00_29_22;
	wire [WIDTH*2-1+0:0] tmp00_29_23;
	wire [WIDTH*2-1+0:0] tmp00_29_24;
	wire [WIDTH*2-1+0:0] tmp00_29_25;
	wire [WIDTH*2-1+0:0] tmp00_29_26;
	wire [WIDTH*2-1+0:0] tmp00_29_27;
	wire [WIDTH*2-1+0:0] tmp00_29_28;
	wire [WIDTH*2-1+0:0] tmp00_29_29;
	wire [WIDTH*2-1+0:0] tmp00_29_30;
	wire [WIDTH*2-1+0:0] tmp00_29_31;
	wire [WIDTH*2-1+0:0] tmp00_29_32;
	wire [WIDTH*2-1+0:0] tmp00_29_33;
	wire [WIDTH*2-1+0:0] tmp00_29_34;
	wire [WIDTH*2-1+0:0] tmp00_29_35;
	wire [WIDTH*2-1+0:0] tmp00_29_36;
	wire [WIDTH*2-1+0:0] tmp00_29_37;
	wire [WIDTH*2-1+0:0] tmp00_29_38;
	wire [WIDTH*2-1+0:0] tmp00_29_39;
	wire [WIDTH*2-1+0:0] tmp00_29_40;
	wire [WIDTH*2-1+0:0] tmp00_29_41;
	wire [WIDTH*2-1+0:0] tmp00_29_42;
	wire [WIDTH*2-1+0:0] tmp00_29_43;
	wire [WIDTH*2-1+0:0] tmp00_29_44;
	wire [WIDTH*2-1+0:0] tmp00_29_45;
	wire [WIDTH*2-1+0:0] tmp00_29_46;
	wire [WIDTH*2-1+0:0] tmp00_29_47;
	wire [WIDTH*2-1+0:0] tmp00_29_48;
	wire [WIDTH*2-1+0:0] tmp00_29_49;
	wire [WIDTH*2-1+0:0] tmp00_29_50;
	wire [WIDTH*2-1+0:0] tmp00_29_51;
	wire [WIDTH*2-1+0:0] tmp00_29_52;
	wire [WIDTH*2-1+0:0] tmp00_29_53;
	wire [WIDTH*2-1+0:0] tmp00_29_54;
	wire [WIDTH*2-1+0:0] tmp00_29_55;
	wire [WIDTH*2-1+0:0] tmp00_29_56;
	wire [WIDTH*2-1+0:0] tmp00_29_57;
	wire [WIDTH*2-1+0:0] tmp00_29_58;
	wire [WIDTH*2-1+0:0] tmp00_29_59;
	wire [WIDTH*2-1+0:0] tmp00_29_60;
	wire [WIDTH*2-1+0:0] tmp00_29_61;
	wire [WIDTH*2-1+0:0] tmp00_29_62;
	wire [WIDTH*2-1+0:0] tmp00_29_63;
	wire [WIDTH*2-1+0:0] tmp00_29_64;
	wire [WIDTH*2-1+0:0] tmp00_29_65;
	wire [WIDTH*2-1+0:0] tmp00_29_66;
	wire [WIDTH*2-1+0:0] tmp00_29_67;
	wire [WIDTH*2-1+0:0] tmp00_29_68;
	wire [WIDTH*2-1+0:0] tmp00_29_69;
	wire [WIDTH*2-1+0:0] tmp00_29_70;
	wire [WIDTH*2-1+0:0] tmp00_29_71;
	wire [WIDTH*2-1+0:0] tmp00_29_72;
	wire [WIDTH*2-1+0:0] tmp00_29_73;
	wire [WIDTH*2-1+0:0] tmp00_29_74;
	wire [WIDTH*2-1+0:0] tmp00_29_75;
	wire [WIDTH*2-1+0:0] tmp00_29_76;
	wire [WIDTH*2-1+0:0] tmp00_29_77;
	wire [WIDTH*2-1+0:0] tmp00_29_78;
	wire [WIDTH*2-1+0:0] tmp00_29_79;
	wire [WIDTH*2-1+0:0] tmp00_29_80;
	wire [WIDTH*2-1+0:0] tmp00_29_81;
	wire [WIDTH*2-1+0:0] tmp00_29_82;
	wire [WIDTH*2-1+0:0] tmp00_29_83;
	wire [WIDTH*2-1+0:0] tmp00_30_0;
	wire [WIDTH*2-1+0:0] tmp00_30_1;
	wire [WIDTH*2-1+0:0] tmp00_30_2;
	wire [WIDTH*2-1+0:0] tmp00_30_3;
	wire [WIDTH*2-1+0:0] tmp00_30_4;
	wire [WIDTH*2-1+0:0] tmp00_30_5;
	wire [WIDTH*2-1+0:0] tmp00_30_6;
	wire [WIDTH*2-1+0:0] tmp00_30_7;
	wire [WIDTH*2-1+0:0] tmp00_30_8;
	wire [WIDTH*2-1+0:0] tmp00_30_9;
	wire [WIDTH*2-1+0:0] tmp00_30_10;
	wire [WIDTH*2-1+0:0] tmp00_30_11;
	wire [WIDTH*2-1+0:0] tmp00_30_12;
	wire [WIDTH*2-1+0:0] tmp00_30_13;
	wire [WIDTH*2-1+0:0] tmp00_30_14;
	wire [WIDTH*2-1+0:0] tmp00_30_15;
	wire [WIDTH*2-1+0:0] tmp00_30_16;
	wire [WIDTH*2-1+0:0] tmp00_30_17;
	wire [WIDTH*2-1+0:0] tmp00_30_18;
	wire [WIDTH*2-1+0:0] tmp00_30_19;
	wire [WIDTH*2-1+0:0] tmp00_30_20;
	wire [WIDTH*2-1+0:0] tmp00_30_21;
	wire [WIDTH*2-1+0:0] tmp00_30_22;
	wire [WIDTH*2-1+0:0] tmp00_30_23;
	wire [WIDTH*2-1+0:0] tmp00_30_24;
	wire [WIDTH*2-1+0:0] tmp00_30_25;
	wire [WIDTH*2-1+0:0] tmp00_30_26;
	wire [WIDTH*2-1+0:0] tmp00_30_27;
	wire [WIDTH*2-1+0:0] tmp00_30_28;
	wire [WIDTH*2-1+0:0] tmp00_30_29;
	wire [WIDTH*2-1+0:0] tmp00_30_30;
	wire [WIDTH*2-1+0:0] tmp00_30_31;
	wire [WIDTH*2-1+0:0] tmp00_30_32;
	wire [WIDTH*2-1+0:0] tmp00_30_33;
	wire [WIDTH*2-1+0:0] tmp00_30_34;
	wire [WIDTH*2-1+0:0] tmp00_30_35;
	wire [WIDTH*2-1+0:0] tmp00_30_36;
	wire [WIDTH*2-1+0:0] tmp00_30_37;
	wire [WIDTH*2-1+0:0] tmp00_30_38;
	wire [WIDTH*2-1+0:0] tmp00_30_39;
	wire [WIDTH*2-1+0:0] tmp00_30_40;
	wire [WIDTH*2-1+0:0] tmp00_30_41;
	wire [WIDTH*2-1+0:0] tmp00_30_42;
	wire [WIDTH*2-1+0:0] tmp00_30_43;
	wire [WIDTH*2-1+0:0] tmp00_30_44;
	wire [WIDTH*2-1+0:0] tmp00_30_45;
	wire [WIDTH*2-1+0:0] tmp00_30_46;
	wire [WIDTH*2-1+0:0] tmp00_30_47;
	wire [WIDTH*2-1+0:0] tmp00_30_48;
	wire [WIDTH*2-1+0:0] tmp00_30_49;
	wire [WIDTH*2-1+0:0] tmp00_30_50;
	wire [WIDTH*2-1+0:0] tmp00_30_51;
	wire [WIDTH*2-1+0:0] tmp00_30_52;
	wire [WIDTH*2-1+0:0] tmp00_30_53;
	wire [WIDTH*2-1+0:0] tmp00_30_54;
	wire [WIDTH*2-1+0:0] tmp00_30_55;
	wire [WIDTH*2-1+0:0] tmp00_30_56;
	wire [WIDTH*2-1+0:0] tmp00_30_57;
	wire [WIDTH*2-1+0:0] tmp00_30_58;
	wire [WIDTH*2-1+0:0] tmp00_30_59;
	wire [WIDTH*2-1+0:0] tmp00_30_60;
	wire [WIDTH*2-1+0:0] tmp00_30_61;
	wire [WIDTH*2-1+0:0] tmp00_30_62;
	wire [WIDTH*2-1+0:0] tmp00_30_63;
	wire [WIDTH*2-1+0:0] tmp00_30_64;
	wire [WIDTH*2-1+0:0] tmp00_30_65;
	wire [WIDTH*2-1+0:0] tmp00_30_66;
	wire [WIDTH*2-1+0:0] tmp00_30_67;
	wire [WIDTH*2-1+0:0] tmp00_30_68;
	wire [WIDTH*2-1+0:0] tmp00_30_69;
	wire [WIDTH*2-1+0:0] tmp00_30_70;
	wire [WIDTH*2-1+0:0] tmp00_30_71;
	wire [WIDTH*2-1+0:0] tmp00_30_72;
	wire [WIDTH*2-1+0:0] tmp00_30_73;
	wire [WIDTH*2-1+0:0] tmp00_30_74;
	wire [WIDTH*2-1+0:0] tmp00_30_75;
	wire [WIDTH*2-1+0:0] tmp00_30_76;
	wire [WIDTH*2-1+0:0] tmp00_30_77;
	wire [WIDTH*2-1+0:0] tmp00_30_78;
	wire [WIDTH*2-1+0:0] tmp00_30_79;
	wire [WIDTH*2-1+0:0] tmp00_30_80;
	wire [WIDTH*2-1+0:0] tmp00_30_81;
	wire [WIDTH*2-1+0:0] tmp00_30_82;
	wire [WIDTH*2-1+0:0] tmp00_30_83;
	wire [WIDTH*2-1+0:0] tmp00_31_0;
	wire [WIDTH*2-1+0:0] tmp00_31_1;
	wire [WIDTH*2-1+0:0] tmp00_31_2;
	wire [WIDTH*2-1+0:0] tmp00_31_3;
	wire [WIDTH*2-1+0:0] tmp00_31_4;
	wire [WIDTH*2-1+0:0] tmp00_31_5;
	wire [WIDTH*2-1+0:0] tmp00_31_6;
	wire [WIDTH*2-1+0:0] tmp00_31_7;
	wire [WIDTH*2-1+0:0] tmp00_31_8;
	wire [WIDTH*2-1+0:0] tmp00_31_9;
	wire [WIDTH*2-1+0:0] tmp00_31_10;
	wire [WIDTH*2-1+0:0] tmp00_31_11;
	wire [WIDTH*2-1+0:0] tmp00_31_12;
	wire [WIDTH*2-1+0:0] tmp00_31_13;
	wire [WIDTH*2-1+0:0] tmp00_31_14;
	wire [WIDTH*2-1+0:0] tmp00_31_15;
	wire [WIDTH*2-1+0:0] tmp00_31_16;
	wire [WIDTH*2-1+0:0] tmp00_31_17;
	wire [WIDTH*2-1+0:0] tmp00_31_18;
	wire [WIDTH*2-1+0:0] tmp00_31_19;
	wire [WIDTH*2-1+0:0] tmp00_31_20;
	wire [WIDTH*2-1+0:0] tmp00_31_21;
	wire [WIDTH*2-1+0:0] tmp00_31_22;
	wire [WIDTH*2-1+0:0] tmp00_31_23;
	wire [WIDTH*2-1+0:0] tmp00_31_24;
	wire [WIDTH*2-1+0:0] tmp00_31_25;
	wire [WIDTH*2-1+0:0] tmp00_31_26;
	wire [WIDTH*2-1+0:0] tmp00_31_27;
	wire [WIDTH*2-1+0:0] tmp00_31_28;
	wire [WIDTH*2-1+0:0] tmp00_31_29;
	wire [WIDTH*2-1+0:0] tmp00_31_30;
	wire [WIDTH*2-1+0:0] tmp00_31_31;
	wire [WIDTH*2-1+0:0] tmp00_31_32;
	wire [WIDTH*2-1+0:0] tmp00_31_33;
	wire [WIDTH*2-1+0:0] tmp00_31_34;
	wire [WIDTH*2-1+0:0] tmp00_31_35;
	wire [WIDTH*2-1+0:0] tmp00_31_36;
	wire [WIDTH*2-1+0:0] tmp00_31_37;
	wire [WIDTH*2-1+0:0] tmp00_31_38;
	wire [WIDTH*2-1+0:0] tmp00_31_39;
	wire [WIDTH*2-1+0:0] tmp00_31_40;
	wire [WIDTH*2-1+0:0] tmp00_31_41;
	wire [WIDTH*2-1+0:0] tmp00_31_42;
	wire [WIDTH*2-1+0:0] tmp00_31_43;
	wire [WIDTH*2-1+0:0] tmp00_31_44;
	wire [WIDTH*2-1+0:0] tmp00_31_45;
	wire [WIDTH*2-1+0:0] tmp00_31_46;
	wire [WIDTH*2-1+0:0] tmp00_31_47;
	wire [WIDTH*2-1+0:0] tmp00_31_48;
	wire [WIDTH*2-1+0:0] tmp00_31_49;
	wire [WIDTH*2-1+0:0] tmp00_31_50;
	wire [WIDTH*2-1+0:0] tmp00_31_51;
	wire [WIDTH*2-1+0:0] tmp00_31_52;
	wire [WIDTH*2-1+0:0] tmp00_31_53;
	wire [WIDTH*2-1+0:0] tmp00_31_54;
	wire [WIDTH*2-1+0:0] tmp00_31_55;
	wire [WIDTH*2-1+0:0] tmp00_31_56;
	wire [WIDTH*2-1+0:0] tmp00_31_57;
	wire [WIDTH*2-1+0:0] tmp00_31_58;
	wire [WIDTH*2-1+0:0] tmp00_31_59;
	wire [WIDTH*2-1+0:0] tmp00_31_60;
	wire [WIDTH*2-1+0:0] tmp00_31_61;
	wire [WIDTH*2-1+0:0] tmp00_31_62;
	wire [WIDTH*2-1+0:0] tmp00_31_63;
	wire [WIDTH*2-1+0:0] tmp00_31_64;
	wire [WIDTH*2-1+0:0] tmp00_31_65;
	wire [WIDTH*2-1+0:0] tmp00_31_66;
	wire [WIDTH*2-1+0:0] tmp00_31_67;
	wire [WIDTH*2-1+0:0] tmp00_31_68;
	wire [WIDTH*2-1+0:0] tmp00_31_69;
	wire [WIDTH*2-1+0:0] tmp00_31_70;
	wire [WIDTH*2-1+0:0] tmp00_31_71;
	wire [WIDTH*2-1+0:0] tmp00_31_72;
	wire [WIDTH*2-1+0:0] tmp00_31_73;
	wire [WIDTH*2-1+0:0] tmp00_31_74;
	wire [WIDTH*2-1+0:0] tmp00_31_75;
	wire [WIDTH*2-1+0:0] tmp00_31_76;
	wire [WIDTH*2-1+0:0] tmp00_31_77;
	wire [WIDTH*2-1+0:0] tmp00_31_78;
	wire [WIDTH*2-1+0:0] tmp00_31_79;
	wire [WIDTH*2-1+0:0] tmp00_31_80;
	wire [WIDTH*2-1+0:0] tmp00_31_81;
	wire [WIDTH*2-1+0:0] tmp00_31_82;
	wire [WIDTH*2-1+0:0] tmp00_31_83;
	wire [WIDTH*2-1+0:0] tmp00_32_0;
	wire [WIDTH*2-1+0:0] tmp00_32_1;
	wire [WIDTH*2-1+0:0] tmp00_32_2;
	wire [WIDTH*2-1+0:0] tmp00_32_3;
	wire [WIDTH*2-1+0:0] tmp00_32_4;
	wire [WIDTH*2-1+0:0] tmp00_32_5;
	wire [WIDTH*2-1+0:0] tmp00_32_6;
	wire [WIDTH*2-1+0:0] tmp00_32_7;
	wire [WIDTH*2-1+0:0] tmp00_32_8;
	wire [WIDTH*2-1+0:0] tmp00_32_9;
	wire [WIDTH*2-1+0:0] tmp00_32_10;
	wire [WIDTH*2-1+0:0] tmp00_32_11;
	wire [WIDTH*2-1+0:0] tmp00_32_12;
	wire [WIDTH*2-1+0:0] tmp00_32_13;
	wire [WIDTH*2-1+0:0] tmp00_32_14;
	wire [WIDTH*2-1+0:0] tmp00_32_15;
	wire [WIDTH*2-1+0:0] tmp00_32_16;
	wire [WIDTH*2-1+0:0] tmp00_32_17;
	wire [WIDTH*2-1+0:0] tmp00_32_18;
	wire [WIDTH*2-1+0:0] tmp00_32_19;
	wire [WIDTH*2-1+0:0] tmp00_32_20;
	wire [WIDTH*2-1+0:0] tmp00_32_21;
	wire [WIDTH*2-1+0:0] tmp00_32_22;
	wire [WIDTH*2-1+0:0] tmp00_32_23;
	wire [WIDTH*2-1+0:0] tmp00_32_24;
	wire [WIDTH*2-1+0:0] tmp00_32_25;
	wire [WIDTH*2-1+0:0] tmp00_32_26;
	wire [WIDTH*2-1+0:0] tmp00_32_27;
	wire [WIDTH*2-1+0:0] tmp00_32_28;
	wire [WIDTH*2-1+0:0] tmp00_32_29;
	wire [WIDTH*2-1+0:0] tmp00_32_30;
	wire [WIDTH*2-1+0:0] tmp00_32_31;
	wire [WIDTH*2-1+0:0] tmp00_32_32;
	wire [WIDTH*2-1+0:0] tmp00_32_33;
	wire [WIDTH*2-1+0:0] tmp00_32_34;
	wire [WIDTH*2-1+0:0] tmp00_32_35;
	wire [WIDTH*2-1+0:0] tmp00_32_36;
	wire [WIDTH*2-1+0:0] tmp00_32_37;
	wire [WIDTH*2-1+0:0] tmp00_32_38;
	wire [WIDTH*2-1+0:0] tmp00_32_39;
	wire [WIDTH*2-1+0:0] tmp00_32_40;
	wire [WIDTH*2-1+0:0] tmp00_32_41;
	wire [WIDTH*2-1+0:0] tmp00_32_42;
	wire [WIDTH*2-1+0:0] tmp00_32_43;
	wire [WIDTH*2-1+0:0] tmp00_32_44;
	wire [WIDTH*2-1+0:0] tmp00_32_45;
	wire [WIDTH*2-1+0:0] tmp00_32_46;
	wire [WIDTH*2-1+0:0] tmp00_32_47;
	wire [WIDTH*2-1+0:0] tmp00_32_48;
	wire [WIDTH*2-1+0:0] tmp00_32_49;
	wire [WIDTH*2-1+0:0] tmp00_32_50;
	wire [WIDTH*2-1+0:0] tmp00_32_51;
	wire [WIDTH*2-1+0:0] tmp00_32_52;
	wire [WIDTH*2-1+0:0] tmp00_32_53;
	wire [WIDTH*2-1+0:0] tmp00_32_54;
	wire [WIDTH*2-1+0:0] tmp00_32_55;
	wire [WIDTH*2-1+0:0] tmp00_32_56;
	wire [WIDTH*2-1+0:0] tmp00_32_57;
	wire [WIDTH*2-1+0:0] tmp00_32_58;
	wire [WIDTH*2-1+0:0] tmp00_32_59;
	wire [WIDTH*2-1+0:0] tmp00_32_60;
	wire [WIDTH*2-1+0:0] tmp00_32_61;
	wire [WIDTH*2-1+0:0] tmp00_32_62;
	wire [WIDTH*2-1+0:0] tmp00_32_63;
	wire [WIDTH*2-1+0:0] tmp00_32_64;
	wire [WIDTH*2-1+0:0] tmp00_32_65;
	wire [WIDTH*2-1+0:0] tmp00_32_66;
	wire [WIDTH*2-1+0:0] tmp00_32_67;
	wire [WIDTH*2-1+0:0] tmp00_32_68;
	wire [WIDTH*2-1+0:0] tmp00_32_69;
	wire [WIDTH*2-1+0:0] tmp00_32_70;
	wire [WIDTH*2-1+0:0] tmp00_32_71;
	wire [WIDTH*2-1+0:0] tmp00_32_72;
	wire [WIDTH*2-1+0:0] tmp00_32_73;
	wire [WIDTH*2-1+0:0] tmp00_32_74;
	wire [WIDTH*2-1+0:0] tmp00_32_75;
	wire [WIDTH*2-1+0:0] tmp00_32_76;
	wire [WIDTH*2-1+0:0] tmp00_32_77;
	wire [WIDTH*2-1+0:0] tmp00_32_78;
	wire [WIDTH*2-1+0:0] tmp00_32_79;
	wire [WIDTH*2-1+0:0] tmp00_32_80;
	wire [WIDTH*2-1+0:0] tmp00_32_81;
	wire [WIDTH*2-1+0:0] tmp00_32_82;
	wire [WIDTH*2-1+0:0] tmp00_32_83;
	wire [WIDTH*2-1+0:0] tmp00_33_0;
	wire [WIDTH*2-1+0:0] tmp00_33_1;
	wire [WIDTH*2-1+0:0] tmp00_33_2;
	wire [WIDTH*2-1+0:0] tmp00_33_3;
	wire [WIDTH*2-1+0:0] tmp00_33_4;
	wire [WIDTH*2-1+0:0] tmp00_33_5;
	wire [WIDTH*2-1+0:0] tmp00_33_6;
	wire [WIDTH*2-1+0:0] tmp00_33_7;
	wire [WIDTH*2-1+0:0] tmp00_33_8;
	wire [WIDTH*2-1+0:0] tmp00_33_9;
	wire [WIDTH*2-1+0:0] tmp00_33_10;
	wire [WIDTH*2-1+0:0] tmp00_33_11;
	wire [WIDTH*2-1+0:0] tmp00_33_12;
	wire [WIDTH*2-1+0:0] tmp00_33_13;
	wire [WIDTH*2-1+0:0] tmp00_33_14;
	wire [WIDTH*2-1+0:0] tmp00_33_15;
	wire [WIDTH*2-1+0:0] tmp00_33_16;
	wire [WIDTH*2-1+0:0] tmp00_33_17;
	wire [WIDTH*2-1+0:0] tmp00_33_18;
	wire [WIDTH*2-1+0:0] tmp00_33_19;
	wire [WIDTH*2-1+0:0] tmp00_33_20;
	wire [WIDTH*2-1+0:0] tmp00_33_21;
	wire [WIDTH*2-1+0:0] tmp00_33_22;
	wire [WIDTH*2-1+0:0] tmp00_33_23;
	wire [WIDTH*2-1+0:0] tmp00_33_24;
	wire [WIDTH*2-1+0:0] tmp00_33_25;
	wire [WIDTH*2-1+0:0] tmp00_33_26;
	wire [WIDTH*2-1+0:0] tmp00_33_27;
	wire [WIDTH*2-1+0:0] tmp00_33_28;
	wire [WIDTH*2-1+0:0] tmp00_33_29;
	wire [WIDTH*2-1+0:0] tmp00_33_30;
	wire [WIDTH*2-1+0:0] tmp00_33_31;
	wire [WIDTH*2-1+0:0] tmp00_33_32;
	wire [WIDTH*2-1+0:0] tmp00_33_33;
	wire [WIDTH*2-1+0:0] tmp00_33_34;
	wire [WIDTH*2-1+0:0] tmp00_33_35;
	wire [WIDTH*2-1+0:0] tmp00_33_36;
	wire [WIDTH*2-1+0:0] tmp00_33_37;
	wire [WIDTH*2-1+0:0] tmp00_33_38;
	wire [WIDTH*2-1+0:0] tmp00_33_39;
	wire [WIDTH*2-1+0:0] tmp00_33_40;
	wire [WIDTH*2-1+0:0] tmp00_33_41;
	wire [WIDTH*2-1+0:0] tmp00_33_42;
	wire [WIDTH*2-1+0:0] tmp00_33_43;
	wire [WIDTH*2-1+0:0] tmp00_33_44;
	wire [WIDTH*2-1+0:0] tmp00_33_45;
	wire [WIDTH*2-1+0:0] tmp00_33_46;
	wire [WIDTH*2-1+0:0] tmp00_33_47;
	wire [WIDTH*2-1+0:0] tmp00_33_48;
	wire [WIDTH*2-1+0:0] tmp00_33_49;
	wire [WIDTH*2-1+0:0] tmp00_33_50;
	wire [WIDTH*2-1+0:0] tmp00_33_51;
	wire [WIDTH*2-1+0:0] tmp00_33_52;
	wire [WIDTH*2-1+0:0] tmp00_33_53;
	wire [WIDTH*2-1+0:0] tmp00_33_54;
	wire [WIDTH*2-1+0:0] tmp00_33_55;
	wire [WIDTH*2-1+0:0] tmp00_33_56;
	wire [WIDTH*2-1+0:0] tmp00_33_57;
	wire [WIDTH*2-1+0:0] tmp00_33_58;
	wire [WIDTH*2-1+0:0] tmp00_33_59;
	wire [WIDTH*2-1+0:0] tmp00_33_60;
	wire [WIDTH*2-1+0:0] tmp00_33_61;
	wire [WIDTH*2-1+0:0] tmp00_33_62;
	wire [WIDTH*2-1+0:0] tmp00_33_63;
	wire [WIDTH*2-1+0:0] tmp00_33_64;
	wire [WIDTH*2-1+0:0] tmp00_33_65;
	wire [WIDTH*2-1+0:0] tmp00_33_66;
	wire [WIDTH*2-1+0:0] tmp00_33_67;
	wire [WIDTH*2-1+0:0] tmp00_33_68;
	wire [WIDTH*2-1+0:0] tmp00_33_69;
	wire [WIDTH*2-1+0:0] tmp00_33_70;
	wire [WIDTH*2-1+0:0] tmp00_33_71;
	wire [WIDTH*2-1+0:0] tmp00_33_72;
	wire [WIDTH*2-1+0:0] tmp00_33_73;
	wire [WIDTH*2-1+0:0] tmp00_33_74;
	wire [WIDTH*2-1+0:0] tmp00_33_75;
	wire [WIDTH*2-1+0:0] tmp00_33_76;
	wire [WIDTH*2-1+0:0] tmp00_33_77;
	wire [WIDTH*2-1+0:0] tmp00_33_78;
	wire [WIDTH*2-1+0:0] tmp00_33_79;
	wire [WIDTH*2-1+0:0] tmp00_33_80;
	wire [WIDTH*2-1+0:0] tmp00_33_81;
	wire [WIDTH*2-1+0:0] tmp00_33_82;
	wire [WIDTH*2-1+0:0] tmp00_33_83;
	wire [WIDTH*2-1+0:0] tmp00_34_0;
	wire [WIDTH*2-1+0:0] tmp00_34_1;
	wire [WIDTH*2-1+0:0] tmp00_34_2;
	wire [WIDTH*2-1+0:0] tmp00_34_3;
	wire [WIDTH*2-1+0:0] tmp00_34_4;
	wire [WIDTH*2-1+0:0] tmp00_34_5;
	wire [WIDTH*2-1+0:0] tmp00_34_6;
	wire [WIDTH*2-1+0:0] tmp00_34_7;
	wire [WIDTH*2-1+0:0] tmp00_34_8;
	wire [WIDTH*2-1+0:0] tmp00_34_9;
	wire [WIDTH*2-1+0:0] tmp00_34_10;
	wire [WIDTH*2-1+0:0] tmp00_34_11;
	wire [WIDTH*2-1+0:0] tmp00_34_12;
	wire [WIDTH*2-1+0:0] tmp00_34_13;
	wire [WIDTH*2-1+0:0] tmp00_34_14;
	wire [WIDTH*2-1+0:0] tmp00_34_15;
	wire [WIDTH*2-1+0:0] tmp00_34_16;
	wire [WIDTH*2-1+0:0] tmp00_34_17;
	wire [WIDTH*2-1+0:0] tmp00_34_18;
	wire [WIDTH*2-1+0:0] tmp00_34_19;
	wire [WIDTH*2-1+0:0] tmp00_34_20;
	wire [WIDTH*2-1+0:0] tmp00_34_21;
	wire [WIDTH*2-1+0:0] tmp00_34_22;
	wire [WIDTH*2-1+0:0] tmp00_34_23;
	wire [WIDTH*2-1+0:0] tmp00_34_24;
	wire [WIDTH*2-1+0:0] tmp00_34_25;
	wire [WIDTH*2-1+0:0] tmp00_34_26;
	wire [WIDTH*2-1+0:0] tmp00_34_27;
	wire [WIDTH*2-1+0:0] tmp00_34_28;
	wire [WIDTH*2-1+0:0] tmp00_34_29;
	wire [WIDTH*2-1+0:0] tmp00_34_30;
	wire [WIDTH*2-1+0:0] tmp00_34_31;
	wire [WIDTH*2-1+0:0] tmp00_34_32;
	wire [WIDTH*2-1+0:0] tmp00_34_33;
	wire [WIDTH*2-1+0:0] tmp00_34_34;
	wire [WIDTH*2-1+0:0] tmp00_34_35;
	wire [WIDTH*2-1+0:0] tmp00_34_36;
	wire [WIDTH*2-1+0:0] tmp00_34_37;
	wire [WIDTH*2-1+0:0] tmp00_34_38;
	wire [WIDTH*2-1+0:0] tmp00_34_39;
	wire [WIDTH*2-1+0:0] tmp00_34_40;
	wire [WIDTH*2-1+0:0] tmp00_34_41;
	wire [WIDTH*2-1+0:0] tmp00_34_42;
	wire [WIDTH*2-1+0:0] tmp00_34_43;
	wire [WIDTH*2-1+0:0] tmp00_34_44;
	wire [WIDTH*2-1+0:0] tmp00_34_45;
	wire [WIDTH*2-1+0:0] tmp00_34_46;
	wire [WIDTH*2-1+0:0] tmp00_34_47;
	wire [WIDTH*2-1+0:0] tmp00_34_48;
	wire [WIDTH*2-1+0:0] tmp00_34_49;
	wire [WIDTH*2-1+0:0] tmp00_34_50;
	wire [WIDTH*2-1+0:0] tmp00_34_51;
	wire [WIDTH*2-1+0:0] tmp00_34_52;
	wire [WIDTH*2-1+0:0] tmp00_34_53;
	wire [WIDTH*2-1+0:0] tmp00_34_54;
	wire [WIDTH*2-1+0:0] tmp00_34_55;
	wire [WIDTH*2-1+0:0] tmp00_34_56;
	wire [WIDTH*2-1+0:0] tmp00_34_57;
	wire [WIDTH*2-1+0:0] tmp00_34_58;
	wire [WIDTH*2-1+0:0] tmp00_34_59;
	wire [WIDTH*2-1+0:0] tmp00_34_60;
	wire [WIDTH*2-1+0:0] tmp00_34_61;
	wire [WIDTH*2-1+0:0] tmp00_34_62;
	wire [WIDTH*2-1+0:0] tmp00_34_63;
	wire [WIDTH*2-1+0:0] tmp00_34_64;
	wire [WIDTH*2-1+0:0] tmp00_34_65;
	wire [WIDTH*2-1+0:0] tmp00_34_66;
	wire [WIDTH*2-1+0:0] tmp00_34_67;
	wire [WIDTH*2-1+0:0] tmp00_34_68;
	wire [WIDTH*2-1+0:0] tmp00_34_69;
	wire [WIDTH*2-1+0:0] tmp00_34_70;
	wire [WIDTH*2-1+0:0] tmp00_34_71;
	wire [WIDTH*2-1+0:0] tmp00_34_72;
	wire [WIDTH*2-1+0:0] tmp00_34_73;
	wire [WIDTH*2-1+0:0] tmp00_34_74;
	wire [WIDTH*2-1+0:0] tmp00_34_75;
	wire [WIDTH*2-1+0:0] tmp00_34_76;
	wire [WIDTH*2-1+0:0] tmp00_34_77;
	wire [WIDTH*2-1+0:0] tmp00_34_78;
	wire [WIDTH*2-1+0:0] tmp00_34_79;
	wire [WIDTH*2-1+0:0] tmp00_34_80;
	wire [WIDTH*2-1+0:0] tmp00_34_81;
	wire [WIDTH*2-1+0:0] tmp00_34_82;
	wire [WIDTH*2-1+0:0] tmp00_34_83;
	wire [WIDTH*2-1+0:0] tmp00_35_0;
	wire [WIDTH*2-1+0:0] tmp00_35_1;
	wire [WIDTH*2-1+0:0] tmp00_35_2;
	wire [WIDTH*2-1+0:0] tmp00_35_3;
	wire [WIDTH*2-1+0:0] tmp00_35_4;
	wire [WIDTH*2-1+0:0] tmp00_35_5;
	wire [WIDTH*2-1+0:0] tmp00_35_6;
	wire [WIDTH*2-1+0:0] tmp00_35_7;
	wire [WIDTH*2-1+0:0] tmp00_35_8;
	wire [WIDTH*2-1+0:0] tmp00_35_9;
	wire [WIDTH*2-1+0:0] tmp00_35_10;
	wire [WIDTH*2-1+0:0] tmp00_35_11;
	wire [WIDTH*2-1+0:0] tmp00_35_12;
	wire [WIDTH*2-1+0:0] tmp00_35_13;
	wire [WIDTH*2-1+0:0] tmp00_35_14;
	wire [WIDTH*2-1+0:0] tmp00_35_15;
	wire [WIDTH*2-1+0:0] tmp00_35_16;
	wire [WIDTH*2-1+0:0] tmp00_35_17;
	wire [WIDTH*2-1+0:0] tmp00_35_18;
	wire [WIDTH*2-1+0:0] tmp00_35_19;
	wire [WIDTH*2-1+0:0] tmp00_35_20;
	wire [WIDTH*2-1+0:0] tmp00_35_21;
	wire [WIDTH*2-1+0:0] tmp00_35_22;
	wire [WIDTH*2-1+0:0] tmp00_35_23;
	wire [WIDTH*2-1+0:0] tmp00_35_24;
	wire [WIDTH*2-1+0:0] tmp00_35_25;
	wire [WIDTH*2-1+0:0] tmp00_35_26;
	wire [WIDTH*2-1+0:0] tmp00_35_27;
	wire [WIDTH*2-1+0:0] tmp00_35_28;
	wire [WIDTH*2-1+0:0] tmp00_35_29;
	wire [WIDTH*2-1+0:0] tmp00_35_30;
	wire [WIDTH*2-1+0:0] tmp00_35_31;
	wire [WIDTH*2-1+0:0] tmp00_35_32;
	wire [WIDTH*2-1+0:0] tmp00_35_33;
	wire [WIDTH*2-1+0:0] tmp00_35_34;
	wire [WIDTH*2-1+0:0] tmp00_35_35;
	wire [WIDTH*2-1+0:0] tmp00_35_36;
	wire [WIDTH*2-1+0:0] tmp00_35_37;
	wire [WIDTH*2-1+0:0] tmp00_35_38;
	wire [WIDTH*2-1+0:0] tmp00_35_39;
	wire [WIDTH*2-1+0:0] tmp00_35_40;
	wire [WIDTH*2-1+0:0] tmp00_35_41;
	wire [WIDTH*2-1+0:0] tmp00_35_42;
	wire [WIDTH*2-1+0:0] tmp00_35_43;
	wire [WIDTH*2-1+0:0] tmp00_35_44;
	wire [WIDTH*2-1+0:0] tmp00_35_45;
	wire [WIDTH*2-1+0:0] tmp00_35_46;
	wire [WIDTH*2-1+0:0] tmp00_35_47;
	wire [WIDTH*2-1+0:0] tmp00_35_48;
	wire [WIDTH*2-1+0:0] tmp00_35_49;
	wire [WIDTH*2-1+0:0] tmp00_35_50;
	wire [WIDTH*2-1+0:0] tmp00_35_51;
	wire [WIDTH*2-1+0:0] tmp00_35_52;
	wire [WIDTH*2-1+0:0] tmp00_35_53;
	wire [WIDTH*2-1+0:0] tmp00_35_54;
	wire [WIDTH*2-1+0:0] tmp00_35_55;
	wire [WIDTH*2-1+0:0] tmp00_35_56;
	wire [WIDTH*2-1+0:0] tmp00_35_57;
	wire [WIDTH*2-1+0:0] tmp00_35_58;
	wire [WIDTH*2-1+0:0] tmp00_35_59;
	wire [WIDTH*2-1+0:0] tmp00_35_60;
	wire [WIDTH*2-1+0:0] tmp00_35_61;
	wire [WIDTH*2-1+0:0] tmp00_35_62;
	wire [WIDTH*2-1+0:0] tmp00_35_63;
	wire [WIDTH*2-1+0:0] tmp00_35_64;
	wire [WIDTH*2-1+0:0] tmp00_35_65;
	wire [WIDTH*2-1+0:0] tmp00_35_66;
	wire [WIDTH*2-1+0:0] tmp00_35_67;
	wire [WIDTH*2-1+0:0] tmp00_35_68;
	wire [WIDTH*2-1+0:0] tmp00_35_69;
	wire [WIDTH*2-1+0:0] tmp00_35_70;
	wire [WIDTH*2-1+0:0] tmp00_35_71;
	wire [WIDTH*2-1+0:0] tmp00_35_72;
	wire [WIDTH*2-1+0:0] tmp00_35_73;
	wire [WIDTH*2-1+0:0] tmp00_35_74;
	wire [WIDTH*2-1+0:0] tmp00_35_75;
	wire [WIDTH*2-1+0:0] tmp00_35_76;
	wire [WIDTH*2-1+0:0] tmp00_35_77;
	wire [WIDTH*2-1+0:0] tmp00_35_78;
	wire [WIDTH*2-1+0:0] tmp00_35_79;
	wire [WIDTH*2-1+0:0] tmp00_35_80;
	wire [WIDTH*2-1+0:0] tmp00_35_81;
	wire [WIDTH*2-1+0:0] tmp00_35_82;
	wire [WIDTH*2-1+0:0] tmp00_35_83;
	wire [WIDTH*2-1+0:0] tmp00_36_0;
	wire [WIDTH*2-1+0:0] tmp00_36_1;
	wire [WIDTH*2-1+0:0] tmp00_36_2;
	wire [WIDTH*2-1+0:0] tmp00_36_3;
	wire [WIDTH*2-1+0:0] tmp00_36_4;
	wire [WIDTH*2-1+0:0] tmp00_36_5;
	wire [WIDTH*2-1+0:0] tmp00_36_6;
	wire [WIDTH*2-1+0:0] tmp00_36_7;
	wire [WIDTH*2-1+0:0] tmp00_36_8;
	wire [WIDTH*2-1+0:0] tmp00_36_9;
	wire [WIDTH*2-1+0:0] tmp00_36_10;
	wire [WIDTH*2-1+0:0] tmp00_36_11;
	wire [WIDTH*2-1+0:0] tmp00_36_12;
	wire [WIDTH*2-1+0:0] tmp00_36_13;
	wire [WIDTH*2-1+0:0] tmp00_36_14;
	wire [WIDTH*2-1+0:0] tmp00_36_15;
	wire [WIDTH*2-1+0:0] tmp00_36_16;
	wire [WIDTH*2-1+0:0] tmp00_36_17;
	wire [WIDTH*2-1+0:0] tmp00_36_18;
	wire [WIDTH*2-1+0:0] tmp00_36_19;
	wire [WIDTH*2-1+0:0] tmp00_36_20;
	wire [WIDTH*2-1+0:0] tmp00_36_21;
	wire [WIDTH*2-1+0:0] tmp00_36_22;
	wire [WIDTH*2-1+0:0] tmp00_36_23;
	wire [WIDTH*2-1+0:0] tmp00_36_24;
	wire [WIDTH*2-1+0:0] tmp00_36_25;
	wire [WIDTH*2-1+0:0] tmp00_36_26;
	wire [WIDTH*2-1+0:0] tmp00_36_27;
	wire [WIDTH*2-1+0:0] tmp00_36_28;
	wire [WIDTH*2-1+0:0] tmp00_36_29;
	wire [WIDTH*2-1+0:0] tmp00_36_30;
	wire [WIDTH*2-1+0:0] tmp00_36_31;
	wire [WIDTH*2-1+0:0] tmp00_36_32;
	wire [WIDTH*2-1+0:0] tmp00_36_33;
	wire [WIDTH*2-1+0:0] tmp00_36_34;
	wire [WIDTH*2-1+0:0] tmp00_36_35;
	wire [WIDTH*2-1+0:0] tmp00_36_36;
	wire [WIDTH*2-1+0:0] tmp00_36_37;
	wire [WIDTH*2-1+0:0] tmp00_36_38;
	wire [WIDTH*2-1+0:0] tmp00_36_39;
	wire [WIDTH*2-1+0:0] tmp00_36_40;
	wire [WIDTH*2-1+0:0] tmp00_36_41;
	wire [WIDTH*2-1+0:0] tmp00_36_42;
	wire [WIDTH*2-1+0:0] tmp00_36_43;
	wire [WIDTH*2-1+0:0] tmp00_36_44;
	wire [WIDTH*2-1+0:0] tmp00_36_45;
	wire [WIDTH*2-1+0:0] tmp00_36_46;
	wire [WIDTH*2-1+0:0] tmp00_36_47;
	wire [WIDTH*2-1+0:0] tmp00_36_48;
	wire [WIDTH*2-1+0:0] tmp00_36_49;
	wire [WIDTH*2-1+0:0] tmp00_36_50;
	wire [WIDTH*2-1+0:0] tmp00_36_51;
	wire [WIDTH*2-1+0:0] tmp00_36_52;
	wire [WIDTH*2-1+0:0] tmp00_36_53;
	wire [WIDTH*2-1+0:0] tmp00_36_54;
	wire [WIDTH*2-1+0:0] tmp00_36_55;
	wire [WIDTH*2-1+0:0] tmp00_36_56;
	wire [WIDTH*2-1+0:0] tmp00_36_57;
	wire [WIDTH*2-1+0:0] tmp00_36_58;
	wire [WIDTH*2-1+0:0] tmp00_36_59;
	wire [WIDTH*2-1+0:0] tmp00_36_60;
	wire [WIDTH*2-1+0:0] tmp00_36_61;
	wire [WIDTH*2-1+0:0] tmp00_36_62;
	wire [WIDTH*2-1+0:0] tmp00_36_63;
	wire [WIDTH*2-1+0:0] tmp00_36_64;
	wire [WIDTH*2-1+0:0] tmp00_36_65;
	wire [WIDTH*2-1+0:0] tmp00_36_66;
	wire [WIDTH*2-1+0:0] tmp00_36_67;
	wire [WIDTH*2-1+0:0] tmp00_36_68;
	wire [WIDTH*2-1+0:0] tmp00_36_69;
	wire [WIDTH*2-1+0:0] tmp00_36_70;
	wire [WIDTH*2-1+0:0] tmp00_36_71;
	wire [WIDTH*2-1+0:0] tmp00_36_72;
	wire [WIDTH*2-1+0:0] tmp00_36_73;
	wire [WIDTH*2-1+0:0] tmp00_36_74;
	wire [WIDTH*2-1+0:0] tmp00_36_75;
	wire [WIDTH*2-1+0:0] tmp00_36_76;
	wire [WIDTH*2-1+0:0] tmp00_36_77;
	wire [WIDTH*2-1+0:0] tmp00_36_78;
	wire [WIDTH*2-1+0:0] tmp00_36_79;
	wire [WIDTH*2-1+0:0] tmp00_36_80;
	wire [WIDTH*2-1+0:0] tmp00_36_81;
	wire [WIDTH*2-1+0:0] tmp00_36_82;
	wire [WIDTH*2-1+0:0] tmp00_36_83;
	wire [WIDTH*2-1+0:0] tmp00_37_0;
	wire [WIDTH*2-1+0:0] tmp00_37_1;
	wire [WIDTH*2-1+0:0] tmp00_37_2;
	wire [WIDTH*2-1+0:0] tmp00_37_3;
	wire [WIDTH*2-1+0:0] tmp00_37_4;
	wire [WIDTH*2-1+0:0] tmp00_37_5;
	wire [WIDTH*2-1+0:0] tmp00_37_6;
	wire [WIDTH*2-1+0:0] tmp00_37_7;
	wire [WIDTH*2-1+0:0] tmp00_37_8;
	wire [WIDTH*2-1+0:0] tmp00_37_9;
	wire [WIDTH*2-1+0:0] tmp00_37_10;
	wire [WIDTH*2-1+0:0] tmp00_37_11;
	wire [WIDTH*2-1+0:0] tmp00_37_12;
	wire [WIDTH*2-1+0:0] tmp00_37_13;
	wire [WIDTH*2-1+0:0] tmp00_37_14;
	wire [WIDTH*2-1+0:0] tmp00_37_15;
	wire [WIDTH*2-1+0:0] tmp00_37_16;
	wire [WIDTH*2-1+0:0] tmp00_37_17;
	wire [WIDTH*2-1+0:0] tmp00_37_18;
	wire [WIDTH*2-1+0:0] tmp00_37_19;
	wire [WIDTH*2-1+0:0] tmp00_37_20;
	wire [WIDTH*2-1+0:0] tmp00_37_21;
	wire [WIDTH*2-1+0:0] tmp00_37_22;
	wire [WIDTH*2-1+0:0] tmp00_37_23;
	wire [WIDTH*2-1+0:0] tmp00_37_24;
	wire [WIDTH*2-1+0:0] tmp00_37_25;
	wire [WIDTH*2-1+0:0] tmp00_37_26;
	wire [WIDTH*2-1+0:0] tmp00_37_27;
	wire [WIDTH*2-1+0:0] tmp00_37_28;
	wire [WIDTH*2-1+0:0] tmp00_37_29;
	wire [WIDTH*2-1+0:0] tmp00_37_30;
	wire [WIDTH*2-1+0:0] tmp00_37_31;
	wire [WIDTH*2-1+0:0] tmp00_37_32;
	wire [WIDTH*2-1+0:0] tmp00_37_33;
	wire [WIDTH*2-1+0:0] tmp00_37_34;
	wire [WIDTH*2-1+0:0] tmp00_37_35;
	wire [WIDTH*2-1+0:0] tmp00_37_36;
	wire [WIDTH*2-1+0:0] tmp00_37_37;
	wire [WIDTH*2-1+0:0] tmp00_37_38;
	wire [WIDTH*2-1+0:0] tmp00_37_39;
	wire [WIDTH*2-1+0:0] tmp00_37_40;
	wire [WIDTH*2-1+0:0] tmp00_37_41;
	wire [WIDTH*2-1+0:0] tmp00_37_42;
	wire [WIDTH*2-1+0:0] tmp00_37_43;
	wire [WIDTH*2-1+0:0] tmp00_37_44;
	wire [WIDTH*2-1+0:0] tmp00_37_45;
	wire [WIDTH*2-1+0:0] tmp00_37_46;
	wire [WIDTH*2-1+0:0] tmp00_37_47;
	wire [WIDTH*2-1+0:0] tmp00_37_48;
	wire [WIDTH*2-1+0:0] tmp00_37_49;
	wire [WIDTH*2-1+0:0] tmp00_37_50;
	wire [WIDTH*2-1+0:0] tmp00_37_51;
	wire [WIDTH*2-1+0:0] tmp00_37_52;
	wire [WIDTH*2-1+0:0] tmp00_37_53;
	wire [WIDTH*2-1+0:0] tmp00_37_54;
	wire [WIDTH*2-1+0:0] tmp00_37_55;
	wire [WIDTH*2-1+0:0] tmp00_37_56;
	wire [WIDTH*2-1+0:0] tmp00_37_57;
	wire [WIDTH*2-1+0:0] tmp00_37_58;
	wire [WIDTH*2-1+0:0] tmp00_37_59;
	wire [WIDTH*2-1+0:0] tmp00_37_60;
	wire [WIDTH*2-1+0:0] tmp00_37_61;
	wire [WIDTH*2-1+0:0] tmp00_37_62;
	wire [WIDTH*2-1+0:0] tmp00_37_63;
	wire [WIDTH*2-1+0:0] tmp00_37_64;
	wire [WIDTH*2-1+0:0] tmp00_37_65;
	wire [WIDTH*2-1+0:0] tmp00_37_66;
	wire [WIDTH*2-1+0:0] tmp00_37_67;
	wire [WIDTH*2-1+0:0] tmp00_37_68;
	wire [WIDTH*2-1+0:0] tmp00_37_69;
	wire [WIDTH*2-1+0:0] tmp00_37_70;
	wire [WIDTH*2-1+0:0] tmp00_37_71;
	wire [WIDTH*2-1+0:0] tmp00_37_72;
	wire [WIDTH*2-1+0:0] tmp00_37_73;
	wire [WIDTH*2-1+0:0] tmp00_37_74;
	wire [WIDTH*2-1+0:0] tmp00_37_75;
	wire [WIDTH*2-1+0:0] tmp00_37_76;
	wire [WIDTH*2-1+0:0] tmp00_37_77;
	wire [WIDTH*2-1+0:0] tmp00_37_78;
	wire [WIDTH*2-1+0:0] tmp00_37_79;
	wire [WIDTH*2-1+0:0] tmp00_37_80;
	wire [WIDTH*2-1+0:0] tmp00_37_81;
	wire [WIDTH*2-1+0:0] tmp00_37_82;
	wire [WIDTH*2-1+0:0] tmp00_37_83;
	wire [WIDTH*2-1+0:0] tmp00_38_0;
	wire [WIDTH*2-1+0:0] tmp00_38_1;
	wire [WIDTH*2-1+0:0] tmp00_38_2;
	wire [WIDTH*2-1+0:0] tmp00_38_3;
	wire [WIDTH*2-1+0:0] tmp00_38_4;
	wire [WIDTH*2-1+0:0] tmp00_38_5;
	wire [WIDTH*2-1+0:0] tmp00_38_6;
	wire [WIDTH*2-1+0:0] tmp00_38_7;
	wire [WIDTH*2-1+0:0] tmp00_38_8;
	wire [WIDTH*2-1+0:0] tmp00_38_9;
	wire [WIDTH*2-1+0:0] tmp00_38_10;
	wire [WIDTH*2-1+0:0] tmp00_38_11;
	wire [WIDTH*2-1+0:0] tmp00_38_12;
	wire [WIDTH*2-1+0:0] tmp00_38_13;
	wire [WIDTH*2-1+0:0] tmp00_38_14;
	wire [WIDTH*2-1+0:0] tmp00_38_15;
	wire [WIDTH*2-1+0:0] tmp00_38_16;
	wire [WIDTH*2-1+0:0] tmp00_38_17;
	wire [WIDTH*2-1+0:0] tmp00_38_18;
	wire [WIDTH*2-1+0:0] tmp00_38_19;
	wire [WIDTH*2-1+0:0] tmp00_38_20;
	wire [WIDTH*2-1+0:0] tmp00_38_21;
	wire [WIDTH*2-1+0:0] tmp00_38_22;
	wire [WIDTH*2-1+0:0] tmp00_38_23;
	wire [WIDTH*2-1+0:0] tmp00_38_24;
	wire [WIDTH*2-1+0:0] tmp00_38_25;
	wire [WIDTH*2-1+0:0] tmp00_38_26;
	wire [WIDTH*2-1+0:0] tmp00_38_27;
	wire [WIDTH*2-1+0:0] tmp00_38_28;
	wire [WIDTH*2-1+0:0] tmp00_38_29;
	wire [WIDTH*2-1+0:0] tmp00_38_30;
	wire [WIDTH*2-1+0:0] tmp00_38_31;
	wire [WIDTH*2-1+0:0] tmp00_38_32;
	wire [WIDTH*2-1+0:0] tmp00_38_33;
	wire [WIDTH*2-1+0:0] tmp00_38_34;
	wire [WIDTH*2-1+0:0] tmp00_38_35;
	wire [WIDTH*2-1+0:0] tmp00_38_36;
	wire [WIDTH*2-1+0:0] tmp00_38_37;
	wire [WIDTH*2-1+0:0] tmp00_38_38;
	wire [WIDTH*2-1+0:0] tmp00_38_39;
	wire [WIDTH*2-1+0:0] tmp00_38_40;
	wire [WIDTH*2-1+0:0] tmp00_38_41;
	wire [WIDTH*2-1+0:0] tmp00_38_42;
	wire [WIDTH*2-1+0:0] tmp00_38_43;
	wire [WIDTH*2-1+0:0] tmp00_38_44;
	wire [WIDTH*2-1+0:0] tmp00_38_45;
	wire [WIDTH*2-1+0:0] tmp00_38_46;
	wire [WIDTH*2-1+0:0] tmp00_38_47;
	wire [WIDTH*2-1+0:0] tmp00_38_48;
	wire [WIDTH*2-1+0:0] tmp00_38_49;
	wire [WIDTH*2-1+0:0] tmp00_38_50;
	wire [WIDTH*2-1+0:0] tmp00_38_51;
	wire [WIDTH*2-1+0:0] tmp00_38_52;
	wire [WIDTH*2-1+0:0] tmp00_38_53;
	wire [WIDTH*2-1+0:0] tmp00_38_54;
	wire [WIDTH*2-1+0:0] tmp00_38_55;
	wire [WIDTH*2-1+0:0] tmp00_38_56;
	wire [WIDTH*2-1+0:0] tmp00_38_57;
	wire [WIDTH*2-1+0:0] tmp00_38_58;
	wire [WIDTH*2-1+0:0] tmp00_38_59;
	wire [WIDTH*2-1+0:0] tmp00_38_60;
	wire [WIDTH*2-1+0:0] tmp00_38_61;
	wire [WIDTH*2-1+0:0] tmp00_38_62;
	wire [WIDTH*2-1+0:0] tmp00_38_63;
	wire [WIDTH*2-1+0:0] tmp00_38_64;
	wire [WIDTH*2-1+0:0] tmp00_38_65;
	wire [WIDTH*2-1+0:0] tmp00_38_66;
	wire [WIDTH*2-1+0:0] tmp00_38_67;
	wire [WIDTH*2-1+0:0] tmp00_38_68;
	wire [WIDTH*2-1+0:0] tmp00_38_69;
	wire [WIDTH*2-1+0:0] tmp00_38_70;
	wire [WIDTH*2-1+0:0] tmp00_38_71;
	wire [WIDTH*2-1+0:0] tmp00_38_72;
	wire [WIDTH*2-1+0:0] tmp00_38_73;
	wire [WIDTH*2-1+0:0] tmp00_38_74;
	wire [WIDTH*2-1+0:0] tmp00_38_75;
	wire [WIDTH*2-1+0:0] tmp00_38_76;
	wire [WIDTH*2-1+0:0] tmp00_38_77;
	wire [WIDTH*2-1+0:0] tmp00_38_78;
	wire [WIDTH*2-1+0:0] tmp00_38_79;
	wire [WIDTH*2-1+0:0] tmp00_38_80;
	wire [WIDTH*2-1+0:0] tmp00_38_81;
	wire [WIDTH*2-1+0:0] tmp00_38_82;
	wire [WIDTH*2-1+0:0] tmp00_38_83;
	wire [WIDTH*2-1+0:0] tmp00_39_0;
	wire [WIDTH*2-1+0:0] tmp00_39_1;
	wire [WIDTH*2-1+0:0] tmp00_39_2;
	wire [WIDTH*2-1+0:0] tmp00_39_3;
	wire [WIDTH*2-1+0:0] tmp00_39_4;
	wire [WIDTH*2-1+0:0] tmp00_39_5;
	wire [WIDTH*2-1+0:0] tmp00_39_6;
	wire [WIDTH*2-1+0:0] tmp00_39_7;
	wire [WIDTH*2-1+0:0] tmp00_39_8;
	wire [WIDTH*2-1+0:0] tmp00_39_9;
	wire [WIDTH*2-1+0:0] tmp00_39_10;
	wire [WIDTH*2-1+0:0] tmp00_39_11;
	wire [WIDTH*2-1+0:0] tmp00_39_12;
	wire [WIDTH*2-1+0:0] tmp00_39_13;
	wire [WIDTH*2-1+0:0] tmp00_39_14;
	wire [WIDTH*2-1+0:0] tmp00_39_15;
	wire [WIDTH*2-1+0:0] tmp00_39_16;
	wire [WIDTH*2-1+0:0] tmp00_39_17;
	wire [WIDTH*2-1+0:0] tmp00_39_18;
	wire [WIDTH*2-1+0:0] tmp00_39_19;
	wire [WIDTH*2-1+0:0] tmp00_39_20;
	wire [WIDTH*2-1+0:0] tmp00_39_21;
	wire [WIDTH*2-1+0:0] tmp00_39_22;
	wire [WIDTH*2-1+0:0] tmp00_39_23;
	wire [WIDTH*2-1+0:0] tmp00_39_24;
	wire [WIDTH*2-1+0:0] tmp00_39_25;
	wire [WIDTH*2-1+0:0] tmp00_39_26;
	wire [WIDTH*2-1+0:0] tmp00_39_27;
	wire [WIDTH*2-1+0:0] tmp00_39_28;
	wire [WIDTH*2-1+0:0] tmp00_39_29;
	wire [WIDTH*2-1+0:0] tmp00_39_30;
	wire [WIDTH*2-1+0:0] tmp00_39_31;
	wire [WIDTH*2-1+0:0] tmp00_39_32;
	wire [WIDTH*2-1+0:0] tmp00_39_33;
	wire [WIDTH*2-1+0:0] tmp00_39_34;
	wire [WIDTH*2-1+0:0] tmp00_39_35;
	wire [WIDTH*2-1+0:0] tmp00_39_36;
	wire [WIDTH*2-1+0:0] tmp00_39_37;
	wire [WIDTH*2-1+0:0] tmp00_39_38;
	wire [WIDTH*2-1+0:0] tmp00_39_39;
	wire [WIDTH*2-1+0:0] tmp00_39_40;
	wire [WIDTH*2-1+0:0] tmp00_39_41;
	wire [WIDTH*2-1+0:0] tmp00_39_42;
	wire [WIDTH*2-1+0:0] tmp00_39_43;
	wire [WIDTH*2-1+0:0] tmp00_39_44;
	wire [WIDTH*2-1+0:0] tmp00_39_45;
	wire [WIDTH*2-1+0:0] tmp00_39_46;
	wire [WIDTH*2-1+0:0] tmp00_39_47;
	wire [WIDTH*2-1+0:0] tmp00_39_48;
	wire [WIDTH*2-1+0:0] tmp00_39_49;
	wire [WIDTH*2-1+0:0] tmp00_39_50;
	wire [WIDTH*2-1+0:0] tmp00_39_51;
	wire [WIDTH*2-1+0:0] tmp00_39_52;
	wire [WIDTH*2-1+0:0] tmp00_39_53;
	wire [WIDTH*2-1+0:0] tmp00_39_54;
	wire [WIDTH*2-1+0:0] tmp00_39_55;
	wire [WIDTH*2-1+0:0] tmp00_39_56;
	wire [WIDTH*2-1+0:0] tmp00_39_57;
	wire [WIDTH*2-1+0:0] tmp00_39_58;
	wire [WIDTH*2-1+0:0] tmp00_39_59;
	wire [WIDTH*2-1+0:0] tmp00_39_60;
	wire [WIDTH*2-1+0:0] tmp00_39_61;
	wire [WIDTH*2-1+0:0] tmp00_39_62;
	wire [WIDTH*2-1+0:0] tmp00_39_63;
	wire [WIDTH*2-1+0:0] tmp00_39_64;
	wire [WIDTH*2-1+0:0] tmp00_39_65;
	wire [WIDTH*2-1+0:0] tmp00_39_66;
	wire [WIDTH*2-1+0:0] tmp00_39_67;
	wire [WIDTH*2-1+0:0] tmp00_39_68;
	wire [WIDTH*2-1+0:0] tmp00_39_69;
	wire [WIDTH*2-1+0:0] tmp00_39_70;
	wire [WIDTH*2-1+0:0] tmp00_39_71;
	wire [WIDTH*2-1+0:0] tmp00_39_72;
	wire [WIDTH*2-1+0:0] tmp00_39_73;
	wire [WIDTH*2-1+0:0] tmp00_39_74;
	wire [WIDTH*2-1+0:0] tmp00_39_75;
	wire [WIDTH*2-1+0:0] tmp00_39_76;
	wire [WIDTH*2-1+0:0] tmp00_39_77;
	wire [WIDTH*2-1+0:0] tmp00_39_78;
	wire [WIDTH*2-1+0:0] tmp00_39_79;
	wire [WIDTH*2-1+0:0] tmp00_39_80;
	wire [WIDTH*2-1+0:0] tmp00_39_81;
	wire [WIDTH*2-1+0:0] tmp00_39_82;
	wire [WIDTH*2-1+0:0] tmp00_39_83;
	wire [WIDTH*2-1+0:0] tmp00_40_0;
	wire [WIDTH*2-1+0:0] tmp00_40_1;
	wire [WIDTH*2-1+0:0] tmp00_40_2;
	wire [WIDTH*2-1+0:0] tmp00_40_3;
	wire [WIDTH*2-1+0:0] tmp00_40_4;
	wire [WIDTH*2-1+0:0] tmp00_40_5;
	wire [WIDTH*2-1+0:0] tmp00_40_6;
	wire [WIDTH*2-1+0:0] tmp00_40_7;
	wire [WIDTH*2-1+0:0] tmp00_40_8;
	wire [WIDTH*2-1+0:0] tmp00_40_9;
	wire [WIDTH*2-1+0:0] tmp00_40_10;
	wire [WIDTH*2-1+0:0] tmp00_40_11;
	wire [WIDTH*2-1+0:0] tmp00_40_12;
	wire [WIDTH*2-1+0:0] tmp00_40_13;
	wire [WIDTH*2-1+0:0] tmp00_40_14;
	wire [WIDTH*2-1+0:0] tmp00_40_15;
	wire [WIDTH*2-1+0:0] tmp00_40_16;
	wire [WIDTH*2-1+0:0] tmp00_40_17;
	wire [WIDTH*2-1+0:0] tmp00_40_18;
	wire [WIDTH*2-1+0:0] tmp00_40_19;
	wire [WIDTH*2-1+0:0] tmp00_40_20;
	wire [WIDTH*2-1+0:0] tmp00_40_21;
	wire [WIDTH*2-1+0:0] tmp00_40_22;
	wire [WIDTH*2-1+0:0] tmp00_40_23;
	wire [WIDTH*2-1+0:0] tmp00_40_24;
	wire [WIDTH*2-1+0:0] tmp00_40_25;
	wire [WIDTH*2-1+0:0] tmp00_40_26;
	wire [WIDTH*2-1+0:0] tmp00_40_27;
	wire [WIDTH*2-1+0:0] tmp00_40_28;
	wire [WIDTH*2-1+0:0] tmp00_40_29;
	wire [WIDTH*2-1+0:0] tmp00_40_30;
	wire [WIDTH*2-1+0:0] tmp00_40_31;
	wire [WIDTH*2-1+0:0] tmp00_40_32;
	wire [WIDTH*2-1+0:0] tmp00_40_33;
	wire [WIDTH*2-1+0:0] tmp00_40_34;
	wire [WIDTH*2-1+0:0] tmp00_40_35;
	wire [WIDTH*2-1+0:0] tmp00_40_36;
	wire [WIDTH*2-1+0:0] tmp00_40_37;
	wire [WIDTH*2-1+0:0] tmp00_40_38;
	wire [WIDTH*2-1+0:0] tmp00_40_39;
	wire [WIDTH*2-1+0:0] tmp00_40_40;
	wire [WIDTH*2-1+0:0] tmp00_40_41;
	wire [WIDTH*2-1+0:0] tmp00_40_42;
	wire [WIDTH*2-1+0:0] tmp00_40_43;
	wire [WIDTH*2-1+0:0] tmp00_40_44;
	wire [WIDTH*2-1+0:0] tmp00_40_45;
	wire [WIDTH*2-1+0:0] tmp00_40_46;
	wire [WIDTH*2-1+0:0] tmp00_40_47;
	wire [WIDTH*2-1+0:0] tmp00_40_48;
	wire [WIDTH*2-1+0:0] tmp00_40_49;
	wire [WIDTH*2-1+0:0] tmp00_40_50;
	wire [WIDTH*2-1+0:0] tmp00_40_51;
	wire [WIDTH*2-1+0:0] tmp00_40_52;
	wire [WIDTH*2-1+0:0] tmp00_40_53;
	wire [WIDTH*2-1+0:0] tmp00_40_54;
	wire [WIDTH*2-1+0:0] tmp00_40_55;
	wire [WIDTH*2-1+0:0] tmp00_40_56;
	wire [WIDTH*2-1+0:0] tmp00_40_57;
	wire [WIDTH*2-1+0:0] tmp00_40_58;
	wire [WIDTH*2-1+0:0] tmp00_40_59;
	wire [WIDTH*2-1+0:0] tmp00_40_60;
	wire [WIDTH*2-1+0:0] tmp00_40_61;
	wire [WIDTH*2-1+0:0] tmp00_40_62;
	wire [WIDTH*2-1+0:0] tmp00_40_63;
	wire [WIDTH*2-1+0:0] tmp00_40_64;
	wire [WIDTH*2-1+0:0] tmp00_40_65;
	wire [WIDTH*2-1+0:0] tmp00_40_66;
	wire [WIDTH*2-1+0:0] tmp00_40_67;
	wire [WIDTH*2-1+0:0] tmp00_40_68;
	wire [WIDTH*2-1+0:0] tmp00_40_69;
	wire [WIDTH*2-1+0:0] tmp00_40_70;
	wire [WIDTH*2-1+0:0] tmp00_40_71;
	wire [WIDTH*2-1+0:0] tmp00_40_72;
	wire [WIDTH*2-1+0:0] tmp00_40_73;
	wire [WIDTH*2-1+0:0] tmp00_40_74;
	wire [WIDTH*2-1+0:0] tmp00_40_75;
	wire [WIDTH*2-1+0:0] tmp00_40_76;
	wire [WIDTH*2-1+0:0] tmp00_40_77;
	wire [WIDTH*2-1+0:0] tmp00_40_78;
	wire [WIDTH*2-1+0:0] tmp00_40_79;
	wire [WIDTH*2-1+0:0] tmp00_40_80;
	wire [WIDTH*2-1+0:0] tmp00_40_81;
	wire [WIDTH*2-1+0:0] tmp00_40_82;
	wire [WIDTH*2-1+0:0] tmp00_40_83;
	wire [WIDTH*2-1+0:0] tmp00_41_0;
	wire [WIDTH*2-1+0:0] tmp00_41_1;
	wire [WIDTH*2-1+0:0] tmp00_41_2;
	wire [WIDTH*2-1+0:0] tmp00_41_3;
	wire [WIDTH*2-1+0:0] tmp00_41_4;
	wire [WIDTH*2-1+0:0] tmp00_41_5;
	wire [WIDTH*2-1+0:0] tmp00_41_6;
	wire [WIDTH*2-1+0:0] tmp00_41_7;
	wire [WIDTH*2-1+0:0] tmp00_41_8;
	wire [WIDTH*2-1+0:0] tmp00_41_9;
	wire [WIDTH*2-1+0:0] tmp00_41_10;
	wire [WIDTH*2-1+0:0] tmp00_41_11;
	wire [WIDTH*2-1+0:0] tmp00_41_12;
	wire [WIDTH*2-1+0:0] tmp00_41_13;
	wire [WIDTH*2-1+0:0] tmp00_41_14;
	wire [WIDTH*2-1+0:0] tmp00_41_15;
	wire [WIDTH*2-1+0:0] tmp00_41_16;
	wire [WIDTH*2-1+0:0] tmp00_41_17;
	wire [WIDTH*2-1+0:0] tmp00_41_18;
	wire [WIDTH*2-1+0:0] tmp00_41_19;
	wire [WIDTH*2-1+0:0] tmp00_41_20;
	wire [WIDTH*2-1+0:0] tmp00_41_21;
	wire [WIDTH*2-1+0:0] tmp00_41_22;
	wire [WIDTH*2-1+0:0] tmp00_41_23;
	wire [WIDTH*2-1+0:0] tmp00_41_24;
	wire [WIDTH*2-1+0:0] tmp00_41_25;
	wire [WIDTH*2-1+0:0] tmp00_41_26;
	wire [WIDTH*2-1+0:0] tmp00_41_27;
	wire [WIDTH*2-1+0:0] tmp00_41_28;
	wire [WIDTH*2-1+0:0] tmp00_41_29;
	wire [WIDTH*2-1+0:0] tmp00_41_30;
	wire [WIDTH*2-1+0:0] tmp00_41_31;
	wire [WIDTH*2-1+0:0] tmp00_41_32;
	wire [WIDTH*2-1+0:0] tmp00_41_33;
	wire [WIDTH*2-1+0:0] tmp00_41_34;
	wire [WIDTH*2-1+0:0] tmp00_41_35;
	wire [WIDTH*2-1+0:0] tmp00_41_36;
	wire [WIDTH*2-1+0:0] tmp00_41_37;
	wire [WIDTH*2-1+0:0] tmp00_41_38;
	wire [WIDTH*2-1+0:0] tmp00_41_39;
	wire [WIDTH*2-1+0:0] tmp00_41_40;
	wire [WIDTH*2-1+0:0] tmp00_41_41;
	wire [WIDTH*2-1+0:0] tmp00_41_42;
	wire [WIDTH*2-1+0:0] tmp00_41_43;
	wire [WIDTH*2-1+0:0] tmp00_41_44;
	wire [WIDTH*2-1+0:0] tmp00_41_45;
	wire [WIDTH*2-1+0:0] tmp00_41_46;
	wire [WIDTH*2-1+0:0] tmp00_41_47;
	wire [WIDTH*2-1+0:0] tmp00_41_48;
	wire [WIDTH*2-1+0:0] tmp00_41_49;
	wire [WIDTH*2-1+0:0] tmp00_41_50;
	wire [WIDTH*2-1+0:0] tmp00_41_51;
	wire [WIDTH*2-1+0:0] tmp00_41_52;
	wire [WIDTH*2-1+0:0] tmp00_41_53;
	wire [WIDTH*2-1+0:0] tmp00_41_54;
	wire [WIDTH*2-1+0:0] tmp00_41_55;
	wire [WIDTH*2-1+0:0] tmp00_41_56;
	wire [WIDTH*2-1+0:0] tmp00_41_57;
	wire [WIDTH*2-1+0:0] tmp00_41_58;
	wire [WIDTH*2-1+0:0] tmp00_41_59;
	wire [WIDTH*2-1+0:0] tmp00_41_60;
	wire [WIDTH*2-1+0:0] tmp00_41_61;
	wire [WIDTH*2-1+0:0] tmp00_41_62;
	wire [WIDTH*2-1+0:0] tmp00_41_63;
	wire [WIDTH*2-1+0:0] tmp00_41_64;
	wire [WIDTH*2-1+0:0] tmp00_41_65;
	wire [WIDTH*2-1+0:0] tmp00_41_66;
	wire [WIDTH*2-1+0:0] tmp00_41_67;
	wire [WIDTH*2-1+0:0] tmp00_41_68;
	wire [WIDTH*2-1+0:0] tmp00_41_69;
	wire [WIDTH*2-1+0:0] tmp00_41_70;
	wire [WIDTH*2-1+0:0] tmp00_41_71;
	wire [WIDTH*2-1+0:0] tmp00_41_72;
	wire [WIDTH*2-1+0:0] tmp00_41_73;
	wire [WIDTH*2-1+0:0] tmp00_41_74;
	wire [WIDTH*2-1+0:0] tmp00_41_75;
	wire [WIDTH*2-1+0:0] tmp00_41_76;
	wire [WIDTH*2-1+0:0] tmp00_41_77;
	wire [WIDTH*2-1+0:0] tmp00_41_78;
	wire [WIDTH*2-1+0:0] tmp00_41_79;
	wire [WIDTH*2-1+0:0] tmp00_41_80;
	wire [WIDTH*2-1+0:0] tmp00_41_81;
	wire [WIDTH*2-1+0:0] tmp00_41_82;
	wire [WIDTH*2-1+0:0] tmp00_41_83;
	wire [WIDTH*2-1+0:0] tmp00_42_0;
	wire [WIDTH*2-1+0:0] tmp00_42_1;
	wire [WIDTH*2-1+0:0] tmp00_42_2;
	wire [WIDTH*2-1+0:0] tmp00_42_3;
	wire [WIDTH*2-1+0:0] tmp00_42_4;
	wire [WIDTH*2-1+0:0] tmp00_42_5;
	wire [WIDTH*2-1+0:0] tmp00_42_6;
	wire [WIDTH*2-1+0:0] tmp00_42_7;
	wire [WIDTH*2-1+0:0] tmp00_42_8;
	wire [WIDTH*2-1+0:0] tmp00_42_9;
	wire [WIDTH*2-1+0:0] tmp00_42_10;
	wire [WIDTH*2-1+0:0] tmp00_42_11;
	wire [WIDTH*2-1+0:0] tmp00_42_12;
	wire [WIDTH*2-1+0:0] tmp00_42_13;
	wire [WIDTH*2-1+0:0] tmp00_42_14;
	wire [WIDTH*2-1+0:0] tmp00_42_15;
	wire [WIDTH*2-1+0:0] tmp00_42_16;
	wire [WIDTH*2-1+0:0] tmp00_42_17;
	wire [WIDTH*2-1+0:0] tmp00_42_18;
	wire [WIDTH*2-1+0:0] tmp00_42_19;
	wire [WIDTH*2-1+0:0] tmp00_42_20;
	wire [WIDTH*2-1+0:0] tmp00_42_21;
	wire [WIDTH*2-1+0:0] tmp00_42_22;
	wire [WIDTH*2-1+0:0] tmp00_42_23;
	wire [WIDTH*2-1+0:0] tmp00_42_24;
	wire [WIDTH*2-1+0:0] tmp00_42_25;
	wire [WIDTH*2-1+0:0] tmp00_42_26;
	wire [WIDTH*2-1+0:0] tmp00_42_27;
	wire [WIDTH*2-1+0:0] tmp00_42_28;
	wire [WIDTH*2-1+0:0] tmp00_42_29;
	wire [WIDTH*2-1+0:0] tmp00_42_30;
	wire [WIDTH*2-1+0:0] tmp00_42_31;
	wire [WIDTH*2-1+0:0] tmp00_42_32;
	wire [WIDTH*2-1+0:0] tmp00_42_33;
	wire [WIDTH*2-1+0:0] tmp00_42_34;
	wire [WIDTH*2-1+0:0] tmp00_42_35;
	wire [WIDTH*2-1+0:0] tmp00_42_36;
	wire [WIDTH*2-1+0:0] tmp00_42_37;
	wire [WIDTH*2-1+0:0] tmp00_42_38;
	wire [WIDTH*2-1+0:0] tmp00_42_39;
	wire [WIDTH*2-1+0:0] tmp00_42_40;
	wire [WIDTH*2-1+0:0] tmp00_42_41;
	wire [WIDTH*2-1+0:0] tmp00_42_42;
	wire [WIDTH*2-1+0:0] tmp00_42_43;
	wire [WIDTH*2-1+0:0] tmp00_42_44;
	wire [WIDTH*2-1+0:0] tmp00_42_45;
	wire [WIDTH*2-1+0:0] tmp00_42_46;
	wire [WIDTH*2-1+0:0] tmp00_42_47;
	wire [WIDTH*2-1+0:0] tmp00_42_48;
	wire [WIDTH*2-1+0:0] tmp00_42_49;
	wire [WIDTH*2-1+0:0] tmp00_42_50;
	wire [WIDTH*2-1+0:0] tmp00_42_51;
	wire [WIDTH*2-1+0:0] tmp00_42_52;
	wire [WIDTH*2-1+0:0] tmp00_42_53;
	wire [WIDTH*2-1+0:0] tmp00_42_54;
	wire [WIDTH*2-1+0:0] tmp00_42_55;
	wire [WIDTH*2-1+0:0] tmp00_42_56;
	wire [WIDTH*2-1+0:0] tmp00_42_57;
	wire [WIDTH*2-1+0:0] tmp00_42_58;
	wire [WIDTH*2-1+0:0] tmp00_42_59;
	wire [WIDTH*2-1+0:0] tmp00_42_60;
	wire [WIDTH*2-1+0:0] tmp00_42_61;
	wire [WIDTH*2-1+0:0] tmp00_42_62;
	wire [WIDTH*2-1+0:0] tmp00_42_63;
	wire [WIDTH*2-1+0:0] tmp00_42_64;
	wire [WIDTH*2-1+0:0] tmp00_42_65;
	wire [WIDTH*2-1+0:0] tmp00_42_66;
	wire [WIDTH*2-1+0:0] tmp00_42_67;
	wire [WIDTH*2-1+0:0] tmp00_42_68;
	wire [WIDTH*2-1+0:0] tmp00_42_69;
	wire [WIDTH*2-1+0:0] tmp00_42_70;
	wire [WIDTH*2-1+0:0] tmp00_42_71;
	wire [WIDTH*2-1+0:0] tmp00_42_72;
	wire [WIDTH*2-1+0:0] tmp00_42_73;
	wire [WIDTH*2-1+0:0] tmp00_42_74;
	wire [WIDTH*2-1+0:0] tmp00_42_75;
	wire [WIDTH*2-1+0:0] tmp00_42_76;
	wire [WIDTH*2-1+0:0] tmp00_42_77;
	wire [WIDTH*2-1+0:0] tmp00_42_78;
	wire [WIDTH*2-1+0:0] tmp00_42_79;
	wire [WIDTH*2-1+0:0] tmp00_42_80;
	wire [WIDTH*2-1+0:0] tmp00_42_81;
	wire [WIDTH*2-1+0:0] tmp00_42_82;
	wire [WIDTH*2-1+0:0] tmp00_42_83;
	wire [WIDTH*2-1+0:0] tmp00_43_0;
	wire [WIDTH*2-1+0:0] tmp00_43_1;
	wire [WIDTH*2-1+0:0] tmp00_43_2;
	wire [WIDTH*2-1+0:0] tmp00_43_3;
	wire [WIDTH*2-1+0:0] tmp00_43_4;
	wire [WIDTH*2-1+0:0] tmp00_43_5;
	wire [WIDTH*2-1+0:0] tmp00_43_6;
	wire [WIDTH*2-1+0:0] tmp00_43_7;
	wire [WIDTH*2-1+0:0] tmp00_43_8;
	wire [WIDTH*2-1+0:0] tmp00_43_9;
	wire [WIDTH*2-1+0:0] tmp00_43_10;
	wire [WIDTH*2-1+0:0] tmp00_43_11;
	wire [WIDTH*2-1+0:0] tmp00_43_12;
	wire [WIDTH*2-1+0:0] tmp00_43_13;
	wire [WIDTH*2-1+0:0] tmp00_43_14;
	wire [WIDTH*2-1+0:0] tmp00_43_15;
	wire [WIDTH*2-1+0:0] tmp00_43_16;
	wire [WIDTH*2-1+0:0] tmp00_43_17;
	wire [WIDTH*2-1+0:0] tmp00_43_18;
	wire [WIDTH*2-1+0:0] tmp00_43_19;
	wire [WIDTH*2-1+0:0] tmp00_43_20;
	wire [WIDTH*2-1+0:0] tmp00_43_21;
	wire [WIDTH*2-1+0:0] tmp00_43_22;
	wire [WIDTH*2-1+0:0] tmp00_43_23;
	wire [WIDTH*2-1+0:0] tmp00_43_24;
	wire [WIDTH*2-1+0:0] tmp00_43_25;
	wire [WIDTH*2-1+0:0] tmp00_43_26;
	wire [WIDTH*2-1+0:0] tmp00_43_27;
	wire [WIDTH*2-1+0:0] tmp00_43_28;
	wire [WIDTH*2-1+0:0] tmp00_43_29;
	wire [WIDTH*2-1+0:0] tmp00_43_30;
	wire [WIDTH*2-1+0:0] tmp00_43_31;
	wire [WIDTH*2-1+0:0] tmp00_43_32;
	wire [WIDTH*2-1+0:0] tmp00_43_33;
	wire [WIDTH*2-1+0:0] tmp00_43_34;
	wire [WIDTH*2-1+0:0] tmp00_43_35;
	wire [WIDTH*2-1+0:0] tmp00_43_36;
	wire [WIDTH*2-1+0:0] tmp00_43_37;
	wire [WIDTH*2-1+0:0] tmp00_43_38;
	wire [WIDTH*2-1+0:0] tmp00_43_39;
	wire [WIDTH*2-1+0:0] tmp00_43_40;
	wire [WIDTH*2-1+0:0] tmp00_43_41;
	wire [WIDTH*2-1+0:0] tmp00_43_42;
	wire [WIDTH*2-1+0:0] tmp00_43_43;
	wire [WIDTH*2-1+0:0] tmp00_43_44;
	wire [WIDTH*2-1+0:0] tmp00_43_45;
	wire [WIDTH*2-1+0:0] tmp00_43_46;
	wire [WIDTH*2-1+0:0] tmp00_43_47;
	wire [WIDTH*2-1+0:0] tmp00_43_48;
	wire [WIDTH*2-1+0:0] tmp00_43_49;
	wire [WIDTH*2-1+0:0] tmp00_43_50;
	wire [WIDTH*2-1+0:0] tmp00_43_51;
	wire [WIDTH*2-1+0:0] tmp00_43_52;
	wire [WIDTH*2-1+0:0] tmp00_43_53;
	wire [WIDTH*2-1+0:0] tmp00_43_54;
	wire [WIDTH*2-1+0:0] tmp00_43_55;
	wire [WIDTH*2-1+0:0] tmp00_43_56;
	wire [WIDTH*2-1+0:0] tmp00_43_57;
	wire [WIDTH*2-1+0:0] tmp00_43_58;
	wire [WIDTH*2-1+0:0] tmp00_43_59;
	wire [WIDTH*2-1+0:0] tmp00_43_60;
	wire [WIDTH*2-1+0:0] tmp00_43_61;
	wire [WIDTH*2-1+0:0] tmp00_43_62;
	wire [WIDTH*2-1+0:0] tmp00_43_63;
	wire [WIDTH*2-1+0:0] tmp00_43_64;
	wire [WIDTH*2-1+0:0] tmp00_43_65;
	wire [WIDTH*2-1+0:0] tmp00_43_66;
	wire [WIDTH*2-1+0:0] tmp00_43_67;
	wire [WIDTH*2-1+0:0] tmp00_43_68;
	wire [WIDTH*2-1+0:0] tmp00_43_69;
	wire [WIDTH*2-1+0:0] tmp00_43_70;
	wire [WIDTH*2-1+0:0] tmp00_43_71;
	wire [WIDTH*2-1+0:0] tmp00_43_72;
	wire [WIDTH*2-1+0:0] tmp00_43_73;
	wire [WIDTH*2-1+0:0] tmp00_43_74;
	wire [WIDTH*2-1+0:0] tmp00_43_75;
	wire [WIDTH*2-1+0:0] tmp00_43_76;
	wire [WIDTH*2-1+0:0] tmp00_43_77;
	wire [WIDTH*2-1+0:0] tmp00_43_78;
	wire [WIDTH*2-1+0:0] tmp00_43_79;
	wire [WIDTH*2-1+0:0] tmp00_43_80;
	wire [WIDTH*2-1+0:0] tmp00_43_81;
	wire [WIDTH*2-1+0:0] tmp00_43_82;
	wire [WIDTH*2-1+0:0] tmp00_43_83;
	wire [WIDTH*2-1+0:0] tmp00_44_0;
	wire [WIDTH*2-1+0:0] tmp00_44_1;
	wire [WIDTH*2-1+0:0] tmp00_44_2;
	wire [WIDTH*2-1+0:0] tmp00_44_3;
	wire [WIDTH*2-1+0:0] tmp00_44_4;
	wire [WIDTH*2-1+0:0] tmp00_44_5;
	wire [WIDTH*2-1+0:0] tmp00_44_6;
	wire [WIDTH*2-1+0:0] tmp00_44_7;
	wire [WIDTH*2-1+0:0] tmp00_44_8;
	wire [WIDTH*2-1+0:0] tmp00_44_9;
	wire [WIDTH*2-1+0:0] tmp00_44_10;
	wire [WIDTH*2-1+0:0] tmp00_44_11;
	wire [WIDTH*2-1+0:0] tmp00_44_12;
	wire [WIDTH*2-1+0:0] tmp00_44_13;
	wire [WIDTH*2-1+0:0] tmp00_44_14;
	wire [WIDTH*2-1+0:0] tmp00_44_15;
	wire [WIDTH*2-1+0:0] tmp00_44_16;
	wire [WIDTH*2-1+0:0] tmp00_44_17;
	wire [WIDTH*2-1+0:0] tmp00_44_18;
	wire [WIDTH*2-1+0:0] tmp00_44_19;
	wire [WIDTH*2-1+0:0] tmp00_44_20;
	wire [WIDTH*2-1+0:0] tmp00_44_21;
	wire [WIDTH*2-1+0:0] tmp00_44_22;
	wire [WIDTH*2-1+0:0] tmp00_44_23;
	wire [WIDTH*2-1+0:0] tmp00_44_24;
	wire [WIDTH*2-1+0:0] tmp00_44_25;
	wire [WIDTH*2-1+0:0] tmp00_44_26;
	wire [WIDTH*2-1+0:0] tmp00_44_27;
	wire [WIDTH*2-1+0:0] tmp00_44_28;
	wire [WIDTH*2-1+0:0] tmp00_44_29;
	wire [WIDTH*2-1+0:0] tmp00_44_30;
	wire [WIDTH*2-1+0:0] tmp00_44_31;
	wire [WIDTH*2-1+0:0] tmp00_44_32;
	wire [WIDTH*2-1+0:0] tmp00_44_33;
	wire [WIDTH*2-1+0:0] tmp00_44_34;
	wire [WIDTH*2-1+0:0] tmp00_44_35;
	wire [WIDTH*2-1+0:0] tmp00_44_36;
	wire [WIDTH*2-1+0:0] tmp00_44_37;
	wire [WIDTH*2-1+0:0] tmp00_44_38;
	wire [WIDTH*2-1+0:0] tmp00_44_39;
	wire [WIDTH*2-1+0:0] tmp00_44_40;
	wire [WIDTH*2-1+0:0] tmp00_44_41;
	wire [WIDTH*2-1+0:0] tmp00_44_42;
	wire [WIDTH*2-1+0:0] tmp00_44_43;
	wire [WIDTH*2-1+0:0] tmp00_44_44;
	wire [WIDTH*2-1+0:0] tmp00_44_45;
	wire [WIDTH*2-1+0:0] tmp00_44_46;
	wire [WIDTH*2-1+0:0] tmp00_44_47;
	wire [WIDTH*2-1+0:0] tmp00_44_48;
	wire [WIDTH*2-1+0:0] tmp00_44_49;
	wire [WIDTH*2-1+0:0] tmp00_44_50;
	wire [WIDTH*2-1+0:0] tmp00_44_51;
	wire [WIDTH*2-1+0:0] tmp00_44_52;
	wire [WIDTH*2-1+0:0] tmp00_44_53;
	wire [WIDTH*2-1+0:0] tmp00_44_54;
	wire [WIDTH*2-1+0:0] tmp00_44_55;
	wire [WIDTH*2-1+0:0] tmp00_44_56;
	wire [WIDTH*2-1+0:0] tmp00_44_57;
	wire [WIDTH*2-1+0:0] tmp00_44_58;
	wire [WIDTH*2-1+0:0] tmp00_44_59;
	wire [WIDTH*2-1+0:0] tmp00_44_60;
	wire [WIDTH*2-1+0:0] tmp00_44_61;
	wire [WIDTH*2-1+0:0] tmp00_44_62;
	wire [WIDTH*2-1+0:0] tmp00_44_63;
	wire [WIDTH*2-1+0:0] tmp00_44_64;
	wire [WIDTH*2-1+0:0] tmp00_44_65;
	wire [WIDTH*2-1+0:0] tmp00_44_66;
	wire [WIDTH*2-1+0:0] tmp00_44_67;
	wire [WIDTH*2-1+0:0] tmp00_44_68;
	wire [WIDTH*2-1+0:0] tmp00_44_69;
	wire [WIDTH*2-1+0:0] tmp00_44_70;
	wire [WIDTH*2-1+0:0] tmp00_44_71;
	wire [WIDTH*2-1+0:0] tmp00_44_72;
	wire [WIDTH*2-1+0:0] tmp00_44_73;
	wire [WIDTH*2-1+0:0] tmp00_44_74;
	wire [WIDTH*2-1+0:0] tmp00_44_75;
	wire [WIDTH*2-1+0:0] tmp00_44_76;
	wire [WIDTH*2-1+0:0] tmp00_44_77;
	wire [WIDTH*2-1+0:0] tmp00_44_78;
	wire [WIDTH*2-1+0:0] tmp00_44_79;
	wire [WIDTH*2-1+0:0] tmp00_44_80;
	wire [WIDTH*2-1+0:0] tmp00_44_81;
	wire [WIDTH*2-1+0:0] tmp00_44_82;
	wire [WIDTH*2-1+0:0] tmp00_44_83;
	wire [WIDTH*2-1+0:0] tmp00_45_0;
	wire [WIDTH*2-1+0:0] tmp00_45_1;
	wire [WIDTH*2-1+0:0] tmp00_45_2;
	wire [WIDTH*2-1+0:0] tmp00_45_3;
	wire [WIDTH*2-1+0:0] tmp00_45_4;
	wire [WIDTH*2-1+0:0] tmp00_45_5;
	wire [WIDTH*2-1+0:0] tmp00_45_6;
	wire [WIDTH*2-1+0:0] tmp00_45_7;
	wire [WIDTH*2-1+0:0] tmp00_45_8;
	wire [WIDTH*2-1+0:0] tmp00_45_9;
	wire [WIDTH*2-1+0:0] tmp00_45_10;
	wire [WIDTH*2-1+0:0] tmp00_45_11;
	wire [WIDTH*2-1+0:0] tmp00_45_12;
	wire [WIDTH*2-1+0:0] tmp00_45_13;
	wire [WIDTH*2-1+0:0] tmp00_45_14;
	wire [WIDTH*2-1+0:0] tmp00_45_15;
	wire [WIDTH*2-1+0:0] tmp00_45_16;
	wire [WIDTH*2-1+0:0] tmp00_45_17;
	wire [WIDTH*2-1+0:0] tmp00_45_18;
	wire [WIDTH*2-1+0:0] tmp00_45_19;
	wire [WIDTH*2-1+0:0] tmp00_45_20;
	wire [WIDTH*2-1+0:0] tmp00_45_21;
	wire [WIDTH*2-1+0:0] tmp00_45_22;
	wire [WIDTH*2-1+0:0] tmp00_45_23;
	wire [WIDTH*2-1+0:0] tmp00_45_24;
	wire [WIDTH*2-1+0:0] tmp00_45_25;
	wire [WIDTH*2-1+0:0] tmp00_45_26;
	wire [WIDTH*2-1+0:0] tmp00_45_27;
	wire [WIDTH*2-1+0:0] tmp00_45_28;
	wire [WIDTH*2-1+0:0] tmp00_45_29;
	wire [WIDTH*2-1+0:0] tmp00_45_30;
	wire [WIDTH*2-1+0:0] tmp00_45_31;
	wire [WIDTH*2-1+0:0] tmp00_45_32;
	wire [WIDTH*2-1+0:0] tmp00_45_33;
	wire [WIDTH*2-1+0:0] tmp00_45_34;
	wire [WIDTH*2-1+0:0] tmp00_45_35;
	wire [WIDTH*2-1+0:0] tmp00_45_36;
	wire [WIDTH*2-1+0:0] tmp00_45_37;
	wire [WIDTH*2-1+0:0] tmp00_45_38;
	wire [WIDTH*2-1+0:0] tmp00_45_39;
	wire [WIDTH*2-1+0:0] tmp00_45_40;
	wire [WIDTH*2-1+0:0] tmp00_45_41;
	wire [WIDTH*2-1+0:0] tmp00_45_42;
	wire [WIDTH*2-1+0:0] tmp00_45_43;
	wire [WIDTH*2-1+0:0] tmp00_45_44;
	wire [WIDTH*2-1+0:0] tmp00_45_45;
	wire [WIDTH*2-1+0:0] tmp00_45_46;
	wire [WIDTH*2-1+0:0] tmp00_45_47;
	wire [WIDTH*2-1+0:0] tmp00_45_48;
	wire [WIDTH*2-1+0:0] tmp00_45_49;
	wire [WIDTH*2-1+0:0] tmp00_45_50;
	wire [WIDTH*2-1+0:0] tmp00_45_51;
	wire [WIDTH*2-1+0:0] tmp00_45_52;
	wire [WIDTH*2-1+0:0] tmp00_45_53;
	wire [WIDTH*2-1+0:0] tmp00_45_54;
	wire [WIDTH*2-1+0:0] tmp00_45_55;
	wire [WIDTH*2-1+0:0] tmp00_45_56;
	wire [WIDTH*2-1+0:0] tmp00_45_57;
	wire [WIDTH*2-1+0:0] tmp00_45_58;
	wire [WIDTH*2-1+0:0] tmp00_45_59;
	wire [WIDTH*2-1+0:0] tmp00_45_60;
	wire [WIDTH*2-1+0:0] tmp00_45_61;
	wire [WIDTH*2-1+0:0] tmp00_45_62;
	wire [WIDTH*2-1+0:0] tmp00_45_63;
	wire [WIDTH*2-1+0:0] tmp00_45_64;
	wire [WIDTH*2-1+0:0] tmp00_45_65;
	wire [WIDTH*2-1+0:0] tmp00_45_66;
	wire [WIDTH*2-1+0:0] tmp00_45_67;
	wire [WIDTH*2-1+0:0] tmp00_45_68;
	wire [WIDTH*2-1+0:0] tmp00_45_69;
	wire [WIDTH*2-1+0:0] tmp00_45_70;
	wire [WIDTH*2-1+0:0] tmp00_45_71;
	wire [WIDTH*2-1+0:0] tmp00_45_72;
	wire [WIDTH*2-1+0:0] tmp00_45_73;
	wire [WIDTH*2-1+0:0] tmp00_45_74;
	wire [WIDTH*2-1+0:0] tmp00_45_75;
	wire [WIDTH*2-1+0:0] tmp00_45_76;
	wire [WIDTH*2-1+0:0] tmp00_45_77;
	wire [WIDTH*2-1+0:0] tmp00_45_78;
	wire [WIDTH*2-1+0:0] tmp00_45_79;
	wire [WIDTH*2-1+0:0] tmp00_45_80;
	wire [WIDTH*2-1+0:0] tmp00_45_81;
	wire [WIDTH*2-1+0:0] tmp00_45_82;
	wire [WIDTH*2-1+0:0] tmp00_45_83;
	wire [WIDTH*2-1+0:0] tmp00_46_0;
	wire [WIDTH*2-1+0:0] tmp00_46_1;
	wire [WIDTH*2-1+0:0] tmp00_46_2;
	wire [WIDTH*2-1+0:0] tmp00_46_3;
	wire [WIDTH*2-1+0:0] tmp00_46_4;
	wire [WIDTH*2-1+0:0] tmp00_46_5;
	wire [WIDTH*2-1+0:0] tmp00_46_6;
	wire [WIDTH*2-1+0:0] tmp00_46_7;
	wire [WIDTH*2-1+0:0] tmp00_46_8;
	wire [WIDTH*2-1+0:0] tmp00_46_9;
	wire [WIDTH*2-1+0:0] tmp00_46_10;
	wire [WIDTH*2-1+0:0] tmp00_46_11;
	wire [WIDTH*2-1+0:0] tmp00_46_12;
	wire [WIDTH*2-1+0:0] tmp00_46_13;
	wire [WIDTH*2-1+0:0] tmp00_46_14;
	wire [WIDTH*2-1+0:0] tmp00_46_15;
	wire [WIDTH*2-1+0:0] tmp00_46_16;
	wire [WIDTH*2-1+0:0] tmp00_46_17;
	wire [WIDTH*2-1+0:0] tmp00_46_18;
	wire [WIDTH*2-1+0:0] tmp00_46_19;
	wire [WIDTH*2-1+0:0] tmp00_46_20;
	wire [WIDTH*2-1+0:0] tmp00_46_21;
	wire [WIDTH*2-1+0:0] tmp00_46_22;
	wire [WIDTH*2-1+0:0] tmp00_46_23;
	wire [WIDTH*2-1+0:0] tmp00_46_24;
	wire [WIDTH*2-1+0:0] tmp00_46_25;
	wire [WIDTH*2-1+0:0] tmp00_46_26;
	wire [WIDTH*2-1+0:0] tmp00_46_27;
	wire [WIDTH*2-1+0:0] tmp00_46_28;
	wire [WIDTH*2-1+0:0] tmp00_46_29;
	wire [WIDTH*2-1+0:0] tmp00_46_30;
	wire [WIDTH*2-1+0:0] tmp00_46_31;
	wire [WIDTH*2-1+0:0] tmp00_46_32;
	wire [WIDTH*2-1+0:0] tmp00_46_33;
	wire [WIDTH*2-1+0:0] tmp00_46_34;
	wire [WIDTH*2-1+0:0] tmp00_46_35;
	wire [WIDTH*2-1+0:0] tmp00_46_36;
	wire [WIDTH*2-1+0:0] tmp00_46_37;
	wire [WIDTH*2-1+0:0] tmp00_46_38;
	wire [WIDTH*2-1+0:0] tmp00_46_39;
	wire [WIDTH*2-1+0:0] tmp00_46_40;
	wire [WIDTH*2-1+0:0] tmp00_46_41;
	wire [WIDTH*2-1+0:0] tmp00_46_42;
	wire [WIDTH*2-1+0:0] tmp00_46_43;
	wire [WIDTH*2-1+0:0] tmp00_46_44;
	wire [WIDTH*2-1+0:0] tmp00_46_45;
	wire [WIDTH*2-1+0:0] tmp00_46_46;
	wire [WIDTH*2-1+0:0] tmp00_46_47;
	wire [WIDTH*2-1+0:0] tmp00_46_48;
	wire [WIDTH*2-1+0:0] tmp00_46_49;
	wire [WIDTH*2-1+0:0] tmp00_46_50;
	wire [WIDTH*2-1+0:0] tmp00_46_51;
	wire [WIDTH*2-1+0:0] tmp00_46_52;
	wire [WIDTH*2-1+0:0] tmp00_46_53;
	wire [WIDTH*2-1+0:0] tmp00_46_54;
	wire [WIDTH*2-1+0:0] tmp00_46_55;
	wire [WIDTH*2-1+0:0] tmp00_46_56;
	wire [WIDTH*2-1+0:0] tmp00_46_57;
	wire [WIDTH*2-1+0:0] tmp00_46_58;
	wire [WIDTH*2-1+0:0] tmp00_46_59;
	wire [WIDTH*2-1+0:0] tmp00_46_60;
	wire [WIDTH*2-1+0:0] tmp00_46_61;
	wire [WIDTH*2-1+0:0] tmp00_46_62;
	wire [WIDTH*2-1+0:0] tmp00_46_63;
	wire [WIDTH*2-1+0:0] tmp00_46_64;
	wire [WIDTH*2-1+0:0] tmp00_46_65;
	wire [WIDTH*2-1+0:0] tmp00_46_66;
	wire [WIDTH*2-1+0:0] tmp00_46_67;
	wire [WIDTH*2-1+0:0] tmp00_46_68;
	wire [WIDTH*2-1+0:0] tmp00_46_69;
	wire [WIDTH*2-1+0:0] tmp00_46_70;
	wire [WIDTH*2-1+0:0] tmp00_46_71;
	wire [WIDTH*2-1+0:0] tmp00_46_72;
	wire [WIDTH*2-1+0:0] tmp00_46_73;
	wire [WIDTH*2-1+0:0] tmp00_46_74;
	wire [WIDTH*2-1+0:0] tmp00_46_75;
	wire [WIDTH*2-1+0:0] tmp00_46_76;
	wire [WIDTH*2-1+0:0] tmp00_46_77;
	wire [WIDTH*2-1+0:0] tmp00_46_78;
	wire [WIDTH*2-1+0:0] tmp00_46_79;
	wire [WIDTH*2-1+0:0] tmp00_46_80;
	wire [WIDTH*2-1+0:0] tmp00_46_81;
	wire [WIDTH*2-1+0:0] tmp00_46_82;
	wire [WIDTH*2-1+0:0] tmp00_46_83;
	wire [WIDTH*2-1+0:0] tmp00_47_0;
	wire [WIDTH*2-1+0:0] tmp00_47_1;
	wire [WIDTH*2-1+0:0] tmp00_47_2;
	wire [WIDTH*2-1+0:0] tmp00_47_3;
	wire [WIDTH*2-1+0:0] tmp00_47_4;
	wire [WIDTH*2-1+0:0] tmp00_47_5;
	wire [WIDTH*2-1+0:0] tmp00_47_6;
	wire [WIDTH*2-1+0:0] tmp00_47_7;
	wire [WIDTH*2-1+0:0] tmp00_47_8;
	wire [WIDTH*2-1+0:0] tmp00_47_9;
	wire [WIDTH*2-1+0:0] tmp00_47_10;
	wire [WIDTH*2-1+0:0] tmp00_47_11;
	wire [WIDTH*2-1+0:0] tmp00_47_12;
	wire [WIDTH*2-1+0:0] tmp00_47_13;
	wire [WIDTH*2-1+0:0] tmp00_47_14;
	wire [WIDTH*2-1+0:0] tmp00_47_15;
	wire [WIDTH*2-1+0:0] tmp00_47_16;
	wire [WIDTH*2-1+0:0] tmp00_47_17;
	wire [WIDTH*2-1+0:0] tmp00_47_18;
	wire [WIDTH*2-1+0:0] tmp00_47_19;
	wire [WIDTH*2-1+0:0] tmp00_47_20;
	wire [WIDTH*2-1+0:0] tmp00_47_21;
	wire [WIDTH*2-1+0:0] tmp00_47_22;
	wire [WIDTH*2-1+0:0] tmp00_47_23;
	wire [WIDTH*2-1+0:0] tmp00_47_24;
	wire [WIDTH*2-1+0:0] tmp00_47_25;
	wire [WIDTH*2-1+0:0] tmp00_47_26;
	wire [WIDTH*2-1+0:0] tmp00_47_27;
	wire [WIDTH*2-1+0:0] tmp00_47_28;
	wire [WIDTH*2-1+0:0] tmp00_47_29;
	wire [WIDTH*2-1+0:0] tmp00_47_30;
	wire [WIDTH*2-1+0:0] tmp00_47_31;
	wire [WIDTH*2-1+0:0] tmp00_47_32;
	wire [WIDTH*2-1+0:0] tmp00_47_33;
	wire [WIDTH*2-1+0:0] tmp00_47_34;
	wire [WIDTH*2-1+0:0] tmp00_47_35;
	wire [WIDTH*2-1+0:0] tmp00_47_36;
	wire [WIDTH*2-1+0:0] tmp00_47_37;
	wire [WIDTH*2-1+0:0] tmp00_47_38;
	wire [WIDTH*2-1+0:0] tmp00_47_39;
	wire [WIDTH*2-1+0:0] tmp00_47_40;
	wire [WIDTH*2-1+0:0] tmp00_47_41;
	wire [WIDTH*2-1+0:0] tmp00_47_42;
	wire [WIDTH*2-1+0:0] tmp00_47_43;
	wire [WIDTH*2-1+0:0] tmp00_47_44;
	wire [WIDTH*2-1+0:0] tmp00_47_45;
	wire [WIDTH*2-1+0:0] tmp00_47_46;
	wire [WIDTH*2-1+0:0] tmp00_47_47;
	wire [WIDTH*2-1+0:0] tmp00_47_48;
	wire [WIDTH*2-1+0:0] tmp00_47_49;
	wire [WIDTH*2-1+0:0] tmp00_47_50;
	wire [WIDTH*2-1+0:0] tmp00_47_51;
	wire [WIDTH*2-1+0:0] tmp00_47_52;
	wire [WIDTH*2-1+0:0] tmp00_47_53;
	wire [WIDTH*2-1+0:0] tmp00_47_54;
	wire [WIDTH*2-1+0:0] tmp00_47_55;
	wire [WIDTH*2-1+0:0] tmp00_47_56;
	wire [WIDTH*2-1+0:0] tmp00_47_57;
	wire [WIDTH*2-1+0:0] tmp00_47_58;
	wire [WIDTH*2-1+0:0] tmp00_47_59;
	wire [WIDTH*2-1+0:0] tmp00_47_60;
	wire [WIDTH*2-1+0:0] tmp00_47_61;
	wire [WIDTH*2-1+0:0] tmp00_47_62;
	wire [WIDTH*2-1+0:0] tmp00_47_63;
	wire [WIDTH*2-1+0:0] tmp00_47_64;
	wire [WIDTH*2-1+0:0] tmp00_47_65;
	wire [WIDTH*2-1+0:0] tmp00_47_66;
	wire [WIDTH*2-1+0:0] tmp00_47_67;
	wire [WIDTH*2-1+0:0] tmp00_47_68;
	wire [WIDTH*2-1+0:0] tmp00_47_69;
	wire [WIDTH*2-1+0:0] tmp00_47_70;
	wire [WIDTH*2-1+0:0] tmp00_47_71;
	wire [WIDTH*2-1+0:0] tmp00_47_72;
	wire [WIDTH*2-1+0:0] tmp00_47_73;
	wire [WIDTH*2-1+0:0] tmp00_47_74;
	wire [WIDTH*2-1+0:0] tmp00_47_75;
	wire [WIDTH*2-1+0:0] tmp00_47_76;
	wire [WIDTH*2-1+0:0] tmp00_47_77;
	wire [WIDTH*2-1+0:0] tmp00_47_78;
	wire [WIDTH*2-1+0:0] tmp00_47_79;
	wire [WIDTH*2-1+0:0] tmp00_47_80;
	wire [WIDTH*2-1+0:0] tmp00_47_81;
	wire [WIDTH*2-1+0:0] tmp00_47_82;
	wire [WIDTH*2-1+0:0] tmp00_47_83;
	wire [WIDTH*2-1+0:0] tmp00_48_0;
	wire [WIDTH*2-1+0:0] tmp00_48_1;
	wire [WIDTH*2-1+0:0] tmp00_48_2;
	wire [WIDTH*2-1+0:0] tmp00_48_3;
	wire [WIDTH*2-1+0:0] tmp00_48_4;
	wire [WIDTH*2-1+0:0] tmp00_48_5;
	wire [WIDTH*2-1+0:0] tmp00_48_6;
	wire [WIDTH*2-1+0:0] tmp00_48_7;
	wire [WIDTH*2-1+0:0] tmp00_48_8;
	wire [WIDTH*2-1+0:0] tmp00_48_9;
	wire [WIDTH*2-1+0:0] tmp00_48_10;
	wire [WIDTH*2-1+0:0] tmp00_48_11;
	wire [WIDTH*2-1+0:0] tmp00_48_12;
	wire [WIDTH*2-1+0:0] tmp00_48_13;
	wire [WIDTH*2-1+0:0] tmp00_48_14;
	wire [WIDTH*2-1+0:0] tmp00_48_15;
	wire [WIDTH*2-1+0:0] tmp00_48_16;
	wire [WIDTH*2-1+0:0] tmp00_48_17;
	wire [WIDTH*2-1+0:0] tmp00_48_18;
	wire [WIDTH*2-1+0:0] tmp00_48_19;
	wire [WIDTH*2-1+0:0] tmp00_48_20;
	wire [WIDTH*2-1+0:0] tmp00_48_21;
	wire [WIDTH*2-1+0:0] tmp00_48_22;
	wire [WIDTH*2-1+0:0] tmp00_48_23;
	wire [WIDTH*2-1+0:0] tmp00_48_24;
	wire [WIDTH*2-1+0:0] tmp00_48_25;
	wire [WIDTH*2-1+0:0] tmp00_48_26;
	wire [WIDTH*2-1+0:0] tmp00_48_27;
	wire [WIDTH*2-1+0:0] tmp00_48_28;
	wire [WIDTH*2-1+0:0] tmp00_48_29;
	wire [WIDTH*2-1+0:0] tmp00_48_30;
	wire [WIDTH*2-1+0:0] tmp00_48_31;
	wire [WIDTH*2-1+0:0] tmp00_48_32;
	wire [WIDTH*2-1+0:0] tmp00_48_33;
	wire [WIDTH*2-1+0:0] tmp00_48_34;
	wire [WIDTH*2-1+0:0] tmp00_48_35;
	wire [WIDTH*2-1+0:0] tmp00_48_36;
	wire [WIDTH*2-1+0:0] tmp00_48_37;
	wire [WIDTH*2-1+0:0] tmp00_48_38;
	wire [WIDTH*2-1+0:0] tmp00_48_39;
	wire [WIDTH*2-1+0:0] tmp00_48_40;
	wire [WIDTH*2-1+0:0] tmp00_48_41;
	wire [WIDTH*2-1+0:0] tmp00_48_42;
	wire [WIDTH*2-1+0:0] tmp00_48_43;
	wire [WIDTH*2-1+0:0] tmp00_48_44;
	wire [WIDTH*2-1+0:0] tmp00_48_45;
	wire [WIDTH*2-1+0:0] tmp00_48_46;
	wire [WIDTH*2-1+0:0] tmp00_48_47;
	wire [WIDTH*2-1+0:0] tmp00_48_48;
	wire [WIDTH*2-1+0:0] tmp00_48_49;
	wire [WIDTH*2-1+0:0] tmp00_48_50;
	wire [WIDTH*2-1+0:0] tmp00_48_51;
	wire [WIDTH*2-1+0:0] tmp00_48_52;
	wire [WIDTH*2-1+0:0] tmp00_48_53;
	wire [WIDTH*2-1+0:0] tmp00_48_54;
	wire [WIDTH*2-1+0:0] tmp00_48_55;
	wire [WIDTH*2-1+0:0] tmp00_48_56;
	wire [WIDTH*2-1+0:0] tmp00_48_57;
	wire [WIDTH*2-1+0:0] tmp00_48_58;
	wire [WIDTH*2-1+0:0] tmp00_48_59;
	wire [WIDTH*2-1+0:0] tmp00_48_60;
	wire [WIDTH*2-1+0:0] tmp00_48_61;
	wire [WIDTH*2-1+0:0] tmp00_48_62;
	wire [WIDTH*2-1+0:0] tmp00_48_63;
	wire [WIDTH*2-1+0:0] tmp00_48_64;
	wire [WIDTH*2-1+0:0] tmp00_48_65;
	wire [WIDTH*2-1+0:0] tmp00_48_66;
	wire [WIDTH*2-1+0:0] tmp00_48_67;
	wire [WIDTH*2-1+0:0] tmp00_48_68;
	wire [WIDTH*2-1+0:0] tmp00_48_69;
	wire [WIDTH*2-1+0:0] tmp00_48_70;
	wire [WIDTH*2-1+0:0] tmp00_48_71;
	wire [WIDTH*2-1+0:0] tmp00_48_72;
	wire [WIDTH*2-1+0:0] tmp00_48_73;
	wire [WIDTH*2-1+0:0] tmp00_48_74;
	wire [WIDTH*2-1+0:0] tmp00_48_75;
	wire [WIDTH*2-1+0:0] tmp00_48_76;
	wire [WIDTH*2-1+0:0] tmp00_48_77;
	wire [WIDTH*2-1+0:0] tmp00_48_78;
	wire [WIDTH*2-1+0:0] tmp00_48_79;
	wire [WIDTH*2-1+0:0] tmp00_48_80;
	wire [WIDTH*2-1+0:0] tmp00_48_81;
	wire [WIDTH*2-1+0:0] tmp00_48_82;
	wire [WIDTH*2-1+0:0] tmp00_48_83;
	wire [WIDTH*2-1+0:0] tmp00_49_0;
	wire [WIDTH*2-1+0:0] tmp00_49_1;
	wire [WIDTH*2-1+0:0] tmp00_49_2;
	wire [WIDTH*2-1+0:0] tmp00_49_3;
	wire [WIDTH*2-1+0:0] tmp00_49_4;
	wire [WIDTH*2-1+0:0] tmp00_49_5;
	wire [WIDTH*2-1+0:0] tmp00_49_6;
	wire [WIDTH*2-1+0:0] tmp00_49_7;
	wire [WIDTH*2-1+0:0] tmp00_49_8;
	wire [WIDTH*2-1+0:0] tmp00_49_9;
	wire [WIDTH*2-1+0:0] tmp00_49_10;
	wire [WIDTH*2-1+0:0] tmp00_49_11;
	wire [WIDTH*2-1+0:0] tmp00_49_12;
	wire [WIDTH*2-1+0:0] tmp00_49_13;
	wire [WIDTH*2-1+0:0] tmp00_49_14;
	wire [WIDTH*2-1+0:0] tmp00_49_15;
	wire [WIDTH*2-1+0:0] tmp00_49_16;
	wire [WIDTH*2-1+0:0] tmp00_49_17;
	wire [WIDTH*2-1+0:0] tmp00_49_18;
	wire [WIDTH*2-1+0:0] tmp00_49_19;
	wire [WIDTH*2-1+0:0] tmp00_49_20;
	wire [WIDTH*2-1+0:0] tmp00_49_21;
	wire [WIDTH*2-1+0:0] tmp00_49_22;
	wire [WIDTH*2-1+0:0] tmp00_49_23;
	wire [WIDTH*2-1+0:0] tmp00_49_24;
	wire [WIDTH*2-1+0:0] tmp00_49_25;
	wire [WIDTH*2-1+0:0] tmp00_49_26;
	wire [WIDTH*2-1+0:0] tmp00_49_27;
	wire [WIDTH*2-1+0:0] tmp00_49_28;
	wire [WIDTH*2-1+0:0] tmp00_49_29;
	wire [WIDTH*2-1+0:0] tmp00_49_30;
	wire [WIDTH*2-1+0:0] tmp00_49_31;
	wire [WIDTH*2-1+0:0] tmp00_49_32;
	wire [WIDTH*2-1+0:0] tmp00_49_33;
	wire [WIDTH*2-1+0:0] tmp00_49_34;
	wire [WIDTH*2-1+0:0] tmp00_49_35;
	wire [WIDTH*2-1+0:0] tmp00_49_36;
	wire [WIDTH*2-1+0:0] tmp00_49_37;
	wire [WIDTH*2-1+0:0] tmp00_49_38;
	wire [WIDTH*2-1+0:0] tmp00_49_39;
	wire [WIDTH*2-1+0:0] tmp00_49_40;
	wire [WIDTH*2-1+0:0] tmp00_49_41;
	wire [WIDTH*2-1+0:0] tmp00_49_42;
	wire [WIDTH*2-1+0:0] tmp00_49_43;
	wire [WIDTH*2-1+0:0] tmp00_49_44;
	wire [WIDTH*2-1+0:0] tmp00_49_45;
	wire [WIDTH*2-1+0:0] tmp00_49_46;
	wire [WIDTH*2-1+0:0] tmp00_49_47;
	wire [WIDTH*2-1+0:0] tmp00_49_48;
	wire [WIDTH*2-1+0:0] tmp00_49_49;
	wire [WIDTH*2-1+0:0] tmp00_49_50;
	wire [WIDTH*2-1+0:0] tmp00_49_51;
	wire [WIDTH*2-1+0:0] tmp00_49_52;
	wire [WIDTH*2-1+0:0] tmp00_49_53;
	wire [WIDTH*2-1+0:0] tmp00_49_54;
	wire [WIDTH*2-1+0:0] tmp00_49_55;
	wire [WIDTH*2-1+0:0] tmp00_49_56;
	wire [WIDTH*2-1+0:0] tmp00_49_57;
	wire [WIDTH*2-1+0:0] tmp00_49_58;
	wire [WIDTH*2-1+0:0] tmp00_49_59;
	wire [WIDTH*2-1+0:0] tmp00_49_60;
	wire [WIDTH*2-1+0:0] tmp00_49_61;
	wire [WIDTH*2-1+0:0] tmp00_49_62;
	wire [WIDTH*2-1+0:0] tmp00_49_63;
	wire [WIDTH*2-1+0:0] tmp00_49_64;
	wire [WIDTH*2-1+0:0] tmp00_49_65;
	wire [WIDTH*2-1+0:0] tmp00_49_66;
	wire [WIDTH*2-1+0:0] tmp00_49_67;
	wire [WIDTH*2-1+0:0] tmp00_49_68;
	wire [WIDTH*2-1+0:0] tmp00_49_69;
	wire [WIDTH*2-1+0:0] tmp00_49_70;
	wire [WIDTH*2-1+0:0] tmp00_49_71;
	wire [WIDTH*2-1+0:0] tmp00_49_72;
	wire [WIDTH*2-1+0:0] tmp00_49_73;
	wire [WIDTH*2-1+0:0] tmp00_49_74;
	wire [WIDTH*2-1+0:0] tmp00_49_75;
	wire [WIDTH*2-1+0:0] tmp00_49_76;
	wire [WIDTH*2-1+0:0] tmp00_49_77;
	wire [WIDTH*2-1+0:0] tmp00_49_78;
	wire [WIDTH*2-1+0:0] tmp00_49_79;
	wire [WIDTH*2-1+0:0] tmp00_49_80;
	wire [WIDTH*2-1+0:0] tmp00_49_81;
	wire [WIDTH*2-1+0:0] tmp00_49_82;
	wire [WIDTH*2-1+0:0] tmp00_49_83;
	wire [WIDTH*2-1+0:0] tmp00_50_0;
	wire [WIDTH*2-1+0:0] tmp00_50_1;
	wire [WIDTH*2-1+0:0] tmp00_50_2;
	wire [WIDTH*2-1+0:0] tmp00_50_3;
	wire [WIDTH*2-1+0:0] tmp00_50_4;
	wire [WIDTH*2-1+0:0] tmp00_50_5;
	wire [WIDTH*2-1+0:0] tmp00_50_6;
	wire [WIDTH*2-1+0:0] tmp00_50_7;
	wire [WIDTH*2-1+0:0] tmp00_50_8;
	wire [WIDTH*2-1+0:0] tmp00_50_9;
	wire [WIDTH*2-1+0:0] tmp00_50_10;
	wire [WIDTH*2-1+0:0] tmp00_50_11;
	wire [WIDTH*2-1+0:0] tmp00_50_12;
	wire [WIDTH*2-1+0:0] tmp00_50_13;
	wire [WIDTH*2-1+0:0] tmp00_50_14;
	wire [WIDTH*2-1+0:0] tmp00_50_15;
	wire [WIDTH*2-1+0:0] tmp00_50_16;
	wire [WIDTH*2-1+0:0] tmp00_50_17;
	wire [WIDTH*2-1+0:0] tmp00_50_18;
	wire [WIDTH*2-1+0:0] tmp00_50_19;
	wire [WIDTH*2-1+0:0] tmp00_50_20;
	wire [WIDTH*2-1+0:0] tmp00_50_21;
	wire [WIDTH*2-1+0:0] tmp00_50_22;
	wire [WIDTH*2-1+0:0] tmp00_50_23;
	wire [WIDTH*2-1+0:0] tmp00_50_24;
	wire [WIDTH*2-1+0:0] tmp00_50_25;
	wire [WIDTH*2-1+0:0] tmp00_50_26;
	wire [WIDTH*2-1+0:0] tmp00_50_27;
	wire [WIDTH*2-1+0:0] tmp00_50_28;
	wire [WIDTH*2-1+0:0] tmp00_50_29;
	wire [WIDTH*2-1+0:0] tmp00_50_30;
	wire [WIDTH*2-1+0:0] tmp00_50_31;
	wire [WIDTH*2-1+0:0] tmp00_50_32;
	wire [WIDTH*2-1+0:0] tmp00_50_33;
	wire [WIDTH*2-1+0:0] tmp00_50_34;
	wire [WIDTH*2-1+0:0] tmp00_50_35;
	wire [WIDTH*2-1+0:0] tmp00_50_36;
	wire [WIDTH*2-1+0:0] tmp00_50_37;
	wire [WIDTH*2-1+0:0] tmp00_50_38;
	wire [WIDTH*2-1+0:0] tmp00_50_39;
	wire [WIDTH*2-1+0:0] tmp00_50_40;
	wire [WIDTH*2-1+0:0] tmp00_50_41;
	wire [WIDTH*2-1+0:0] tmp00_50_42;
	wire [WIDTH*2-1+0:0] tmp00_50_43;
	wire [WIDTH*2-1+0:0] tmp00_50_44;
	wire [WIDTH*2-1+0:0] tmp00_50_45;
	wire [WIDTH*2-1+0:0] tmp00_50_46;
	wire [WIDTH*2-1+0:0] tmp00_50_47;
	wire [WIDTH*2-1+0:0] tmp00_50_48;
	wire [WIDTH*2-1+0:0] tmp00_50_49;
	wire [WIDTH*2-1+0:0] tmp00_50_50;
	wire [WIDTH*2-1+0:0] tmp00_50_51;
	wire [WIDTH*2-1+0:0] tmp00_50_52;
	wire [WIDTH*2-1+0:0] tmp00_50_53;
	wire [WIDTH*2-1+0:0] tmp00_50_54;
	wire [WIDTH*2-1+0:0] tmp00_50_55;
	wire [WIDTH*2-1+0:0] tmp00_50_56;
	wire [WIDTH*2-1+0:0] tmp00_50_57;
	wire [WIDTH*2-1+0:0] tmp00_50_58;
	wire [WIDTH*2-1+0:0] tmp00_50_59;
	wire [WIDTH*2-1+0:0] tmp00_50_60;
	wire [WIDTH*2-1+0:0] tmp00_50_61;
	wire [WIDTH*2-1+0:0] tmp00_50_62;
	wire [WIDTH*2-1+0:0] tmp00_50_63;
	wire [WIDTH*2-1+0:0] tmp00_50_64;
	wire [WIDTH*2-1+0:0] tmp00_50_65;
	wire [WIDTH*2-1+0:0] tmp00_50_66;
	wire [WIDTH*2-1+0:0] tmp00_50_67;
	wire [WIDTH*2-1+0:0] tmp00_50_68;
	wire [WIDTH*2-1+0:0] tmp00_50_69;
	wire [WIDTH*2-1+0:0] tmp00_50_70;
	wire [WIDTH*2-1+0:0] tmp00_50_71;
	wire [WIDTH*2-1+0:0] tmp00_50_72;
	wire [WIDTH*2-1+0:0] tmp00_50_73;
	wire [WIDTH*2-1+0:0] tmp00_50_74;
	wire [WIDTH*2-1+0:0] tmp00_50_75;
	wire [WIDTH*2-1+0:0] tmp00_50_76;
	wire [WIDTH*2-1+0:0] tmp00_50_77;
	wire [WIDTH*2-1+0:0] tmp00_50_78;
	wire [WIDTH*2-1+0:0] tmp00_50_79;
	wire [WIDTH*2-1+0:0] tmp00_50_80;
	wire [WIDTH*2-1+0:0] tmp00_50_81;
	wire [WIDTH*2-1+0:0] tmp00_50_82;
	wire [WIDTH*2-1+0:0] tmp00_50_83;
	wire [WIDTH*2-1+0:0] tmp00_51_0;
	wire [WIDTH*2-1+0:0] tmp00_51_1;
	wire [WIDTH*2-1+0:0] tmp00_51_2;
	wire [WIDTH*2-1+0:0] tmp00_51_3;
	wire [WIDTH*2-1+0:0] tmp00_51_4;
	wire [WIDTH*2-1+0:0] tmp00_51_5;
	wire [WIDTH*2-1+0:0] tmp00_51_6;
	wire [WIDTH*2-1+0:0] tmp00_51_7;
	wire [WIDTH*2-1+0:0] tmp00_51_8;
	wire [WIDTH*2-1+0:0] tmp00_51_9;
	wire [WIDTH*2-1+0:0] tmp00_51_10;
	wire [WIDTH*2-1+0:0] tmp00_51_11;
	wire [WIDTH*2-1+0:0] tmp00_51_12;
	wire [WIDTH*2-1+0:0] tmp00_51_13;
	wire [WIDTH*2-1+0:0] tmp00_51_14;
	wire [WIDTH*2-1+0:0] tmp00_51_15;
	wire [WIDTH*2-1+0:0] tmp00_51_16;
	wire [WIDTH*2-1+0:0] tmp00_51_17;
	wire [WIDTH*2-1+0:0] tmp00_51_18;
	wire [WIDTH*2-1+0:0] tmp00_51_19;
	wire [WIDTH*2-1+0:0] tmp00_51_20;
	wire [WIDTH*2-1+0:0] tmp00_51_21;
	wire [WIDTH*2-1+0:0] tmp00_51_22;
	wire [WIDTH*2-1+0:0] tmp00_51_23;
	wire [WIDTH*2-1+0:0] tmp00_51_24;
	wire [WIDTH*2-1+0:0] tmp00_51_25;
	wire [WIDTH*2-1+0:0] tmp00_51_26;
	wire [WIDTH*2-1+0:0] tmp00_51_27;
	wire [WIDTH*2-1+0:0] tmp00_51_28;
	wire [WIDTH*2-1+0:0] tmp00_51_29;
	wire [WIDTH*2-1+0:0] tmp00_51_30;
	wire [WIDTH*2-1+0:0] tmp00_51_31;
	wire [WIDTH*2-1+0:0] tmp00_51_32;
	wire [WIDTH*2-1+0:0] tmp00_51_33;
	wire [WIDTH*2-1+0:0] tmp00_51_34;
	wire [WIDTH*2-1+0:0] tmp00_51_35;
	wire [WIDTH*2-1+0:0] tmp00_51_36;
	wire [WIDTH*2-1+0:0] tmp00_51_37;
	wire [WIDTH*2-1+0:0] tmp00_51_38;
	wire [WIDTH*2-1+0:0] tmp00_51_39;
	wire [WIDTH*2-1+0:0] tmp00_51_40;
	wire [WIDTH*2-1+0:0] tmp00_51_41;
	wire [WIDTH*2-1+0:0] tmp00_51_42;
	wire [WIDTH*2-1+0:0] tmp00_51_43;
	wire [WIDTH*2-1+0:0] tmp00_51_44;
	wire [WIDTH*2-1+0:0] tmp00_51_45;
	wire [WIDTH*2-1+0:0] tmp00_51_46;
	wire [WIDTH*2-1+0:0] tmp00_51_47;
	wire [WIDTH*2-1+0:0] tmp00_51_48;
	wire [WIDTH*2-1+0:0] tmp00_51_49;
	wire [WIDTH*2-1+0:0] tmp00_51_50;
	wire [WIDTH*2-1+0:0] tmp00_51_51;
	wire [WIDTH*2-1+0:0] tmp00_51_52;
	wire [WIDTH*2-1+0:0] tmp00_51_53;
	wire [WIDTH*2-1+0:0] tmp00_51_54;
	wire [WIDTH*2-1+0:0] tmp00_51_55;
	wire [WIDTH*2-1+0:0] tmp00_51_56;
	wire [WIDTH*2-1+0:0] tmp00_51_57;
	wire [WIDTH*2-1+0:0] tmp00_51_58;
	wire [WIDTH*2-1+0:0] tmp00_51_59;
	wire [WIDTH*2-1+0:0] tmp00_51_60;
	wire [WIDTH*2-1+0:0] tmp00_51_61;
	wire [WIDTH*2-1+0:0] tmp00_51_62;
	wire [WIDTH*2-1+0:0] tmp00_51_63;
	wire [WIDTH*2-1+0:0] tmp00_51_64;
	wire [WIDTH*2-1+0:0] tmp00_51_65;
	wire [WIDTH*2-1+0:0] tmp00_51_66;
	wire [WIDTH*2-1+0:0] tmp00_51_67;
	wire [WIDTH*2-1+0:0] tmp00_51_68;
	wire [WIDTH*2-1+0:0] tmp00_51_69;
	wire [WIDTH*2-1+0:0] tmp00_51_70;
	wire [WIDTH*2-1+0:0] tmp00_51_71;
	wire [WIDTH*2-1+0:0] tmp00_51_72;
	wire [WIDTH*2-1+0:0] tmp00_51_73;
	wire [WIDTH*2-1+0:0] tmp00_51_74;
	wire [WIDTH*2-1+0:0] tmp00_51_75;
	wire [WIDTH*2-1+0:0] tmp00_51_76;
	wire [WIDTH*2-1+0:0] tmp00_51_77;
	wire [WIDTH*2-1+0:0] tmp00_51_78;
	wire [WIDTH*2-1+0:0] tmp00_51_79;
	wire [WIDTH*2-1+0:0] tmp00_51_80;
	wire [WIDTH*2-1+0:0] tmp00_51_81;
	wire [WIDTH*2-1+0:0] tmp00_51_82;
	wire [WIDTH*2-1+0:0] tmp00_51_83;
	wire [WIDTH*2-1+0:0] tmp00_52_0;
	wire [WIDTH*2-1+0:0] tmp00_52_1;
	wire [WIDTH*2-1+0:0] tmp00_52_2;
	wire [WIDTH*2-1+0:0] tmp00_52_3;
	wire [WIDTH*2-1+0:0] tmp00_52_4;
	wire [WIDTH*2-1+0:0] tmp00_52_5;
	wire [WIDTH*2-1+0:0] tmp00_52_6;
	wire [WIDTH*2-1+0:0] tmp00_52_7;
	wire [WIDTH*2-1+0:0] tmp00_52_8;
	wire [WIDTH*2-1+0:0] tmp00_52_9;
	wire [WIDTH*2-1+0:0] tmp00_52_10;
	wire [WIDTH*2-1+0:0] tmp00_52_11;
	wire [WIDTH*2-1+0:0] tmp00_52_12;
	wire [WIDTH*2-1+0:0] tmp00_52_13;
	wire [WIDTH*2-1+0:0] tmp00_52_14;
	wire [WIDTH*2-1+0:0] tmp00_52_15;
	wire [WIDTH*2-1+0:0] tmp00_52_16;
	wire [WIDTH*2-1+0:0] tmp00_52_17;
	wire [WIDTH*2-1+0:0] tmp00_52_18;
	wire [WIDTH*2-1+0:0] tmp00_52_19;
	wire [WIDTH*2-1+0:0] tmp00_52_20;
	wire [WIDTH*2-1+0:0] tmp00_52_21;
	wire [WIDTH*2-1+0:0] tmp00_52_22;
	wire [WIDTH*2-1+0:0] tmp00_52_23;
	wire [WIDTH*2-1+0:0] tmp00_52_24;
	wire [WIDTH*2-1+0:0] tmp00_52_25;
	wire [WIDTH*2-1+0:0] tmp00_52_26;
	wire [WIDTH*2-1+0:0] tmp00_52_27;
	wire [WIDTH*2-1+0:0] tmp00_52_28;
	wire [WIDTH*2-1+0:0] tmp00_52_29;
	wire [WIDTH*2-1+0:0] tmp00_52_30;
	wire [WIDTH*2-1+0:0] tmp00_52_31;
	wire [WIDTH*2-1+0:0] tmp00_52_32;
	wire [WIDTH*2-1+0:0] tmp00_52_33;
	wire [WIDTH*2-1+0:0] tmp00_52_34;
	wire [WIDTH*2-1+0:0] tmp00_52_35;
	wire [WIDTH*2-1+0:0] tmp00_52_36;
	wire [WIDTH*2-1+0:0] tmp00_52_37;
	wire [WIDTH*2-1+0:0] tmp00_52_38;
	wire [WIDTH*2-1+0:0] tmp00_52_39;
	wire [WIDTH*2-1+0:0] tmp00_52_40;
	wire [WIDTH*2-1+0:0] tmp00_52_41;
	wire [WIDTH*2-1+0:0] tmp00_52_42;
	wire [WIDTH*2-1+0:0] tmp00_52_43;
	wire [WIDTH*2-1+0:0] tmp00_52_44;
	wire [WIDTH*2-1+0:0] tmp00_52_45;
	wire [WIDTH*2-1+0:0] tmp00_52_46;
	wire [WIDTH*2-1+0:0] tmp00_52_47;
	wire [WIDTH*2-1+0:0] tmp00_52_48;
	wire [WIDTH*2-1+0:0] tmp00_52_49;
	wire [WIDTH*2-1+0:0] tmp00_52_50;
	wire [WIDTH*2-1+0:0] tmp00_52_51;
	wire [WIDTH*2-1+0:0] tmp00_52_52;
	wire [WIDTH*2-1+0:0] tmp00_52_53;
	wire [WIDTH*2-1+0:0] tmp00_52_54;
	wire [WIDTH*2-1+0:0] tmp00_52_55;
	wire [WIDTH*2-1+0:0] tmp00_52_56;
	wire [WIDTH*2-1+0:0] tmp00_52_57;
	wire [WIDTH*2-1+0:0] tmp00_52_58;
	wire [WIDTH*2-1+0:0] tmp00_52_59;
	wire [WIDTH*2-1+0:0] tmp00_52_60;
	wire [WIDTH*2-1+0:0] tmp00_52_61;
	wire [WIDTH*2-1+0:0] tmp00_52_62;
	wire [WIDTH*2-1+0:0] tmp00_52_63;
	wire [WIDTH*2-1+0:0] tmp00_52_64;
	wire [WIDTH*2-1+0:0] tmp00_52_65;
	wire [WIDTH*2-1+0:0] tmp00_52_66;
	wire [WIDTH*2-1+0:0] tmp00_52_67;
	wire [WIDTH*2-1+0:0] tmp00_52_68;
	wire [WIDTH*2-1+0:0] tmp00_52_69;
	wire [WIDTH*2-1+0:0] tmp00_52_70;
	wire [WIDTH*2-1+0:0] tmp00_52_71;
	wire [WIDTH*2-1+0:0] tmp00_52_72;
	wire [WIDTH*2-1+0:0] tmp00_52_73;
	wire [WIDTH*2-1+0:0] tmp00_52_74;
	wire [WIDTH*2-1+0:0] tmp00_52_75;
	wire [WIDTH*2-1+0:0] tmp00_52_76;
	wire [WIDTH*2-1+0:0] tmp00_52_77;
	wire [WIDTH*2-1+0:0] tmp00_52_78;
	wire [WIDTH*2-1+0:0] tmp00_52_79;
	wire [WIDTH*2-1+0:0] tmp00_52_80;
	wire [WIDTH*2-1+0:0] tmp00_52_81;
	wire [WIDTH*2-1+0:0] tmp00_52_82;
	wire [WIDTH*2-1+0:0] tmp00_52_83;
	wire [WIDTH*2-1+0:0] tmp00_53_0;
	wire [WIDTH*2-1+0:0] tmp00_53_1;
	wire [WIDTH*2-1+0:0] tmp00_53_2;
	wire [WIDTH*2-1+0:0] tmp00_53_3;
	wire [WIDTH*2-1+0:0] tmp00_53_4;
	wire [WIDTH*2-1+0:0] tmp00_53_5;
	wire [WIDTH*2-1+0:0] tmp00_53_6;
	wire [WIDTH*2-1+0:0] tmp00_53_7;
	wire [WIDTH*2-1+0:0] tmp00_53_8;
	wire [WIDTH*2-1+0:0] tmp00_53_9;
	wire [WIDTH*2-1+0:0] tmp00_53_10;
	wire [WIDTH*2-1+0:0] tmp00_53_11;
	wire [WIDTH*2-1+0:0] tmp00_53_12;
	wire [WIDTH*2-1+0:0] tmp00_53_13;
	wire [WIDTH*2-1+0:0] tmp00_53_14;
	wire [WIDTH*2-1+0:0] tmp00_53_15;
	wire [WIDTH*2-1+0:0] tmp00_53_16;
	wire [WIDTH*2-1+0:0] tmp00_53_17;
	wire [WIDTH*2-1+0:0] tmp00_53_18;
	wire [WIDTH*2-1+0:0] tmp00_53_19;
	wire [WIDTH*2-1+0:0] tmp00_53_20;
	wire [WIDTH*2-1+0:0] tmp00_53_21;
	wire [WIDTH*2-1+0:0] tmp00_53_22;
	wire [WIDTH*2-1+0:0] tmp00_53_23;
	wire [WIDTH*2-1+0:0] tmp00_53_24;
	wire [WIDTH*2-1+0:0] tmp00_53_25;
	wire [WIDTH*2-1+0:0] tmp00_53_26;
	wire [WIDTH*2-1+0:0] tmp00_53_27;
	wire [WIDTH*2-1+0:0] tmp00_53_28;
	wire [WIDTH*2-1+0:0] tmp00_53_29;
	wire [WIDTH*2-1+0:0] tmp00_53_30;
	wire [WIDTH*2-1+0:0] tmp00_53_31;
	wire [WIDTH*2-1+0:0] tmp00_53_32;
	wire [WIDTH*2-1+0:0] tmp00_53_33;
	wire [WIDTH*2-1+0:0] tmp00_53_34;
	wire [WIDTH*2-1+0:0] tmp00_53_35;
	wire [WIDTH*2-1+0:0] tmp00_53_36;
	wire [WIDTH*2-1+0:0] tmp00_53_37;
	wire [WIDTH*2-1+0:0] tmp00_53_38;
	wire [WIDTH*2-1+0:0] tmp00_53_39;
	wire [WIDTH*2-1+0:0] tmp00_53_40;
	wire [WIDTH*2-1+0:0] tmp00_53_41;
	wire [WIDTH*2-1+0:0] tmp00_53_42;
	wire [WIDTH*2-1+0:0] tmp00_53_43;
	wire [WIDTH*2-1+0:0] tmp00_53_44;
	wire [WIDTH*2-1+0:0] tmp00_53_45;
	wire [WIDTH*2-1+0:0] tmp00_53_46;
	wire [WIDTH*2-1+0:0] tmp00_53_47;
	wire [WIDTH*2-1+0:0] tmp00_53_48;
	wire [WIDTH*2-1+0:0] tmp00_53_49;
	wire [WIDTH*2-1+0:0] tmp00_53_50;
	wire [WIDTH*2-1+0:0] tmp00_53_51;
	wire [WIDTH*2-1+0:0] tmp00_53_52;
	wire [WIDTH*2-1+0:0] tmp00_53_53;
	wire [WIDTH*2-1+0:0] tmp00_53_54;
	wire [WIDTH*2-1+0:0] tmp00_53_55;
	wire [WIDTH*2-1+0:0] tmp00_53_56;
	wire [WIDTH*2-1+0:0] tmp00_53_57;
	wire [WIDTH*2-1+0:0] tmp00_53_58;
	wire [WIDTH*2-1+0:0] tmp00_53_59;
	wire [WIDTH*2-1+0:0] tmp00_53_60;
	wire [WIDTH*2-1+0:0] tmp00_53_61;
	wire [WIDTH*2-1+0:0] tmp00_53_62;
	wire [WIDTH*2-1+0:0] tmp00_53_63;
	wire [WIDTH*2-1+0:0] tmp00_53_64;
	wire [WIDTH*2-1+0:0] tmp00_53_65;
	wire [WIDTH*2-1+0:0] tmp00_53_66;
	wire [WIDTH*2-1+0:0] tmp00_53_67;
	wire [WIDTH*2-1+0:0] tmp00_53_68;
	wire [WIDTH*2-1+0:0] tmp00_53_69;
	wire [WIDTH*2-1+0:0] tmp00_53_70;
	wire [WIDTH*2-1+0:0] tmp00_53_71;
	wire [WIDTH*2-1+0:0] tmp00_53_72;
	wire [WIDTH*2-1+0:0] tmp00_53_73;
	wire [WIDTH*2-1+0:0] tmp00_53_74;
	wire [WIDTH*2-1+0:0] tmp00_53_75;
	wire [WIDTH*2-1+0:0] tmp00_53_76;
	wire [WIDTH*2-1+0:0] tmp00_53_77;
	wire [WIDTH*2-1+0:0] tmp00_53_78;
	wire [WIDTH*2-1+0:0] tmp00_53_79;
	wire [WIDTH*2-1+0:0] tmp00_53_80;
	wire [WIDTH*2-1+0:0] tmp00_53_81;
	wire [WIDTH*2-1+0:0] tmp00_53_82;
	wire [WIDTH*2-1+0:0] tmp00_53_83;
	wire [WIDTH*2-1+0:0] tmp00_54_0;
	wire [WIDTH*2-1+0:0] tmp00_54_1;
	wire [WIDTH*2-1+0:0] tmp00_54_2;
	wire [WIDTH*2-1+0:0] tmp00_54_3;
	wire [WIDTH*2-1+0:0] tmp00_54_4;
	wire [WIDTH*2-1+0:0] tmp00_54_5;
	wire [WIDTH*2-1+0:0] tmp00_54_6;
	wire [WIDTH*2-1+0:0] tmp00_54_7;
	wire [WIDTH*2-1+0:0] tmp00_54_8;
	wire [WIDTH*2-1+0:0] tmp00_54_9;
	wire [WIDTH*2-1+0:0] tmp00_54_10;
	wire [WIDTH*2-1+0:0] tmp00_54_11;
	wire [WIDTH*2-1+0:0] tmp00_54_12;
	wire [WIDTH*2-1+0:0] tmp00_54_13;
	wire [WIDTH*2-1+0:0] tmp00_54_14;
	wire [WIDTH*2-1+0:0] tmp00_54_15;
	wire [WIDTH*2-1+0:0] tmp00_54_16;
	wire [WIDTH*2-1+0:0] tmp00_54_17;
	wire [WIDTH*2-1+0:0] tmp00_54_18;
	wire [WIDTH*2-1+0:0] tmp00_54_19;
	wire [WIDTH*2-1+0:0] tmp00_54_20;
	wire [WIDTH*2-1+0:0] tmp00_54_21;
	wire [WIDTH*2-1+0:0] tmp00_54_22;
	wire [WIDTH*2-1+0:0] tmp00_54_23;
	wire [WIDTH*2-1+0:0] tmp00_54_24;
	wire [WIDTH*2-1+0:0] tmp00_54_25;
	wire [WIDTH*2-1+0:0] tmp00_54_26;
	wire [WIDTH*2-1+0:0] tmp00_54_27;
	wire [WIDTH*2-1+0:0] tmp00_54_28;
	wire [WIDTH*2-1+0:0] tmp00_54_29;
	wire [WIDTH*2-1+0:0] tmp00_54_30;
	wire [WIDTH*2-1+0:0] tmp00_54_31;
	wire [WIDTH*2-1+0:0] tmp00_54_32;
	wire [WIDTH*2-1+0:0] tmp00_54_33;
	wire [WIDTH*2-1+0:0] tmp00_54_34;
	wire [WIDTH*2-1+0:0] tmp00_54_35;
	wire [WIDTH*2-1+0:0] tmp00_54_36;
	wire [WIDTH*2-1+0:0] tmp00_54_37;
	wire [WIDTH*2-1+0:0] tmp00_54_38;
	wire [WIDTH*2-1+0:0] tmp00_54_39;
	wire [WIDTH*2-1+0:0] tmp00_54_40;
	wire [WIDTH*2-1+0:0] tmp00_54_41;
	wire [WIDTH*2-1+0:0] tmp00_54_42;
	wire [WIDTH*2-1+0:0] tmp00_54_43;
	wire [WIDTH*2-1+0:0] tmp00_54_44;
	wire [WIDTH*2-1+0:0] tmp00_54_45;
	wire [WIDTH*2-1+0:0] tmp00_54_46;
	wire [WIDTH*2-1+0:0] tmp00_54_47;
	wire [WIDTH*2-1+0:0] tmp00_54_48;
	wire [WIDTH*2-1+0:0] tmp00_54_49;
	wire [WIDTH*2-1+0:0] tmp00_54_50;
	wire [WIDTH*2-1+0:0] tmp00_54_51;
	wire [WIDTH*2-1+0:0] tmp00_54_52;
	wire [WIDTH*2-1+0:0] tmp00_54_53;
	wire [WIDTH*2-1+0:0] tmp00_54_54;
	wire [WIDTH*2-1+0:0] tmp00_54_55;
	wire [WIDTH*2-1+0:0] tmp00_54_56;
	wire [WIDTH*2-1+0:0] tmp00_54_57;
	wire [WIDTH*2-1+0:0] tmp00_54_58;
	wire [WIDTH*2-1+0:0] tmp00_54_59;
	wire [WIDTH*2-1+0:0] tmp00_54_60;
	wire [WIDTH*2-1+0:0] tmp00_54_61;
	wire [WIDTH*2-1+0:0] tmp00_54_62;
	wire [WIDTH*2-1+0:0] tmp00_54_63;
	wire [WIDTH*2-1+0:0] tmp00_54_64;
	wire [WIDTH*2-1+0:0] tmp00_54_65;
	wire [WIDTH*2-1+0:0] tmp00_54_66;
	wire [WIDTH*2-1+0:0] tmp00_54_67;
	wire [WIDTH*2-1+0:0] tmp00_54_68;
	wire [WIDTH*2-1+0:0] tmp00_54_69;
	wire [WIDTH*2-1+0:0] tmp00_54_70;
	wire [WIDTH*2-1+0:0] tmp00_54_71;
	wire [WIDTH*2-1+0:0] tmp00_54_72;
	wire [WIDTH*2-1+0:0] tmp00_54_73;
	wire [WIDTH*2-1+0:0] tmp00_54_74;
	wire [WIDTH*2-1+0:0] tmp00_54_75;
	wire [WIDTH*2-1+0:0] tmp00_54_76;
	wire [WIDTH*2-1+0:0] tmp00_54_77;
	wire [WIDTH*2-1+0:0] tmp00_54_78;
	wire [WIDTH*2-1+0:0] tmp00_54_79;
	wire [WIDTH*2-1+0:0] tmp00_54_80;
	wire [WIDTH*2-1+0:0] tmp00_54_81;
	wire [WIDTH*2-1+0:0] tmp00_54_82;
	wire [WIDTH*2-1+0:0] tmp00_54_83;
	wire [WIDTH*2-1+0:0] tmp00_55_0;
	wire [WIDTH*2-1+0:0] tmp00_55_1;
	wire [WIDTH*2-1+0:0] tmp00_55_2;
	wire [WIDTH*2-1+0:0] tmp00_55_3;
	wire [WIDTH*2-1+0:0] tmp00_55_4;
	wire [WIDTH*2-1+0:0] tmp00_55_5;
	wire [WIDTH*2-1+0:0] tmp00_55_6;
	wire [WIDTH*2-1+0:0] tmp00_55_7;
	wire [WIDTH*2-1+0:0] tmp00_55_8;
	wire [WIDTH*2-1+0:0] tmp00_55_9;
	wire [WIDTH*2-1+0:0] tmp00_55_10;
	wire [WIDTH*2-1+0:0] tmp00_55_11;
	wire [WIDTH*2-1+0:0] tmp00_55_12;
	wire [WIDTH*2-1+0:0] tmp00_55_13;
	wire [WIDTH*2-1+0:0] tmp00_55_14;
	wire [WIDTH*2-1+0:0] tmp00_55_15;
	wire [WIDTH*2-1+0:0] tmp00_55_16;
	wire [WIDTH*2-1+0:0] tmp00_55_17;
	wire [WIDTH*2-1+0:0] tmp00_55_18;
	wire [WIDTH*2-1+0:0] tmp00_55_19;
	wire [WIDTH*2-1+0:0] tmp00_55_20;
	wire [WIDTH*2-1+0:0] tmp00_55_21;
	wire [WIDTH*2-1+0:0] tmp00_55_22;
	wire [WIDTH*2-1+0:0] tmp00_55_23;
	wire [WIDTH*2-1+0:0] tmp00_55_24;
	wire [WIDTH*2-1+0:0] tmp00_55_25;
	wire [WIDTH*2-1+0:0] tmp00_55_26;
	wire [WIDTH*2-1+0:0] tmp00_55_27;
	wire [WIDTH*2-1+0:0] tmp00_55_28;
	wire [WIDTH*2-1+0:0] tmp00_55_29;
	wire [WIDTH*2-1+0:0] tmp00_55_30;
	wire [WIDTH*2-1+0:0] tmp00_55_31;
	wire [WIDTH*2-1+0:0] tmp00_55_32;
	wire [WIDTH*2-1+0:0] tmp00_55_33;
	wire [WIDTH*2-1+0:0] tmp00_55_34;
	wire [WIDTH*2-1+0:0] tmp00_55_35;
	wire [WIDTH*2-1+0:0] tmp00_55_36;
	wire [WIDTH*2-1+0:0] tmp00_55_37;
	wire [WIDTH*2-1+0:0] tmp00_55_38;
	wire [WIDTH*2-1+0:0] tmp00_55_39;
	wire [WIDTH*2-1+0:0] tmp00_55_40;
	wire [WIDTH*2-1+0:0] tmp00_55_41;
	wire [WIDTH*2-1+0:0] tmp00_55_42;
	wire [WIDTH*2-1+0:0] tmp00_55_43;
	wire [WIDTH*2-1+0:0] tmp00_55_44;
	wire [WIDTH*2-1+0:0] tmp00_55_45;
	wire [WIDTH*2-1+0:0] tmp00_55_46;
	wire [WIDTH*2-1+0:0] tmp00_55_47;
	wire [WIDTH*2-1+0:0] tmp00_55_48;
	wire [WIDTH*2-1+0:0] tmp00_55_49;
	wire [WIDTH*2-1+0:0] tmp00_55_50;
	wire [WIDTH*2-1+0:0] tmp00_55_51;
	wire [WIDTH*2-1+0:0] tmp00_55_52;
	wire [WIDTH*2-1+0:0] tmp00_55_53;
	wire [WIDTH*2-1+0:0] tmp00_55_54;
	wire [WIDTH*2-1+0:0] tmp00_55_55;
	wire [WIDTH*2-1+0:0] tmp00_55_56;
	wire [WIDTH*2-1+0:0] tmp00_55_57;
	wire [WIDTH*2-1+0:0] tmp00_55_58;
	wire [WIDTH*2-1+0:0] tmp00_55_59;
	wire [WIDTH*2-1+0:0] tmp00_55_60;
	wire [WIDTH*2-1+0:0] tmp00_55_61;
	wire [WIDTH*2-1+0:0] tmp00_55_62;
	wire [WIDTH*2-1+0:0] tmp00_55_63;
	wire [WIDTH*2-1+0:0] tmp00_55_64;
	wire [WIDTH*2-1+0:0] tmp00_55_65;
	wire [WIDTH*2-1+0:0] tmp00_55_66;
	wire [WIDTH*2-1+0:0] tmp00_55_67;
	wire [WIDTH*2-1+0:0] tmp00_55_68;
	wire [WIDTH*2-1+0:0] tmp00_55_69;
	wire [WIDTH*2-1+0:0] tmp00_55_70;
	wire [WIDTH*2-1+0:0] tmp00_55_71;
	wire [WIDTH*2-1+0:0] tmp00_55_72;
	wire [WIDTH*2-1+0:0] tmp00_55_73;
	wire [WIDTH*2-1+0:0] tmp00_55_74;
	wire [WIDTH*2-1+0:0] tmp00_55_75;
	wire [WIDTH*2-1+0:0] tmp00_55_76;
	wire [WIDTH*2-1+0:0] tmp00_55_77;
	wire [WIDTH*2-1+0:0] tmp00_55_78;
	wire [WIDTH*2-1+0:0] tmp00_55_79;
	wire [WIDTH*2-1+0:0] tmp00_55_80;
	wire [WIDTH*2-1+0:0] tmp00_55_81;
	wire [WIDTH*2-1+0:0] tmp00_55_82;
	wire [WIDTH*2-1+0:0] tmp00_55_83;
	wire [WIDTH*2-1+0:0] tmp00_56_0;
	wire [WIDTH*2-1+0:0] tmp00_56_1;
	wire [WIDTH*2-1+0:0] tmp00_56_2;
	wire [WIDTH*2-1+0:0] tmp00_56_3;
	wire [WIDTH*2-1+0:0] tmp00_56_4;
	wire [WIDTH*2-1+0:0] tmp00_56_5;
	wire [WIDTH*2-1+0:0] tmp00_56_6;
	wire [WIDTH*2-1+0:0] tmp00_56_7;
	wire [WIDTH*2-1+0:0] tmp00_56_8;
	wire [WIDTH*2-1+0:0] tmp00_56_9;
	wire [WIDTH*2-1+0:0] tmp00_56_10;
	wire [WIDTH*2-1+0:0] tmp00_56_11;
	wire [WIDTH*2-1+0:0] tmp00_56_12;
	wire [WIDTH*2-1+0:0] tmp00_56_13;
	wire [WIDTH*2-1+0:0] tmp00_56_14;
	wire [WIDTH*2-1+0:0] tmp00_56_15;
	wire [WIDTH*2-1+0:0] tmp00_56_16;
	wire [WIDTH*2-1+0:0] tmp00_56_17;
	wire [WIDTH*2-1+0:0] tmp00_56_18;
	wire [WIDTH*2-1+0:0] tmp00_56_19;
	wire [WIDTH*2-1+0:0] tmp00_56_20;
	wire [WIDTH*2-1+0:0] tmp00_56_21;
	wire [WIDTH*2-1+0:0] tmp00_56_22;
	wire [WIDTH*2-1+0:0] tmp00_56_23;
	wire [WIDTH*2-1+0:0] tmp00_56_24;
	wire [WIDTH*2-1+0:0] tmp00_56_25;
	wire [WIDTH*2-1+0:0] tmp00_56_26;
	wire [WIDTH*2-1+0:0] tmp00_56_27;
	wire [WIDTH*2-1+0:0] tmp00_56_28;
	wire [WIDTH*2-1+0:0] tmp00_56_29;
	wire [WIDTH*2-1+0:0] tmp00_56_30;
	wire [WIDTH*2-1+0:0] tmp00_56_31;
	wire [WIDTH*2-1+0:0] tmp00_56_32;
	wire [WIDTH*2-1+0:0] tmp00_56_33;
	wire [WIDTH*2-1+0:0] tmp00_56_34;
	wire [WIDTH*2-1+0:0] tmp00_56_35;
	wire [WIDTH*2-1+0:0] tmp00_56_36;
	wire [WIDTH*2-1+0:0] tmp00_56_37;
	wire [WIDTH*2-1+0:0] tmp00_56_38;
	wire [WIDTH*2-1+0:0] tmp00_56_39;
	wire [WIDTH*2-1+0:0] tmp00_56_40;
	wire [WIDTH*2-1+0:0] tmp00_56_41;
	wire [WIDTH*2-1+0:0] tmp00_56_42;
	wire [WIDTH*2-1+0:0] tmp00_56_43;
	wire [WIDTH*2-1+0:0] tmp00_56_44;
	wire [WIDTH*2-1+0:0] tmp00_56_45;
	wire [WIDTH*2-1+0:0] tmp00_56_46;
	wire [WIDTH*2-1+0:0] tmp00_56_47;
	wire [WIDTH*2-1+0:0] tmp00_56_48;
	wire [WIDTH*2-1+0:0] tmp00_56_49;
	wire [WIDTH*2-1+0:0] tmp00_56_50;
	wire [WIDTH*2-1+0:0] tmp00_56_51;
	wire [WIDTH*2-1+0:0] tmp00_56_52;
	wire [WIDTH*2-1+0:0] tmp00_56_53;
	wire [WIDTH*2-1+0:0] tmp00_56_54;
	wire [WIDTH*2-1+0:0] tmp00_56_55;
	wire [WIDTH*2-1+0:0] tmp00_56_56;
	wire [WIDTH*2-1+0:0] tmp00_56_57;
	wire [WIDTH*2-1+0:0] tmp00_56_58;
	wire [WIDTH*2-1+0:0] tmp00_56_59;
	wire [WIDTH*2-1+0:0] tmp00_56_60;
	wire [WIDTH*2-1+0:0] tmp00_56_61;
	wire [WIDTH*2-1+0:0] tmp00_56_62;
	wire [WIDTH*2-1+0:0] tmp00_56_63;
	wire [WIDTH*2-1+0:0] tmp00_56_64;
	wire [WIDTH*2-1+0:0] tmp00_56_65;
	wire [WIDTH*2-1+0:0] tmp00_56_66;
	wire [WIDTH*2-1+0:0] tmp00_56_67;
	wire [WIDTH*2-1+0:0] tmp00_56_68;
	wire [WIDTH*2-1+0:0] tmp00_56_69;
	wire [WIDTH*2-1+0:0] tmp00_56_70;
	wire [WIDTH*2-1+0:0] tmp00_56_71;
	wire [WIDTH*2-1+0:0] tmp00_56_72;
	wire [WIDTH*2-1+0:0] tmp00_56_73;
	wire [WIDTH*2-1+0:0] tmp00_56_74;
	wire [WIDTH*2-1+0:0] tmp00_56_75;
	wire [WIDTH*2-1+0:0] tmp00_56_76;
	wire [WIDTH*2-1+0:0] tmp00_56_77;
	wire [WIDTH*2-1+0:0] tmp00_56_78;
	wire [WIDTH*2-1+0:0] tmp00_56_79;
	wire [WIDTH*2-1+0:0] tmp00_56_80;
	wire [WIDTH*2-1+0:0] tmp00_56_81;
	wire [WIDTH*2-1+0:0] tmp00_56_82;
	wire [WIDTH*2-1+0:0] tmp00_56_83;
	wire [WIDTH*2-1+0:0] tmp00_57_0;
	wire [WIDTH*2-1+0:0] tmp00_57_1;
	wire [WIDTH*2-1+0:0] tmp00_57_2;
	wire [WIDTH*2-1+0:0] tmp00_57_3;
	wire [WIDTH*2-1+0:0] tmp00_57_4;
	wire [WIDTH*2-1+0:0] tmp00_57_5;
	wire [WIDTH*2-1+0:0] tmp00_57_6;
	wire [WIDTH*2-1+0:0] tmp00_57_7;
	wire [WIDTH*2-1+0:0] tmp00_57_8;
	wire [WIDTH*2-1+0:0] tmp00_57_9;
	wire [WIDTH*2-1+0:0] tmp00_57_10;
	wire [WIDTH*2-1+0:0] tmp00_57_11;
	wire [WIDTH*2-1+0:0] tmp00_57_12;
	wire [WIDTH*2-1+0:0] tmp00_57_13;
	wire [WIDTH*2-1+0:0] tmp00_57_14;
	wire [WIDTH*2-1+0:0] tmp00_57_15;
	wire [WIDTH*2-1+0:0] tmp00_57_16;
	wire [WIDTH*2-1+0:0] tmp00_57_17;
	wire [WIDTH*2-1+0:0] tmp00_57_18;
	wire [WIDTH*2-1+0:0] tmp00_57_19;
	wire [WIDTH*2-1+0:0] tmp00_57_20;
	wire [WIDTH*2-1+0:0] tmp00_57_21;
	wire [WIDTH*2-1+0:0] tmp00_57_22;
	wire [WIDTH*2-1+0:0] tmp00_57_23;
	wire [WIDTH*2-1+0:0] tmp00_57_24;
	wire [WIDTH*2-1+0:0] tmp00_57_25;
	wire [WIDTH*2-1+0:0] tmp00_57_26;
	wire [WIDTH*2-1+0:0] tmp00_57_27;
	wire [WIDTH*2-1+0:0] tmp00_57_28;
	wire [WIDTH*2-1+0:0] tmp00_57_29;
	wire [WIDTH*2-1+0:0] tmp00_57_30;
	wire [WIDTH*2-1+0:0] tmp00_57_31;
	wire [WIDTH*2-1+0:0] tmp00_57_32;
	wire [WIDTH*2-1+0:0] tmp00_57_33;
	wire [WIDTH*2-1+0:0] tmp00_57_34;
	wire [WIDTH*2-1+0:0] tmp00_57_35;
	wire [WIDTH*2-1+0:0] tmp00_57_36;
	wire [WIDTH*2-1+0:0] tmp00_57_37;
	wire [WIDTH*2-1+0:0] tmp00_57_38;
	wire [WIDTH*2-1+0:0] tmp00_57_39;
	wire [WIDTH*2-1+0:0] tmp00_57_40;
	wire [WIDTH*2-1+0:0] tmp00_57_41;
	wire [WIDTH*2-1+0:0] tmp00_57_42;
	wire [WIDTH*2-1+0:0] tmp00_57_43;
	wire [WIDTH*2-1+0:0] tmp00_57_44;
	wire [WIDTH*2-1+0:0] tmp00_57_45;
	wire [WIDTH*2-1+0:0] tmp00_57_46;
	wire [WIDTH*2-1+0:0] tmp00_57_47;
	wire [WIDTH*2-1+0:0] tmp00_57_48;
	wire [WIDTH*2-1+0:0] tmp00_57_49;
	wire [WIDTH*2-1+0:0] tmp00_57_50;
	wire [WIDTH*2-1+0:0] tmp00_57_51;
	wire [WIDTH*2-1+0:0] tmp00_57_52;
	wire [WIDTH*2-1+0:0] tmp00_57_53;
	wire [WIDTH*2-1+0:0] tmp00_57_54;
	wire [WIDTH*2-1+0:0] tmp00_57_55;
	wire [WIDTH*2-1+0:0] tmp00_57_56;
	wire [WIDTH*2-1+0:0] tmp00_57_57;
	wire [WIDTH*2-1+0:0] tmp00_57_58;
	wire [WIDTH*2-1+0:0] tmp00_57_59;
	wire [WIDTH*2-1+0:0] tmp00_57_60;
	wire [WIDTH*2-1+0:0] tmp00_57_61;
	wire [WIDTH*2-1+0:0] tmp00_57_62;
	wire [WIDTH*2-1+0:0] tmp00_57_63;
	wire [WIDTH*2-1+0:0] tmp00_57_64;
	wire [WIDTH*2-1+0:0] tmp00_57_65;
	wire [WIDTH*2-1+0:0] tmp00_57_66;
	wire [WIDTH*2-1+0:0] tmp00_57_67;
	wire [WIDTH*2-1+0:0] tmp00_57_68;
	wire [WIDTH*2-1+0:0] tmp00_57_69;
	wire [WIDTH*2-1+0:0] tmp00_57_70;
	wire [WIDTH*2-1+0:0] tmp00_57_71;
	wire [WIDTH*2-1+0:0] tmp00_57_72;
	wire [WIDTH*2-1+0:0] tmp00_57_73;
	wire [WIDTH*2-1+0:0] tmp00_57_74;
	wire [WIDTH*2-1+0:0] tmp00_57_75;
	wire [WIDTH*2-1+0:0] tmp00_57_76;
	wire [WIDTH*2-1+0:0] tmp00_57_77;
	wire [WIDTH*2-1+0:0] tmp00_57_78;
	wire [WIDTH*2-1+0:0] tmp00_57_79;
	wire [WIDTH*2-1+0:0] tmp00_57_80;
	wire [WIDTH*2-1+0:0] tmp00_57_81;
	wire [WIDTH*2-1+0:0] tmp00_57_82;
	wire [WIDTH*2-1+0:0] tmp00_57_83;
	wire [WIDTH*2-1+0:0] tmp00_58_0;
	wire [WIDTH*2-1+0:0] tmp00_58_1;
	wire [WIDTH*2-1+0:0] tmp00_58_2;
	wire [WIDTH*2-1+0:0] tmp00_58_3;
	wire [WIDTH*2-1+0:0] tmp00_58_4;
	wire [WIDTH*2-1+0:0] tmp00_58_5;
	wire [WIDTH*2-1+0:0] tmp00_58_6;
	wire [WIDTH*2-1+0:0] tmp00_58_7;
	wire [WIDTH*2-1+0:0] tmp00_58_8;
	wire [WIDTH*2-1+0:0] tmp00_58_9;
	wire [WIDTH*2-1+0:0] tmp00_58_10;
	wire [WIDTH*2-1+0:0] tmp00_58_11;
	wire [WIDTH*2-1+0:0] tmp00_58_12;
	wire [WIDTH*2-1+0:0] tmp00_58_13;
	wire [WIDTH*2-1+0:0] tmp00_58_14;
	wire [WIDTH*2-1+0:0] tmp00_58_15;
	wire [WIDTH*2-1+0:0] tmp00_58_16;
	wire [WIDTH*2-1+0:0] tmp00_58_17;
	wire [WIDTH*2-1+0:0] tmp00_58_18;
	wire [WIDTH*2-1+0:0] tmp00_58_19;
	wire [WIDTH*2-1+0:0] tmp00_58_20;
	wire [WIDTH*2-1+0:0] tmp00_58_21;
	wire [WIDTH*2-1+0:0] tmp00_58_22;
	wire [WIDTH*2-1+0:0] tmp00_58_23;
	wire [WIDTH*2-1+0:0] tmp00_58_24;
	wire [WIDTH*2-1+0:0] tmp00_58_25;
	wire [WIDTH*2-1+0:0] tmp00_58_26;
	wire [WIDTH*2-1+0:0] tmp00_58_27;
	wire [WIDTH*2-1+0:0] tmp00_58_28;
	wire [WIDTH*2-1+0:0] tmp00_58_29;
	wire [WIDTH*2-1+0:0] tmp00_58_30;
	wire [WIDTH*2-1+0:0] tmp00_58_31;
	wire [WIDTH*2-1+0:0] tmp00_58_32;
	wire [WIDTH*2-1+0:0] tmp00_58_33;
	wire [WIDTH*2-1+0:0] tmp00_58_34;
	wire [WIDTH*2-1+0:0] tmp00_58_35;
	wire [WIDTH*2-1+0:0] tmp00_58_36;
	wire [WIDTH*2-1+0:0] tmp00_58_37;
	wire [WIDTH*2-1+0:0] tmp00_58_38;
	wire [WIDTH*2-1+0:0] tmp00_58_39;
	wire [WIDTH*2-1+0:0] tmp00_58_40;
	wire [WIDTH*2-1+0:0] tmp00_58_41;
	wire [WIDTH*2-1+0:0] tmp00_58_42;
	wire [WIDTH*2-1+0:0] tmp00_58_43;
	wire [WIDTH*2-1+0:0] tmp00_58_44;
	wire [WIDTH*2-1+0:0] tmp00_58_45;
	wire [WIDTH*2-1+0:0] tmp00_58_46;
	wire [WIDTH*2-1+0:0] tmp00_58_47;
	wire [WIDTH*2-1+0:0] tmp00_58_48;
	wire [WIDTH*2-1+0:0] tmp00_58_49;
	wire [WIDTH*2-1+0:0] tmp00_58_50;
	wire [WIDTH*2-1+0:0] tmp00_58_51;
	wire [WIDTH*2-1+0:0] tmp00_58_52;
	wire [WIDTH*2-1+0:0] tmp00_58_53;
	wire [WIDTH*2-1+0:0] tmp00_58_54;
	wire [WIDTH*2-1+0:0] tmp00_58_55;
	wire [WIDTH*2-1+0:0] tmp00_58_56;
	wire [WIDTH*2-1+0:0] tmp00_58_57;
	wire [WIDTH*2-1+0:0] tmp00_58_58;
	wire [WIDTH*2-1+0:0] tmp00_58_59;
	wire [WIDTH*2-1+0:0] tmp00_58_60;
	wire [WIDTH*2-1+0:0] tmp00_58_61;
	wire [WIDTH*2-1+0:0] tmp00_58_62;
	wire [WIDTH*2-1+0:0] tmp00_58_63;
	wire [WIDTH*2-1+0:0] tmp00_58_64;
	wire [WIDTH*2-1+0:0] tmp00_58_65;
	wire [WIDTH*2-1+0:0] tmp00_58_66;
	wire [WIDTH*2-1+0:0] tmp00_58_67;
	wire [WIDTH*2-1+0:0] tmp00_58_68;
	wire [WIDTH*2-1+0:0] tmp00_58_69;
	wire [WIDTH*2-1+0:0] tmp00_58_70;
	wire [WIDTH*2-1+0:0] tmp00_58_71;
	wire [WIDTH*2-1+0:0] tmp00_58_72;
	wire [WIDTH*2-1+0:0] tmp00_58_73;
	wire [WIDTH*2-1+0:0] tmp00_58_74;
	wire [WIDTH*2-1+0:0] tmp00_58_75;
	wire [WIDTH*2-1+0:0] tmp00_58_76;
	wire [WIDTH*2-1+0:0] tmp00_58_77;
	wire [WIDTH*2-1+0:0] tmp00_58_78;
	wire [WIDTH*2-1+0:0] tmp00_58_79;
	wire [WIDTH*2-1+0:0] tmp00_58_80;
	wire [WIDTH*2-1+0:0] tmp00_58_81;
	wire [WIDTH*2-1+0:0] tmp00_58_82;
	wire [WIDTH*2-1+0:0] tmp00_58_83;
	wire [WIDTH*2-1+0:0] tmp00_59_0;
	wire [WIDTH*2-1+0:0] tmp00_59_1;
	wire [WIDTH*2-1+0:0] tmp00_59_2;
	wire [WIDTH*2-1+0:0] tmp00_59_3;
	wire [WIDTH*2-1+0:0] tmp00_59_4;
	wire [WIDTH*2-1+0:0] tmp00_59_5;
	wire [WIDTH*2-1+0:0] tmp00_59_6;
	wire [WIDTH*2-1+0:0] tmp00_59_7;
	wire [WIDTH*2-1+0:0] tmp00_59_8;
	wire [WIDTH*2-1+0:0] tmp00_59_9;
	wire [WIDTH*2-1+0:0] tmp00_59_10;
	wire [WIDTH*2-1+0:0] tmp00_59_11;
	wire [WIDTH*2-1+0:0] tmp00_59_12;
	wire [WIDTH*2-1+0:0] tmp00_59_13;
	wire [WIDTH*2-1+0:0] tmp00_59_14;
	wire [WIDTH*2-1+0:0] tmp00_59_15;
	wire [WIDTH*2-1+0:0] tmp00_59_16;
	wire [WIDTH*2-1+0:0] tmp00_59_17;
	wire [WIDTH*2-1+0:0] tmp00_59_18;
	wire [WIDTH*2-1+0:0] tmp00_59_19;
	wire [WIDTH*2-1+0:0] tmp00_59_20;
	wire [WIDTH*2-1+0:0] tmp00_59_21;
	wire [WIDTH*2-1+0:0] tmp00_59_22;
	wire [WIDTH*2-1+0:0] tmp00_59_23;
	wire [WIDTH*2-1+0:0] tmp00_59_24;
	wire [WIDTH*2-1+0:0] tmp00_59_25;
	wire [WIDTH*2-1+0:0] tmp00_59_26;
	wire [WIDTH*2-1+0:0] tmp00_59_27;
	wire [WIDTH*2-1+0:0] tmp00_59_28;
	wire [WIDTH*2-1+0:0] tmp00_59_29;
	wire [WIDTH*2-1+0:0] tmp00_59_30;
	wire [WIDTH*2-1+0:0] tmp00_59_31;
	wire [WIDTH*2-1+0:0] tmp00_59_32;
	wire [WIDTH*2-1+0:0] tmp00_59_33;
	wire [WIDTH*2-1+0:0] tmp00_59_34;
	wire [WIDTH*2-1+0:0] tmp00_59_35;
	wire [WIDTH*2-1+0:0] tmp00_59_36;
	wire [WIDTH*2-1+0:0] tmp00_59_37;
	wire [WIDTH*2-1+0:0] tmp00_59_38;
	wire [WIDTH*2-1+0:0] tmp00_59_39;
	wire [WIDTH*2-1+0:0] tmp00_59_40;
	wire [WIDTH*2-1+0:0] tmp00_59_41;
	wire [WIDTH*2-1+0:0] tmp00_59_42;
	wire [WIDTH*2-1+0:0] tmp00_59_43;
	wire [WIDTH*2-1+0:0] tmp00_59_44;
	wire [WIDTH*2-1+0:0] tmp00_59_45;
	wire [WIDTH*2-1+0:0] tmp00_59_46;
	wire [WIDTH*2-1+0:0] tmp00_59_47;
	wire [WIDTH*2-1+0:0] tmp00_59_48;
	wire [WIDTH*2-1+0:0] tmp00_59_49;
	wire [WIDTH*2-1+0:0] tmp00_59_50;
	wire [WIDTH*2-1+0:0] tmp00_59_51;
	wire [WIDTH*2-1+0:0] tmp00_59_52;
	wire [WIDTH*2-1+0:0] tmp00_59_53;
	wire [WIDTH*2-1+0:0] tmp00_59_54;
	wire [WIDTH*2-1+0:0] tmp00_59_55;
	wire [WIDTH*2-1+0:0] tmp00_59_56;
	wire [WIDTH*2-1+0:0] tmp00_59_57;
	wire [WIDTH*2-1+0:0] tmp00_59_58;
	wire [WIDTH*2-1+0:0] tmp00_59_59;
	wire [WIDTH*2-1+0:0] tmp00_59_60;
	wire [WIDTH*2-1+0:0] tmp00_59_61;
	wire [WIDTH*2-1+0:0] tmp00_59_62;
	wire [WIDTH*2-1+0:0] tmp00_59_63;
	wire [WIDTH*2-1+0:0] tmp00_59_64;
	wire [WIDTH*2-1+0:0] tmp00_59_65;
	wire [WIDTH*2-1+0:0] tmp00_59_66;
	wire [WIDTH*2-1+0:0] tmp00_59_67;
	wire [WIDTH*2-1+0:0] tmp00_59_68;
	wire [WIDTH*2-1+0:0] tmp00_59_69;
	wire [WIDTH*2-1+0:0] tmp00_59_70;
	wire [WIDTH*2-1+0:0] tmp00_59_71;
	wire [WIDTH*2-1+0:0] tmp00_59_72;
	wire [WIDTH*2-1+0:0] tmp00_59_73;
	wire [WIDTH*2-1+0:0] tmp00_59_74;
	wire [WIDTH*2-1+0:0] tmp00_59_75;
	wire [WIDTH*2-1+0:0] tmp00_59_76;
	wire [WIDTH*2-1+0:0] tmp00_59_77;
	wire [WIDTH*2-1+0:0] tmp00_59_78;
	wire [WIDTH*2-1+0:0] tmp00_59_79;
	wire [WIDTH*2-1+0:0] tmp00_59_80;
	wire [WIDTH*2-1+0:0] tmp00_59_81;
	wire [WIDTH*2-1+0:0] tmp00_59_82;
	wire [WIDTH*2-1+0:0] tmp00_59_83;
	wire [WIDTH*2-1+0:0] tmp00_60_0;
	wire [WIDTH*2-1+0:0] tmp00_60_1;
	wire [WIDTH*2-1+0:0] tmp00_60_2;
	wire [WIDTH*2-1+0:0] tmp00_60_3;
	wire [WIDTH*2-1+0:0] tmp00_60_4;
	wire [WIDTH*2-1+0:0] tmp00_60_5;
	wire [WIDTH*2-1+0:0] tmp00_60_6;
	wire [WIDTH*2-1+0:0] tmp00_60_7;
	wire [WIDTH*2-1+0:0] tmp00_60_8;
	wire [WIDTH*2-1+0:0] tmp00_60_9;
	wire [WIDTH*2-1+0:0] tmp00_60_10;
	wire [WIDTH*2-1+0:0] tmp00_60_11;
	wire [WIDTH*2-1+0:0] tmp00_60_12;
	wire [WIDTH*2-1+0:0] tmp00_60_13;
	wire [WIDTH*2-1+0:0] tmp00_60_14;
	wire [WIDTH*2-1+0:0] tmp00_60_15;
	wire [WIDTH*2-1+0:0] tmp00_60_16;
	wire [WIDTH*2-1+0:0] tmp00_60_17;
	wire [WIDTH*2-1+0:0] tmp00_60_18;
	wire [WIDTH*2-1+0:0] tmp00_60_19;
	wire [WIDTH*2-1+0:0] tmp00_60_20;
	wire [WIDTH*2-1+0:0] tmp00_60_21;
	wire [WIDTH*2-1+0:0] tmp00_60_22;
	wire [WIDTH*2-1+0:0] tmp00_60_23;
	wire [WIDTH*2-1+0:0] tmp00_60_24;
	wire [WIDTH*2-1+0:0] tmp00_60_25;
	wire [WIDTH*2-1+0:0] tmp00_60_26;
	wire [WIDTH*2-1+0:0] tmp00_60_27;
	wire [WIDTH*2-1+0:0] tmp00_60_28;
	wire [WIDTH*2-1+0:0] tmp00_60_29;
	wire [WIDTH*2-1+0:0] tmp00_60_30;
	wire [WIDTH*2-1+0:0] tmp00_60_31;
	wire [WIDTH*2-1+0:0] tmp00_60_32;
	wire [WIDTH*2-1+0:0] tmp00_60_33;
	wire [WIDTH*2-1+0:0] tmp00_60_34;
	wire [WIDTH*2-1+0:0] tmp00_60_35;
	wire [WIDTH*2-1+0:0] tmp00_60_36;
	wire [WIDTH*2-1+0:0] tmp00_60_37;
	wire [WIDTH*2-1+0:0] tmp00_60_38;
	wire [WIDTH*2-1+0:0] tmp00_60_39;
	wire [WIDTH*2-1+0:0] tmp00_60_40;
	wire [WIDTH*2-1+0:0] tmp00_60_41;
	wire [WIDTH*2-1+0:0] tmp00_60_42;
	wire [WIDTH*2-1+0:0] tmp00_60_43;
	wire [WIDTH*2-1+0:0] tmp00_60_44;
	wire [WIDTH*2-1+0:0] tmp00_60_45;
	wire [WIDTH*2-1+0:0] tmp00_60_46;
	wire [WIDTH*2-1+0:0] tmp00_60_47;
	wire [WIDTH*2-1+0:0] tmp00_60_48;
	wire [WIDTH*2-1+0:0] tmp00_60_49;
	wire [WIDTH*2-1+0:0] tmp00_60_50;
	wire [WIDTH*2-1+0:0] tmp00_60_51;
	wire [WIDTH*2-1+0:0] tmp00_60_52;
	wire [WIDTH*2-1+0:0] tmp00_60_53;
	wire [WIDTH*2-1+0:0] tmp00_60_54;
	wire [WIDTH*2-1+0:0] tmp00_60_55;
	wire [WIDTH*2-1+0:0] tmp00_60_56;
	wire [WIDTH*2-1+0:0] tmp00_60_57;
	wire [WIDTH*2-1+0:0] tmp00_60_58;
	wire [WIDTH*2-1+0:0] tmp00_60_59;
	wire [WIDTH*2-1+0:0] tmp00_60_60;
	wire [WIDTH*2-1+0:0] tmp00_60_61;
	wire [WIDTH*2-1+0:0] tmp00_60_62;
	wire [WIDTH*2-1+0:0] tmp00_60_63;
	wire [WIDTH*2-1+0:0] tmp00_60_64;
	wire [WIDTH*2-1+0:0] tmp00_60_65;
	wire [WIDTH*2-1+0:0] tmp00_60_66;
	wire [WIDTH*2-1+0:0] tmp00_60_67;
	wire [WIDTH*2-1+0:0] tmp00_60_68;
	wire [WIDTH*2-1+0:0] tmp00_60_69;
	wire [WIDTH*2-1+0:0] tmp00_60_70;
	wire [WIDTH*2-1+0:0] tmp00_60_71;
	wire [WIDTH*2-1+0:0] tmp00_60_72;
	wire [WIDTH*2-1+0:0] tmp00_60_73;
	wire [WIDTH*2-1+0:0] tmp00_60_74;
	wire [WIDTH*2-1+0:0] tmp00_60_75;
	wire [WIDTH*2-1+0:0] tmp00_60_76;
	wire [WIDTH*2-1+0:0] tmp00_60_77;
	wire [WIDTH*2-1+0:0] tmp00_60_78;
	wire [WIDTH*2-1+0:0] tmp00_60_79;
	wire [WIDTH*2-1+0:0] tmp00_60_80;
	wire [WIDTH*2-1+0:0] tmp00_60_81;
	wire [WIDTH*2-1+0:0] tmp00_60_82;
	wire [WIDTH*2-1+0:0] tmp00_60_83;
	wire [WIDTH*2-1+0:0] tmp00_61_0;
	wire [WIDTH*2-1+0:0] tmp00_61_1;
	wire [WIDTH*2-1+0:0] tmp00_61_2;
	wire [WIDTH*2-1+0:0] tmp00_61_3;
	wire [WIDTH*2-1+0:0] tmp00_61_4;
	wire [WIDTH*2-1+0:0] tmp00_61_5;
	wire [WIDTH*2-1+0:0] tmp00_61_6;
	wire [WIDTH*2-1+0:0] tmp00_61_7;
	wire [WIDTH*2-1+0:0] tmp00_61_8;
	wire [WIDTH*2-1+0:0] tmp00_61_9;
	wire [WIDTH*2-1+0:0] tmp00_61_10;
	wire [WIDTH*2-1+0:0] tmp00_61_11;
	wire [WIDTH*2-1+0:0] tmp00_61_12;
	wire [WIDTH*2-1+0:0] tmp00_61_13;
	wire [WIDTH*2-1+0:0] tmp00_61_14;
	wire [WIDTH*2-1+0:0] tmp00_61_15;
	wire [WIDTH*2-1+0:0] tmp00_61_16;
	wire [WIDTH*2-1+0:0] tmp00_61_17;
	wire [WIDTH*2-1+0:0] tmp00_61_18;
	wire [WIDTH*2-1+0:0] tmp00_61_19;
	wire [WIDTH*2-1+0:0] tmp00_61_20;
	wire [WIDTH*2-1+0:0] tmp00_61_21;
	wire [WIDTH*2-1+0:0] tmp00_61_22;
	wire [WIDTH*2-1+0:0] tmp00_61_23;
	wire [WIDTH*2-1+0:0] tmp00_61_24;
	wire [WIDTH*2-1+0:0] tmp00_61_25;
	wire [WIDTH*2-1+0:0] tmp00_61_26;
	wire [WIDTH*2-1+0:0] tmp00_61_27;
	wire [WIDTH*2-1+0:0] tmp00_61_28;
	wire [WIDTH*2-1+0:0] tmp00_61_29;
	wire [WIDTH*2-1+0:0] tmp00_61_30;
	wire [WIDTH*2-1+0:0] tmp00_61_31;
	wire [WIDTH*2-1+0:0] tmp00_61_32;
	wire [WIDTH*2-1+0:0] tmp00_61_33;
	wire [WIDTH*2-1+0:0] tmp00_61_34;
	wire [WIDTH*2-1+0:0] tmp00_61_35;
	wire [WIDTH*2-1+0:0] tmp00_61_36;
	wire [WIDTH*2-1+0:0] tmp00_61_37;
	wire [WIDTH*2-1+0:0] tmp00_61_38;
	wire [WIDTH*2-1+0:0] tmp00_61_39;
	wire [WIDTH*2-1+0:0] tmp00_61_40;
	wire [WIDTH*2-1+0:0] tmp00_61_41;
	wire [WIDTH*2-1+0:0] tmp00_61_42;
	wire [WIDTH*2-1+0:0] tmp00_61_43;
	wire [WIDTH*2-1+0:0] tmp00_61_44;
	wire [WIDTH*2-1+0:0] tmp00_61_45;
	wire [WIDTH*2-1+0:0] tmp00_61_46;
	wire [WIDTH*2-1+0:0] tmp00_61_47;
	wire [WIDTH*2-1+0:0] tmp00_61_48;
	wire [WIDTH*2-1+0:0] tmp00_61_49;
	wire [WIDTH*2-1+0:0] tmp00_61_50;
	wire [WIDTH*2-1+0:0] tmp00_61_51;
	wire [WIDTH*2-1+0:0] tmp00_61_52;
	wire [WIDTH*2-1+0:0] tmp00_61_53;
	wire [WIDTH*2-1+0:0] tmp00_61_54;
	wire [WIDTH*2-1+0:0] tmp00_61_55;
	wire [WIDTH*2-1+0:0] tmp00_61_56;
	wire [WIDTH*2-1+0:0] tmp00_61_57;
	wire [WIDTH*2-1+0:0] tmp00_61_58;
	wire [WIDTH*2-1+0:0] tmp00_61_59;
	wire [WIDTH*2-1+0:0] tmp00_61_60;
	wire [WIDTH*2-1+0:0] tmp00_61_61;
	wire [WIDTH*2-1+0:0] tmp00_61_62;
	wire [WIDTH*2-1+0:0] tmp00_61_63;
	wire [WIDTH*2-1+0:0] tmp00_61_64;
	wire [WIDTH*2-1+0:0] tmp00_61_65;
	wire [WIDTH*2-1+0:0] tmp00_61_66;
	wire [WIDTH*2-1+0:0] tmp00_61_67;
	wire [WIDTH*2-1+0:0] tmp00_61_68;
	wire [WIDTH*2-1+0:0] tmp00_61_69;
	wire [WIDTH*2-1+0:0] tmp00_61_70;
	wire [WIDTH*2-1+0:0] tmp00_61_71;
	wire [WIDTH*2-1+0:0] tmp00_61_72;
	wire [WIDTH*2-1+0:0] tmp00_61_73;
	wire [WIDTH*2-1+0:0] tmp00_61_74;
	wire [WIDTH*2-1+0:0] tmp00_61_75;
	wire [WIDTH*2-1+0:0] tmp00_61_76;
	wire [WIDTH*2-1+0:0] tmp00_61_77;
	wire [WIDTH*2-1+0:0] tmp00_61_78;
	wire [WIDTH*2-1+0:0] tmp00_61_79;
	wire [WIDTH*2-1+0:0] tmp00_61_80;
	wire [WIDTH*2-1+0:0] tmp00_61_81;
	wire [WIDTH*2-1+0:0] tmp00_61_82;
	wire [WIDTH*2-1+0:0] tmp00_61_83;
	wire [WIDTH*2-1+0:0] tmp00_62_0;
	wire [WIDTH*2-1+0:0] tmp00_62_1;
	wire [WIDTH*2-1+0:0] tmp00_62_2;
	wire [WIDTH*2-1+0:0] tmp00_62_3;
	wire [WIDTH*2-1+0:0] tmp00_62_4;
	wire [WIDTH*2-1+0:0] tmp00_62_5;
	wire [WIDTH*2-1+0:0] tmp00_62_6;
	wire [WIDTH*2-1+0:0] tmp00_62_7;
	wire [WIDTH*2-1+0:0] tmp00_62_8;
	wire [WIDTH*2-1+0:0] tmp00_62_9;
	wire [WIDTH*2-1+0:0] tmp00_62_10;
	wire [WIDTH*2-1+0:0] tmp00_62_11;
	wire [WIDTH*2-1+0:0] tmp00_62_12;
	wire [WIDTH*2-1+0:0] tmp00_62_13;
	wire [WIDTH*2-1+0:0] tmp00_62_14;
	wire [WIDTH*2-1+0:0] tmp00_62_15;
	wire [WIDTH*2-1+0:0] tmp00_62_16;
	wire [WIDTH*2-1+0:0] tmp00_62_17;
	wire [WIDTH*2-1+0:0] tmp00_62_18;
	wire [WIDTH*2-1+0:0] tmp00_62_19;
	wire [WIDTH*2-1+0:0] tmp00_62_20;
	wire [WIDTH*2-1+0:0] tmp00_62_21;
	wire [WIDTH*2-1+0:0] tmp00_62_22;
	wire [WIDTH*2-1+0:0] tmp00_62_23;
	wire [WIDTH*2-1+0:0] tmp00_62_24;
	wire [WIDTH*2-1+0:0] tmp00_62_25;
	wire [WIDTH*2-1+0:0] tmp00_62_26;
	wire [WIDTH*2-1+0:0] tmp00_62_27;
	wire [WIDTH*2-1+0:0] tmp00_62_28;
	wire [WIDTH*2-1+0:0] tmp00_62_29;
	wire [WIDTH*2-1+0:0] tmp00_62_30;
	wire [WIDTH*2-1+0:0] tmp00_62_31;
	wire [WIDTH*2-1+0:0] tmp00_62_32;
	wire [WIDTH*2-1+0:0] tmp00_62_33;
	wire [WIDTH*2-1+0:0] tmp00_62_34;
	wire [WIDTH*2-1+0:0] tmp00_62_35;
	wire [WIDTH*2-1+0:0] tmp00_62_36;
	wire [WIDTH*2-1+0:0] tmp00_62_37;
	wire [WIDTH*2-1+0:0] tmp00_62_38;
	wire [WIDTH*2-1+0:0] tmp00_62_39;
	wire [WIDTH*2-1+0:0] tmp00_62_40;
	wire [WIDTH*2-1+0:0] tmp00_62_41;
	wire [WIDTH*2-1+0:0] tmp00_62_42;
	wire [WIDTH*2-1+0:0] tmp00_62_43;
	wire [WIDTH*2-1+0:0] tmp00_62_44;
	wire [WIDTH*2-1+0:0] tmp00_62_45;
	wire [WIDTH*2-1+0:0] tmp00_62_46;
	wire [WIDTH*2-1+0:0] tmp00_62_47;
	wire [WIDTH*2-1+0:0] tmp00_62_48;
	wire [WIDTH*2-1+0:0] tmp00_62_49;
	wire [WIDTH*2-1+0:0] tmp00_62_50;
	wire [WIDTH*2-1+0:0] tmp00_62_51;
	wire [WIDTH*2-1+0:0] tmp00_62_52;
	wire [WIDTH*2-1+0:0] tmp00_62_53;
	wire [WIDTH*2-1+0:0] tmp00_62_54;
	wire [WIDTH*2-1+0:0] tmp00_62_55;
	wire [WIDTH*2-1+0:0] tmp00_62_56;
	wire [WIDTH*2-1+0:0] tmp00_62_57;
	wire [WIDTH*2-1+0:0] tmp00_62_58;
	wire [WIDTH*2-1+0:0] tmp00_62_59;
	wire [WIDTH*2-1+0:0] tmp00_62_60;
	wire [WIDTH*2-1+0:0] tmp00_62_61;
	wire [WIDTH*2-1+0:0] tmp00_62_62;
	wire [WIDTH*2-1+0:0] tmp00_62_63;
	wire [WIDTH*2-1+0:0] tmp00_62_64;
	wire [WIDTH*2-1+0:0] tmp00_62_65;
	wire [WIDTH*2-1+0:0] tmp00_62_66;
	wire [WIDTH*2-1+0:0] tmp00_62_67;
	wire [WIDTH*2-1+0:0] tmp00_62_68;
	wire [WIDTH*2-1+0:0] tmp00_62_69;
	wire [WIDTH*2-1+0:0] tmp00_62_70;
	wire [WIDTH*2-1+0:0] tmp00_62_71;
	wire [WIDTH*2-1+0:0] tmp00_62_72;
	wire [WIDTH*2-1+0:0] tmp00_62_73;
	wire [WIDTH*2-1+0:0] tmp00_62_74;
	wire [WIDTH*2-1+0:0] tmp00_62_75;
	wire [WIDTH*2-1+0:0] tmp00_62_76;
	wire [WIDTH*2-1+0:0] tmp00_62_77;
	wire [WIDTH*2-1+0:0] tmp00_62_78;
	wire [WIDTH*2-1+0:0] tmp00_62_79;
	wire [WIDTH*2-1+0:0] tmp00_62_80;
	wire [WIDTH*2-1+0:0] tmp00_62_81;
	wire [WIDTH*2-1+0:0] tmp00_62_82;
	wire [WIDTH*2-1+0:0] tmp00_62_83;
	wire [WIDTH*2-1+0:0] tmp00_63_0;
	wire [WIDTH*2-1+0:0] tmp00_63_1;
	wire [WIDTH*2-1+0:0] tmp00_63_2;
	wire [WIDTH*2-1+0:0] tmp00_63_3;
	wire [WIDTH*2-1+0:0] tmp00_63_4;
	wire [WIDTH*2-1+0:0] tmp00_63_5;
	wire [WIDTH*2-1+0:0] tmp00_63_6;
	wire [WIDTH*2-1+0:0] tmp00_63_7;
	wire [WIDTH*2-1+0:0] tmp00_63_8;
	wire [WIDTH*2-1+0:0] tmp00_63_9;
	wire [WIDTH*2-1+0:0] tmp00_63_10;
	wire [WIDTH*2-1+0:0] tmp00_63_11;
	wire [WIDTH*2-1+0:0] tmp00_63_12;
	wire [WIDTH*2-1+0:0] tmp00_63_13;
	wire [WIDTH*2-1+0:0] tmp00_63_14;
	wire [WIDTH*2-1+0:0] tmp00_63_15;
	wire [WIDTH*2-1+0:0] tmp00_63_16;
	wire [WIDTH*2-1+0:0] tmp00_63_17;
	wire [WIDTH*2-1+0:0] tmp00_63_18;
	wire [WIDTH*2-1+0:0] tmp00_63_19;
	wire [WIDTH*2-1+0:0] tmp00_63_20;
	wire [WIDTH*2-1+0:0] tmp00_63_21;
	wire [WIDTH*2-1+0:0] tmp00_63_22;
	wire [WIDTH*2-1+0:0] tmp00_63_23;
	wire [WIDTH*2-1+0:0] tmp00_63_24;
	wire [WIDTH*2-1+0:0] tmp00_63_25;
	wire [WIDTH*2-1+0:0] tmp00_63_26;
	wire [WIDTH*2-1+0:0] tmp00_63_27;
	wire [WIDTH*2-1+0:0] tmp00_63_28;
	wire [WIDTH*2-1+0:0] tmp00_63_29;
	wire [WIDTH*2-1+0:0] tmp00_63_30;
	wire [WIDTH*2-1+0:0] tmp00_63_31;
	wire [WIDTH*2-1+0:0] tmp00_63_32;
	wire [WIDTH*2-1+0:0] tmp00_63_33;
	wire [WIDTH*2-1+0:0] tmp00_63_34;
	wire [WIDTH*2-1+0:0] tmp00_63_35;
	wire [WIDTH*2-1+0:0] tmp00_63_36;
	wire [WIDTH*2-1+0:0] tmp00_63_37;
	wire [WIDTH*2-1+0:0] tmp00_63_38;
	wire [WIDTH*2-1+0:0] tmp00_63_39;
	wire [WIDTH*2-1+0:0] tmp00_63_40;
	wire [WIDTH*2-1+0:0] tmp00_63_41;
	wire [WIDTH*2-1+0:0] tmp00_63_42;
	wire [WIDTH*2-1+0:0] tmp00_63_43;
	wire [WIDTH*2-1+0:0] tmp00_63_44;
	wire [WIDTH*2-1+0:0] tmp00_63_45;
	wire [WIDTH*2-1+0:0] tmp00_63_46;
	wire [WIDTH*2-1+0:0] tmp00_63_47;
	wire [WIDTH*2-1+0:0] tmp00_63_48;
	wire [WIDTH*2-1+0:0] tmp00_63_49;
	wire [WIDTH*2-1+0:0] tmp00_63_50;
	wire [WIDTH*2-1+0:0] tmp00_63_51;
	wire [WIDTH*2-1+0:0] tmp00_63_52;
	wire [WIDTH*2-1+0:0] tmp00_63_53;
	wire [WIDTH*2-1+0:0] tmp00_63_54;
	wire [WIDTH*2-1+0:0] tmp00_63_55;
	wire [WIDTH*2-1+0:0] tmp00_63_56;
	wire [WIDTH*2-1+0:0] tmp00_63_57;
	wire [WIDTH*2-1+0:0] tmp00_63_58;
	wire [WIDTH*2-1+0:0] tmp00_63_59;
	wire [WIDTH*2-1+0:0] tmp00_63_60;
	wire [WIDTH*2-1+0:0] tmp00_63_61;
	wire [WIDTH*2-1+0:0] tmp00_63_62;
	wire [WIDTH*2-1+0:0] tmp00_63_63;
	wire [WIDTH*2-1+0:0] tmp00_63_64;
	wire [WIDTH*2-1+0:0] tmp00_63_65;
	wire [WIDTH*2-1+0:0] tmp00_63_66;
	wire [WIDTH*2-1+0:0] tmp00_63_67;
	wire [WIDTH*2-1+0:0] tmp00_63_68;
	wire [WIDTH*2-1+0:0] tmp00_63_69;
	wire [WIDTH*2-1+0:0] tmp00_63_70;
	wire [WIDTH*2-1+0:0] tmp00_63_71;
	wire [WIDTH*2-1+0:0] tmp00_63_72;
	wire [WIDTH*2-1+0:0] tmp00_63_73;
	wire [WIDTH*2-1+0:0] tmp00_63_74;
	wire [WIDTH*2-1+0:0] tmp00_63_75;
	wire [WIDTH*2-1+0:0] tmp00_63_76;
	wire [WIDTH*2-1+0:0] tmp00_63_77;
	wire [WIDTH*2-1+0:0] tmp00_63_78;
	wire [WIDTH*2-1+0:0] tmp00_63_79;
	wire [WIDTH*2-1+0:0] tmp00_63_80;
	wire [WIDTH*2-1+0:0] tmp00_63_81;
	wire [WIDTH*2-1+0:0] tmp00_63_82;
	wire [WIDTH*2-1+0:0] tmp00_63_83;
	wire [WIDTH*2-1+0:0] tmp00_64_0;
	wire [WIDTH*2-1+0:0] tmp00_64_1;
	wire [WIDTH*2-1+0:0] tmp00_64_2;
	wire [WIDTH*2-1+0:0] tmp00_64_3;
	wire [WIDTH*2-1+0:0] tmp00_64_4;
	wire [WIDTH*2-1+0:0] tmp00_64_5;
	wire [WIDTH*2-1+0:0] tmp00_64_6;
	wire [WIDTH*2-1+0:0] tmp00_64_7;
	wire [WIDTH*2-1+0:0] tmp00_64_8;
	wire [WIDTH*2-1+0:0] tmp00_64_9;
	wire [WIDTH*2-1+0:0] tmp00_64_10;
	wire [WIDTH*2-1+0:0] tmp00_64_11;
	wire [WIDTH*2-1+0:0] tmp00_64_12;
	wire [WIDTH*2-1+0:0] tmp00_64_13;
	wire [WIDTH*2-1+0:0] tmp00_64_14;
	wire [WIDTH*2-1+0:0] tmp00_64_15;
	wire [WIDTH*2-1+0:0] tmp00_64_16;
	wire [WIDTH*2-1+0:0] tmp00_64_17;
	wire [WIDTH*2-1+0:0] tmp00_64_18;
	wire [WIDTH*2-1+0:0] tmp00_64_19;
	wire [WIDTH*2-1+0:0] tmp00_64_20;
	wire [WIDTH*2-1+0:0] tmp00_64_21;
	wire [WIDTH*2-1+0:0] tmp00_64_22;
	wire [WIDTH*2-1+0:0] tmp00_64_23;
	wire [WIDTH*2-1+0:0] tmp00_64_24;
	wire [WIDTH*2-1+0:0] tmp00_64_25;
	wire [WIDTH*2-1+0:0] tmp00_64_26;
	wire [WIDTH*2-1+0:0] tmp00_64_27;
	wire [WIDTH*2-1+0:0] tmp00_64_28;
	wire [WIDTH*2-1+0:0] tmp00_64_29;
	wire [WIDTH*2-1+0:0] tmp00_64_30;
	wire [WIDTH*2-1+0:0] tmp00_64_31;
	wire [WIDTH*2-1+0:0] tmp00_64_32;
	wire [WIDTH*2-1+0:0] tmp00_64_33;
	wire [WIDTH*2-1+0:0] tmp00_64_34;
	wire [WIDTH*2-1+0:0] tmp00_64_35;
	wire [WIDTH*2-1+0:0] tmp00_64_36;
	wire [WIDTH*2-1+0:0] tmp00_64_37;
	wire [WIDTH*2-1+0:0] tmp00_64_38;
	wire [WIDTH*2-1+0:0] tmp00_64_39;
	wire [WIDTH*2-1+0:0] tmp00_64_40;
	wire [WIDTH*2-1+0:0] tmp00_64_41;
	wire [WIDTH*2-1+0:0] tmp00_64_42;
	wire [WIDTH*2-1+0:0] tmp00_64_43;
	wire [WIDTH*2-1+0:0] tmp00_64_44;
	wire [WIDTH*2-1+0:0] tmp00_64_45;
	wire [WIDTH*2-1+0:0] tmp00_64_46;
	wire [WIDTH*2-1+0:0] tmp00_64_47;
	wire [WIDTH*2-1+0:0] tmp00_64_48;
	wire [WIDTH*2-1+0:0] tmp00_64_49;
	wire [WIDTH*2-1+0:0] tmp00_64_50;
	wire [WIDTH*2-1+0:0] tmp00_64_51;
	wire [WIDTH*2-1+0:0] tmp00_64_52;
	wire [WIDTH*2-1+0:0] tmp00_64_53;
	wire [WIDTH*2-1+0:0] tmp00_64_54;
	wire [WIDTH*2-1+0:0] tmp00_64_55;
	wire [WIDTH*2-1+0:0] tmp00_64_56;
	wire [WIDTH*2-1+0:0] tmp00_64_57;
	wire [WIDTH*2-1+0:0] tmp00_64_58;
	wire [WIDTH*2-1+0:0] tmp00_64_59;
	wire [WIDTH*2-1+0:0] tmp00_64_60;
	wire [WIDTH*2-1+0:0] tmp00_64_61;
	wire [WIDTH*2-1+0:0] tmp00_64_62;
	wire [WIDTH*2-1+0:0] tmp00_64_63;
	wire [WIDTH*2-1+0:0] tmp00_64_64;
	wire [WIDTH*2-1+0:0] tmp00_64_65;
	wire [WIDTH*2-1+0:0] tmp00_64_66;
	wire [WIDTH*2-1+0:0] tmp00_64_67;
	wire [WIDTH*2-1+0:0] tmp00_64_68;
	wire [WIDTH*2-1+0:0] tmp00_64_69;
	wire [WIDTH*2-1+0:0] tmp00_64_70;
	wire [WIDTH*2-1+0:0] tmp00_64_71;
	wire [WIDTH*2-1+0:0] tmp00_64_72;
	wire [WIDTH*2-1+0:0] tmp00_64_73;
	wire [WIDTH*2-1+0:0] tmp00_64_74;
	wire [WIDTH*2-1+0:0] tmp00_64_75;
	wire [WIDTH*2-1+0:0] tmp00_64_76;
	wire [WIDTH*2-1+0:0] tmp00_64_77;
	wire [WIDTH*2-1+0:0] tmp00_64_78;
	wire [WIDTH*2-1+0:0] tmp00_64_79;
	wire [WIDTH*2-1+0:0] tmp00_64_80;
	wire [WIDTH*2-1+0:0] tmp00_64_81;
	wire [WIDTH*2-1+0:0] tmp00_64_82;
	wire [WIDTH*2-1+0:0] tmp00_64_83;
	wire [WIDTH*2-1+0:0] tmp00_65_0;
	wire [WIDTH*2-1+0:0] tmp00_65_1;
	wire [WIDTH*2-1+0:0] tmp00_65_2;
	wire [WIDTH*2-1+0:0] tmp00_65_3;
	wire [WIDTH*2-1+0:0] tmp00_65_4;
	wire [WIDTH*2-1+0:0] tmp00_65_5;
	wire [WIDTH*2-1+0:0] tmp00_65_6;
	wire [WIDTH*2-1+0:0] tmp00_65_7;
	wire [WIDTH*2-1+0:0] tmp00_65_8;
	wire [WIDTH*2-1+0:0] tmp00_65_9;
	wire [WIDTH*2-1+0:0] tmp00_65_10;
	wire [WIDTH*2-1+0:0] tmp00_65_11;
	wire [WIDTH*2-1+0:0] tmp00_65_12;
	wire [WIDTH*2-1+0:0] tmp00_65_13;
	wire [WIDTH*2-1+0:0] tmp00_65_14;
	wire [WIDTH*2-1+0:0] tmp00_65_15;
	wire [WIDTH*2-1+0:0] tmp00_65_16;
	wire [WIDTH*2-1+0:0] tmp00_65_17;
	wire [WIDTH*2-1+0:0] tmp00_65_18;
	wire [WIDTH*2-1+0:0] tmp00_65_19;
	wire [WIDTH*2-1+0:0] tmp00_65_20;
	wire [WIDTH*2-1+0:0] tmp00_65_21;
	wire [WIDTH*2-1+0:0] tmp00_65_22;
	wire [WIDTH*2-1+0:0] tmp00_65_23;
	wire [WIDTH*2-1+0:0] tmp00_65_24;
	wire [WIDTH*2-1+0:0] tmp00_65_25;
	wire [WIDTH*2-1+0:0] tmp00_65_26;
	wire [WIDTH*2-1+0:0] tmp00_65_27;
	wire [WIDTH*2-1+0:0] tmp00_65_28;
	wire [WIDTH*2-1+0:0] tmp00_65_29;
	wire [WIDTH*2-1+0:0] tmp00_65_30;
	wire [WIDTH*2-1+0:0] tmp00_65_31;
	wire [WIDTH*2-1+0:0] tmp00_65_32;
	wire [WIDTH*2-1+0:0] tmp00_65_33;
	wire [WIDTH*2-1+0:0] tmp00_65_34;
	wire [WIDTH*2-1+0:0] tmp00_65_35;
	wire [WIDTH*2-1+0:0] tmp00_65_36;
	wire [WIDTH*2-1+0:0] tmp00_65_37;
	wire [WIDTH*2-1+0:0] tmp00_65_38;
	wire [WIDTH*2-1+0:0] tmp00_65_39;
	wire [WIDTH*2-1+0:0] tmp00_65_40;
	wire [WIDTH*2-1+0:0] tmp00_65_41;
	wire [WIDTH*2-1+0:0] tmp00_65_42;
	wire [WIDTH*2-1+0:0] tmp00_65_43;
	wire [WIDTH*2-1+0:0] tmp00_65_44;
	wire [WIDTH*2-1+0:0] tmp00_65_45;
	wire [WIDTH*2-1+0:0] tmp00_65_46;
	wire [WIDTH*2-1+0:0] tmp00_65_47;
	wire [WIDTH*2-1+0:0] tmp00_65_48;
	wire [WIDTH*2-1+0:0] tmp00_65_49;
	wire [WIDTH*2-1+0:0] tmp00_65_50;
	wire [WIDTH*2-1+0:0] tmp00_65_51;
	wire [WIDTH*2-1+0:0] tmp00_65_52;
	wire [WIDTH*2-1+0:0] tmp00_65_53;
	wire [WIDTH*2-1+0:0] tmp00_65_54;
	wire [WIDTH*2-1+0:0] tmp00_65_55;
	wire [WIDTH*2-1+0:0] tmp00_65_56;
	wire [WIDTH*2-1+0:0] tmp00_65_57;
	wire [WIDTH*2-1+0:0] tmp00_65_58;
	wire [WIDTH*2-1+0:0] tmp00_65_59;
	wire [WIDTH*2-1+0:0] tmp00_65_60;
	wire [WIDTH*2-1+0:0] tmp00_65_61;
	wire [WIDTH*2-1+0:0] tmp00_65_62;
	wire [WIDTH*2-1+0:0] tmp00_65_63;
	wire [WIDTH*2-1+0:0] tmp00_65_64;
	wire [WIDTH*2-1+0:0] tmp00_65_65;
	wire [WIDTH*2-1+0:0] tmp00_65_66;
	wire [WIDTH*2-1+0:0] tmp00_65_67;
	wire [WIDTH*2-1+0:0] tmp00_65_68;
	wire [WIDTH*2-1+0:0] tmp00_65_69;
	wire [WIDTH*2-1+0:0] tmp00_65_70;
	wire [WIDTH*2-1+0:0] tmp00_65_71;
	wire [WIDTH*2-1+0:0] tmp00_65_72;
	wire [WIDTH*2-1+0:0] tmp00_65_73;
	wire [WIDTH*2-1+0:0] tmp00_65_74;
	wire [WIDTH*2-1+0:0] tmp00_65_75;
	wire [WIDTH*2-1+0:0] tmp00_65_76;
	wire [WIDTH*2-1+0:0] tmp00_65_77;
	wire [WIDTH*2-1+0:0] tmp00_65_78;
	wire [WIDTH*2-1+0:0] tmp00_65_79;
	wire [WIDTH*2-1+0:0] tmp00_65_80;
	wire [WIDTH*2-1+0:0] tmp00_65_81;
	wire [WIDTH*2-1+0:0] tmp00_65_82;
	wire [WIDTH*2-1+0:0] tmp00_65_83;
	wire [WIDTH*2-1+0:0] tmp00_66_0;
	wire [WIDTH*2-1+0:0] tmp00_66_1;
	wire [WIDTH*2-1+0:0] tmp00_66_2;
	wire [WIDTH*2-1+0:0] tmp00_66_3;
	wire [WIDTH*2-1+0:0] tmp00_66_4;
	wire [WIDTH*2-1+0:0] tmp00_66_5;
	wire [WIDTH*2-1+0:0] tmp00_66_6;
	wire [WIDTH*2-1+0:0] tmp00_66_7;
	wire [WIDTH*2-1+0:0] tmp00_66_8;
	wire [WIDTH*2-1+0:0] tmp00_66_9;
	wire [WIDTH*2-1+0:0] tmp00_66_10;
	wire [WIDTH*2-1+0:0] tmp00_66_11;
	wire [WIDTH*2-1+0:0] tmp00_66_12;
	wire [WIDTH*2-1+0:0] tmp00_66_13;
	wire [WIDTH*2-1+0:0] tmp00_66_14;
	wire [WIDTH*2-1+0:0] tmp00_66_15;
	wire [WIDTH*2-1+0:0] tmp00_66_16;
	wire [WIDTH*2-1+0:0] tmp00_66_17;
	wire [WIDTH*2-1+0:0] tmp00_66_18;
	wire [WIDTH*2-1+0:0] tmp00_66_19;
	wire [WIDTH*2-1+0:0] tmp00_66_20;
	wire [WIDTH*2-1+0:0] tmp00_66_21;
	wire [WIDTH*2-1+0:0] tmp00_66_22;
	wire [WIDTH*2-1+0:0] tmp00_66_23;
	wire [WIDTH*2-1+0:0] tmp00_66_24;
	wire [WIDTH*2-1+0:0] tmp00_66_25;
	wire [WIDTH*2-1+0:0] tmp00_66_26;
	wire [WIDTH*2-1+0:0] tmp00_66_27;
	wire [WIDTH*2-1+0:0] tmp00_66_28;
	wire [WIDTH*2-1+0:0] tmp00_66_29;
	wire [WIDTH*2-1+0:0] tmp00_66_30;
	wire [WIDTH*2-1+0:0] tmp00_66_31;
	wire [WIDTH*2-1+0:0] tmp00_66_32;
	wire [WIDTH*2-1+0:0] tmp00_66_33;
	wire [WIDTH*2-1+0:0] tmp00_66_34;
	wire [WIDTH*2-1+0:0] tmp00_66_35;
	wire [WIDTH*2-1+0:0] tmp00_66_36;
	wire [WIDTH*2-1+0:0] tmp00_66_37;
	wire [WIDTH*2-1+0:0] tmp00_66_38;
	wire [WIDTH*2-1+0:0] tmp00_66_39;
	wire [WIDTH*2-1+0:0] tmp00_66_40;
	wire [WIDTH*2-1+0:0] tmp00_66_41;
	wire [WIDTH*2-1+0:0] tmp00_66_42;
	wire [WIDTH*2-1+0:0] tmp00_66_43;
	wire [WIDTH*2-1+0:0] tmp00_66_44;
	wire [WIDTH*2-1+0:0] tmp00_66_45;
	wire [WIDTH*2-1+0:0] tmp00_66_46;
	wire [WIDTH*2-1+0:0] tmp00_66_47;
	wire [WIDTH*2-1+0:0] tmp00_66_48;
	wire [WIDTH*2-1+0:0] tmp00_66_49;
	wire [WIDTH*2-1+0:0] tmp00_66_50;
	wire [WIDTH*2-1+0:0] tmp00_66_51;
	wire [WIDTH*2-1+0:0] tmp00_66_52;
	wire [WIDTH*2-1+0:0] tmp00_66_53;
	wire [WIDTH*2-1+0:0] tmp00_66_54;
	wire [WIDTH*2-1+0:0] tmp00_66_55;
	wire [WIDTH*2-1+0:0] tmp00_66_56;
	wire [WIDTH*2-1+0:0] tmp00_66_57;
	wire [WIDTH*2-1+0:0] tmp00_66_58;
	wire [WIDTH*2-1+0:0] tmp00_66_59;
	wire [WIDTH*2-1+0:0] tmp00_66_60;
	wire [WIDTH*2-1+0:0] tmp00_66_61;
	wire [WIDTH*2-1+0:0] tmp00_66_62;
	wire [WIDTH*2-1+0:0] tmp00_66_63;
	wire [WIDTH*2-1+0:0] tmp00_66_64;
	wire [WIDTH*2-1+0:0] tmp00_66_65;
	wire [WIDTH*2-1+0:0] tmp00_66_66;
	wire [WIDTH*2-1+0:0] tmp00_66_67;
	wire [WIDTH*2-1+0:0] tmp00_66_68;
	wire [WIDTH*2-1+0:0] tmp00_66_69;
	wire [WIDTH*2-1+0:0] tmp00_66_70;
	wire [WIDTH*2-1+0:0] tmp00_66_71;
	wire [WIDTH*2-1+0:0] tmp00_66_72;
	wire [WIDTH*2-1+0:0] tmp00_66_73;
	wire [WIDTH*2-1+0:0] tmp00_66_74;
	wire [WIDTH*2-1+0:0] tmp00_66_75;
	wire [WIDTH*2-1+0:0] tmp00_66_76;
	wire [WIDTH*2-1+0:0] tmp00_66_77;
	wire [WIDTH*2-1+0:0] tmp00_66_78;
	wire [WIDTH*2-1+0:0] tmp00_66_79;
	wire [WIDTH*2-1+0:0] tmp00_66_80;
	wire [WIDTH*2-1+0:0] tmp00_66_81;
	wire [WIDTH*2-1+0:0] tmp00_66_82;
	wire [WIDTH*2-1+0:0] tmp00_66_83;
	wire [WIDTH*2-1+0:0] tmp00_67_0;
	wire [WIDTH*2-1+0:0] tmp00_67_1;
	wire [WIDTH*2-1+0:0] tmp00_67_2;
	wire [WIDTH*2-1+0:0] tmp00_67_3;
	wire [WIDTH*2-1+0:0] tmp00_67_4;
	wire [WIDTH*2-1+0:0] tmp00_67_5;
	wire [WIDTH*2-1+0:0] tmp00_67_6;
	wire [WIDTH*2-1+0:0] tmp00_67_7;
	wire [WIDTH*2-1+0:0] tmp00_67_8;
	wire [WIDTH*2-1+0:0] tmp00_67_9;
	wire [WIDTH*2-1+0:0] tmp00_67_10;
	wire [WIDTH*2-1+0:0] tmp00_67_11;
	wire [WIDTH*2-1+0:0] tmp00_67_12;
	wire [WIDTH*2-1+0:0] tmp00_67_13;
	wire [WIDTH*2-1+0:0] tmp00_67_14;
	wire [WIDTH*2-1+0:0] tmp00_67_15;
	wire [WIDTH*2-1+0:0] tmp00_67_16;
	wire [WIDTH*2-1+0:0] tmp00_67_17;
	wire [WIDTH*2-1+0:0] tmp00_67_18;
	wire [WIDTH*2-1+0:0] tmp00_67_19;
	wire [WIDTH*2-1+0:0] tmp00_67_20;
	wire [WIDTH*2-1+0:0] tmp00_67_21;
	wire [WIDTH*2-1+0:0] tmp00_67_22;
	wire [WIDTH*2-1+0:0] tmp00_67_23;
	wire [WIDTH*2-1+0:0] tmp00_67_24;
	wire [WIDTH*2-1+0:0] tmp00_67_25;
	wire [WIDTH*2-1+0:0] tmp00_67_26;
	wire [WIDTH*2-1+0:0] tmp00_67_27;
	wire [WIDTH*2-1+0:0] tmp00_67_28;
	wire [WIDTH*2-1+0:0] tmp00_67_29;
	wire [WIDTH*2-1+0:0] tmp00_67_30;
	wire [WIDTH*2-1+0:0] tmp00_67_31;
	wire [WIDTH*2-1+0:0] tmp00_67_32;
	wire [WIDTH*2-1+0:0] tmp00_67_33;
	wire [WIDTH*2-1+0:0] tmp00_67_34;
	wire [WIDTH*2-1+0:0] tmp00_67_35;
	wire [WIDTH*2-1+0:0] tmp00_67_36;
	wire [WIDTH*2-1+0:0] tmp00_67_37;
	wire [WIDTH*2-1+0:0] tmp00_67_38;
	wire [WIDTH*2-1+0:0] tmp00_67_39;
	wire [WIDTH*2-1+0:0] tmp00_67_40;
	wire [WIDTH*2-1+0:0] tmp00_67_41;
	wire [WIDTH*2-1+0:0] tmp00_67_42;
	wire [WIDTH*2-1+0:0] tmp00_67_43;
	wire [WIDTH*2-1+0:0] tmp00_67_44;
	wire [WIDTH*2-1+0:0] tmp00_67_45;
	wire [WIDTH*2-1+0:0] tmp00_67_46;
	wire [WIDTH*2-1+0:0] tmp00_67_47;
	wire [WIDTH*2-1+0:0] tmp00_67_48;
	wire [WIDTH*2-1+0:0] tmp00_67_49;
	wire [WIDTH*2-1+0:0] tmp00_67_50;
	wire [WIDTH*2-1+0:0] tmp00_67_51;
	wire [WIDTH*2-1+0:0] tmp00_67_52;
	wire [WIDTH*2-1+0:0] tmp00_67_53;
	wire [WIDTH*2-1+0:0] tmp00_67_54;
	wire [WIDTH*2-1+0:0] tmp00_67_55;
	wire [WIDTH*2-1+0:0] tmp00_67_56;
	wire [WIDTH*2-1+0:0] tmp00_67_57;
	wire [WIDTH*2-1+0:0] tmp00_67_58;
	wire [WIDTH*2-1+0:0] tmp00_67_59;
	wire [WIDTH*2-1+0:0] tmp00_67_60;
	wire [WIDTH*2-1+0:0] tmp00_67_61;
	wire [WIDTH*2-1+0:0] tmp00_67_62;
	wire [WIDTH*2-1+0:0] tmp00_67_63;
	wire [WIDTH*2-1+0:0] tmp00_67_64;
	wire [WIDTH*2-1+0:0] tmp00_67_65;
	wire [WIDTH*2-1+0:0] tmp00_67_66;
	wire [WIDTH*2-1+0:0] tmp00_67_67;
	wire [WIDTH*2-1+0:0] tmp00_67_68;
	wire [WIDTH*2-1+0:0] tmp00_67_69;
	wire [WIDTH*2-1+0:0] tmp00_67_70;
	wire [WIDTH*2-1+0:0] tmp00_67_71;
	wire [WIDTH*2-1+0:0] tmp00_67_72;
	wire [WIDTH*2-1+0:0] tmp00_67_73;
	wire [WIDTH*2-1+0:0] tmp00_67_74;
	wire [WIDTH*2-1+0:0] tmp00_67_75;
	wire [WIDTH*2-1+0:0] tmp00_67_76;
	wire [WIDTH*2-1+0:0] tmp00_67_77;
	wire [WIDTH*2-1+0:0] tmp00_67_78;
	wire [WIDTH*2-1+0:0] tmp00_67_79;
	wire [WIDTH*2-1+0:0] tmp00_67_80;
	wire [WIDTH*2-1+0:0] tmp00_67_81;
	wire [WIDTH*2-1+0:0] tmp00_67_82;
	wire [WIDTH*2-1+0:0] tmp00_67_83;
	wire [WIDTH*2-1+0:0] tmp00_68_0;
	wire [WIDTH*2-1+0:0] tmp00_68_1;
	wire [WIDTH*2-1+0:0] tmp00_68_2;
	wire [WIDTH*2-1+0:0] tmp00_68_3;
	wire [WIDTH*2-1+0:0] tmp00_68_4;
	wire [WIDTH*2-1+0:0] tmp00_68_5;
	wire [WIDTH*2-1+0:0] tmp00_68_6;
	wire [WIDTH*2-1+0:0] tmp00_68_7;
	wire [WIDTH*2-1+0:0] tmp00_68_8;
	wire [WIDTH*2-1+0:0] tmp00_68_9;
	wire [WIDTH*2-1+0:0] tmp00_68_10;
	wire [WIDTH*2-1+0:0] tmp00_68_11;
	wire [WIDTH*2-1+0:0] tmp00_68_12;
	wire [WIDTH*2-1+0:0] tmp00_68_13;
	wire [WIDTH*2-1+0:0] tmp00_68_14;
	wire [WIDTH*2-1+0:0] tmp00_68_15;
	wire [WIDTH*2-1+0:0] tmp00_68_16;
	wire [WIDTH*2-1+0:0] tmp00_68_17;
	wire [WIDTH*2-1+0:0] tmp00_68_18;
	wire [WIDTH*2-1+0:0] tmp00_68_19;
	wire [WIDTH*2-1+0:0] tmp00_68_20;
	wire [WIDTH*2-1+0:0] tmp00_68_21;
	wire [WIDTH*2-1+0:0] tmp00_68_22;
	wire [WIDTH*2-1+0:0] tmp00_68_23;
	wire [WIDTH*2-1+0:0] tmp00_68_24;
	wire [WIDTH*2-1+0:0] tmp00_68_25;
	wire [WIDTH*2-1+0:0] tmp00_68_26;
	wire [WIDTH*2-1+0:0] tmp00_68_27;
	wire [WIDTH*2-1+0:0] tmp00_68_28;
	wire [WIDTH*2-1+0:0] tmp00_68_29;
	wire [WIDTH*2-1+0:0] tmp00_68_30;
	wire [WIDTH*2-1+0:0] tmp00_68_31;
	wire [WIDTH*2-1+0:0] tmp00_68_32;
	wire [WIDTH*2-1+0:0] tmp00_68_33;
	wire [WIDTH*2-1+0:0] tmp00_68_34;
	wire [WIDTH*2-1+0:0] tmp00_68_35;
	wire [WIDTH*2-1+0:0] tmp00_68_36;
	wire [WIDTH*2-1+0:0] tmp00_68_37;
	wire [WIDTH*2-1+0:0] tmp00_68_38;
	wire [WIDTH*2-1+0:0] tmp00_68_39;
	wire [WIDTH*2-1+0:0] tmp00_68_40;
	wire [WIDTH*2-1+0:0] tmp00_68_41;
	wire [WIDTH*2-1+0:0] tmp00_68_42;
	wire [WIDTH*2-1+0:0] tmp00_68_43;
	wire [WIDTH*2-1+0:0] tmp00_68_44;
	wire [WIDTH*2-1+0:0] tmp00_68_45;
	wire [WIDTH*2-1+0:0] tmp00_68_46;
	wire [WIDTH*2-1+0:0] tmp00_68_47;
	wire [WIDTH*2-1+0:0] tmp00_68_48;
	wire [WIDTH*2-1+0:0] tmp00_68_49;
	wire [WIDTH*2-1+0:0] tmp00_68_50;
	wire [WIDTH*2-1+0:0] tmp00_68_51;
	wire [WIDTH*2-1+0:0] tmp00_68_52;
	wire [WIDTH*2-1+0:0] tmp00_68_53;
	wire [WIDTH*2-1+0:0] tmp00_68_54;
	wire [WIDTH*2-1+0:0] tmp00_68_55;
	wire [WIDTH*2-1+0:0] tmp00_68_56;
	wire [WIDTH*2-1+0:0] tmp00_68_57;
	wire [WIDTH*2-1+0:0] tmp00_68_58;
	wire [WIDTH*2-1+0:0] tmp00_68_59;
	wire [WIDTH*2-1+0:0] tmp00_68_60;
	wire [WIDTH*2-1+0:0] tmp00_68_61;
	wire [WIDTH*2-1+0:0] tmp00_68_62;
	wire [WIDTH*2-1+0:0] tmp00_68_63;
	wire [WIDTH*2-1+0:0] tmp00_68_64;
	wire [WIDTH*2-1+0:0] tmp00_68_65;
	wire [WIDTH*2-1+0:0] tmp00_68_66;
	wire [WIDTH*2-1+0:0] tmp00_68_67;
	wire [WIDTH*2-1+0:0] tmp00_68_68;
	wire [WIDTH*2-1+0:0] tmp00_68_69;
	wire [WIDTH*2-1+0:0] tmp00_68_70;
	wire [WIDTH*2-1+0:0] tmp00_68_71;
	wire [WIDTH*2-1+0:0] tmp00_68_72;
	wire [WIDTH*2-1+0:0] tmp00_68_73;
	wire [WIDTH*2-1+0:0] tmp00_68_74;
	wire [WIDTH*2-1+0:0] tmp00_68_75;
	wire [WIDTH*2-1+0:0] tmp00_68_76;
	wire [WIDTH*2-1+0:0] tmp00_68_77;
	wire [WIDTH*2-1+0:0] tmp00_68_78;
	wire [WIDTH*2-1+0:0] tmp00_68_79;
	wire [WIDTH*2-1+0:0] tmp00_68_80;
	wire [WIDTH*2-1+0:0] tmp00_68_81;
	wire [WIDTH*2-1+0:0] tmp00_68_82;
	wire [WIDTH*2-1+0:0] tmp00_68_83;
	wire [WIDTH*2-1+0:0] tmp00_69_0;
	wire [WIDTH*2-1+0:0] tmp00_69_1;
	wire [WIDTH*2-1+0:0] tmp00_69_2;
	wire [WIDTH*2-1+0:0] tmp00_69_3;
	wire [WIDTH*2-1+0:0] tmp00_69_4;
	wire [WIDTH*2-1+0:0] tmp00_69_5;
	wire [WIDTH*2-1+0:0] tmp00_69_6;
	wire [WIDTH*2-1+0:0] tmp00_69_7;
	wire [WIDTH*2-1+0:0] tmp00_69_8;
	wire [WIDTH*2-1+0:0] tmp00_69_9;
	wire [WIDTH*2-1+0:0] tmp00_69_10;
	wire [WIDTH*2-1+0:0] tmp00_69_11;
	wire [WIDTH*2-1+0:0] tmp00_69_12;
	wire [WIDTH*2-1+0:0] tmp00_69_13;
	wire [WIDTH*2-1+0:0] tmp00_69_14;
	wire [WIDTH*2-1+0:0] tmp00_69_15;
	wire [WIDTH*2-1+0:0] tmp00_69_16;
	wire [WIDTH*2-1+0:0] tmp00_69_17;
	wire [WIDTH*2-1+0:0] tmp00_69_18;
	wire [WIDTH*2-1+0:0] tmp00_69_19;
	wire [WIDTH*2-1+0:0] tmp00_69_20;
	wire [WIDTH*2-1+0:0] tmp00_69_21;
	wire [WIDTH*2-1+0:0] tmp00_69_22;
	wire [WIDTH*2-1+0:0] tmp00_69_23;
	wire [WIDTH*2-1+0:0] tmp00_69_24;
	wire [WIDTH*2-1+0:0] tmp00_69_25;
	wire [WIDTH*2-1+0:0] tmp00_69_26;
	wire [WIDTH*2-1+0:0] tmp00_69_27;
	wire [WIDTH*2-1+0:0] tmp00_69_28;
	wire [WIDTH*2-1+0:0] tmp00_69_29;
	wire [WIDTH*2-1+0:0] tmp00_69_30;
	wire [WIDTH*2-1+0:0] tmp00_69_31;
	wire [WIDTH*2-1+0:0] tmp00_69_32;
	wire [WIDTH*2-1+0:0] tmp00_69_33;
	wire [WIDTH*2-1+0:0] tmp00_69_34;
	wire [WIDTH*2-1+0:0] tmp00_69_35;
	wire [WIDTH*2-1+0:0] tmp00_69_36;
	wire [WIDTH*2-1+0:0] tmp00_69_37;
	wire [WIDTH*2-1+0:0] tmp00_69_38;
	wire [WIDTH*2-1+0:0] tmp00_69_39;
	wire [WIDTH*2-1+0:0] tmp00_69_40;
	wire [WIDTH*2-1+0:0] tmp00_69_41;
	wire [WIDTH*2-1+0:0] tmp00_69_42;
	wire [WIDTH*2-1+0:0] tmp00_69_43;
	wire [WIDTH*2-1+0:0] tmp00_69_44;
	wire [WIDTH*2-1+0:0] tmp00_69_45;
	wire [WIDTH*2-1+0:0] tmp00_69_46;
	wire [WIDTH*2-1+0:0] tmp00_69_47;
	wire [WIDTH*2-1+0:0] tmp00_69_48;
	wire [WIDTH*2-1+0:0] tmp00_69_49;
	wire [WIDTH*2-1+0:0] tmp00_69_50;
	wire [WIDTH*2-1+0:0] tmp00_69_51;
	wire [WIDTH*2-1+0:0] tmp00_69_52;
	wire [WIDTH*2-1+0:0] tmp00_69_53;
	wire [WIDTH*2-1+0:0] tmp00_69_54;
	wire [WIDTH*2-1+0:0] tmp00_69_55;
	wire [WIDTH*2-1+0:0] tmp00_69_56;
	wire [WIDTH*2-1+0:0] tmp00_69_57;
	wire [WIDTH*2-1+0:0] tmp00_69_58;
	wire [WIDTH*2-1+0:0] tmp00_69_59;
	wire [WIDTH*2-1+0:0] tmp00_69_60;
	wire [WIDTH*2-1+0:0] tmp00_69_61;
	wire [WIDTH*2-1+0:0] tmp00_69_62;
	wire [WIDTH*2-1+0:0] tmp00_69_63;
	wire [WIDTH*2-1+0:0] tmp00_69_64;
	wire [WIDTH*2-1+0:0] tmp00_69_65;
	wire [WIDTH*2-1+0:0] tmp00_69_66;
	wire [WIDTH*2-1+0:0] tmp00_69_67;
	wire [WIDTH*2-1+0:0] tmp00_69_68;
	wire [WIDTH*2-1+0:0] tmp00_69_69;
	wire [WIDTH*2-1+0:0] tmp00_69_70;
	wire [WIDTH*2-1+0:0] tmp00_69_71;
	wire [WIDTH*2-1+0:0] tmp00_69_72;
	wire [WIDTH*2-1+0:0] tmp00_69_73;
	wire [WIDTH*2-1+0:0] tmp00_69_74;
	wire [WIDTH*2-1+0:0] tmp00_69_75;
	wire [WIDTH*2-1+0:0] tmp00_69_76;
	wire [WIDTH*2-1+0:0] tmp00_69_77;
	wire [WIDTH*2-1+0:0] tmp00_69_78;
	wire [WIDTH*2-1+0:0] tmp00_69_79;
	wire [WIDTH*2-1+0:0] tmp00_69_80;
	wire [WIDTH*2-1+0:0] tmp00_69_81;
	wire [WIDTH*2-1+0:0] tmp00_69_82;
	wire [WIDTH*2-1+0:0] tmp00_69_83;
	wire [WIDTH*2-1+0:0] tmp00_70_0;
	wire [WIDTH*2-1+0:0] tmp00_70_1;
	wire [WIDTH*2-1+0:0] tmp00_70_2;
	wire [WIDTH*2-1+0:0] tmp00_70_3;
	wire [WIDTH*2-1+0:0] tmp00_70_4;
	wire [WIDTH*2-1+0:0] tmp00_70_5;
	wire [WIDTH*2-1+0:0] tmp00_70_6;
	wire [WIDTH*2-1+0:0] tmp00_70_7;
	wire [WIDTH*2-1+0:0] tmp00_70_8;
	wire [WIDTH*2-1+0:0] tmp00_70_9;
	wire [WIDTH*2-1+0:0] tmp00_70_10;
	wire [WIDTH*2-1+0:0] tmp00_70_11;
	wire [WIDTH*2-1+0:0] tmp00_70_12;
	wire [WIDTH*2-1+0:0] tmp00_70_13;
	wire [WIDTH*2-1+0:0] tmp00_70_14;
	wire [WIDTH*2-1+0:0] tmp00_70_15;
	wire [WIDTH*2-1+0:0] tmp00_70_16;
	wire [WIDTH*2-1+0:0] tmp00_70_17;
	wire [WIDTH*2-1+0:0] tmp00_70_18;
	wire [WIDTH*2-1+0:0] tmp00_70_19;
	wire [WIDTH*2-1+0:0] tmp00_70_20;
	wire [WIDTH*2-1+0:0] tmp00_70_21;
	wire [WIDTH*2-1+0:0] tmp00_70_22;
	wire [WIDTH*2-1+0:0] tmp00_70_23;
	wire [WIDTH*2-1+0:0] tmp00_70_24;
	wire [WIDTH*2-1+0:0] tmp00_70_25;
	wire [WIDTH*2-1+0:0] tmp00_70_26;
	wire [WIDTH*2-1+0:0] tmp00_70_27;
	wire [WIDTH*2-1+0:0] tmp00_70_28;
	wire [WIDTH*2-1+0:0] tmp00_70_29;
	wire [WIDTH*2-1+0:0] tmp00_70_30;
	wire [WIDTH*2-1+0:0] tmp00_70_31;
	wire [WIDTH*2-1+0:0] tmp00_70_32;
	wire [WIDTH*2-1+0:0] tmp00_70_33;
	wire [WIDTH*2-1+0:0] tmp00_70_34;
	wire [WIDTH*2-1+0:0] tmp00_70_35;
	wire [WIDTH*2-1+0:0] tmp00_70_36;
	wire [WIDTH*2-1+0:0] tmp00_70_37;
	wire [WIDTH*2-1+0:0] tmp00_70_38;
	wire [WIDTH*2-1+0:0] tmp00_70_39;
	wire [WIDTH*2-1+0:0] tmp00_70_40;
	wire [WIDTH*2-1+0:0] tmp00_70_41;
	wire [WIDTH*2-1+0:0] tmp00_70_42;
	wire [WIDTH*2-1+0:0] tmp00_70_43;
	wire [WIDTH*2-1+0:0] tmp00_70_44;
	wire [WIDTH*2-1+0:0] tmp00_70_45;
	wire [WIDTH*2-1+0:0] tmp00_70_46;
	wire [WIDTH*2-1+0:0] tmp00_70_47;
	wire [WIDTH*2-1+0:0] tmp00_70_48;
	wire [WIDTH*2-1+0:0] tmp00_70_49;
	wire [WIDTH*2-1+0:0] tmp00_70_50;
	wire [WIDTH*2-1+0:0] tmp00_70_51;
	wire [WIDTH*2-1+0:0] tmp00_70_52;
	wire [WIDTH*2-1+0:0] tmp00_70_53;
	wire [WIDTH*2-1+0:0] tmp00_70_54;
	wire [WIDTH*2-1+0:0] tmp00_70_55;
	wire [WIDTH*2-1+0:0] tmp00_70_56;
	wire [WIDTH*2-1+0:0] tmp00_70_57;
	wire [WIDTH*2-1+0:0] tmp00_70_58;
	wire [WIDTH*2-1+0:0] tmp00_70_59;
	wire [WIDTH*2-1+0:0] tmp00_70_60;
	wire [WIDTH*2-1+0:0] tmp00_70_61;
	wire [WIDTH*2-1+0:0] tmp00_70_62;
	wire [WIDTH*2-1+0:0] tmp00_70_63;
	wire [WIDTH*2-1+0:0] tmp00_70_64;
	wire [WIDTH*2-1+0:0] tmp00_70_65;
	wire [WIDTH*2-1+0:0] tmp00_70_66;
	wire [WIDTH*2-1+0:0] tmp00_70_67;
	wire [WIDTH*2-1+0:0] tmp00_70_68;
	wire [WIDTH*2-1+0:0] tmp00_70_69;
	wire [WIDTH*2-1+0:0] tmp00_70_70;
	wire [WIDTH*2-1+0:0] tmp00_70_71;
	wire [WIDTH*2-1+0:0] tmp00_70_72;
	wire [WIDTH*2-1+0:0] tmp00_70_73;
	wire [WIDTH*2-1+0:0] tmp00_70_74;
	wire [WIDTH*2-1+0:0] tmp00_70_75;
	wire [WIDTH*2-1+0:0] tmp00_70_76;
	wire [WIDTH*2-1+0:0] tmp00_70_77;
	wire [WIDTH*2-1+0:0] tmp00_70_78;
	wire [WIDTH*2-1+0:0] tmp00_70_79;
	wire [WIDTH*2-1+0:0] tmp00_70_80;
	wire [WIDTH*2-1+0:0] tmp00_70_81;
	wire [WIDTH*2-1+0:0] tmp00_70_82;
	wire [WIDTH*2-1+0:0] tmp00_70_83;
	wire [WIDTH*2-1+0:0] tmp00_71_0;
	wire [WIDTH*2-1+0:0] tmp00_71_1;
	wire [WIDTH*2-1+0:0] tmp00_71_2;
	wire [WIDTH*2-1+0:0] tmp00_71_3;
	wire [WIDTH*2-1+0:0] tmp00_71_4;
	wire [WIDTH*2-1+0:0] tmp00_71_5;
	wire [WIDTH*2-1+0:0] tmp00_71_6;
	wire [WIDTH*2-1+0:0] tmp00_71_7;
	wire [WIDTH*2-1+0:0] tmp00_71_8;
	wire [WIDTH*2-1+0:0] tmp00_71_9;
	wire [WIDTH*2-1+0:0] tmp00_71_10;
	wire [WIDTH*2-1+0:0] tmp00_71_11;
	wire [WIDTH*2-1+0:0] tmp00_71_12;
	wire [WIDTH*2-1+0:0] tmp00_71_13;
	wire [WIDTH*2-1+0:0] tmp00_71_14;
	wire [WIDTH*2-1+0:0] tmp00_71_15;
	wire [WIDTH*2-1+0:0] tmp00_71_16;
	wire [WIDTH*2-1+0:0] tmp00_71_17;
	wire [WIDTH*2-1+0:0] tmp00_71_18;
	wire [WIDTH*2-1+0:0] tmp00_71_19;
	wire [WIDTH*2-1+0:0] tmp00_71_20;
	wire [WIDTH*2-1+0:0] tmp00_71_21;
	wire [WIDTH*2-1+0:0] tmp00_71_22;
	wire [WIDTH*2-1+0:0] tmp00_71_23;
	wire [WIDTH*2-1+0:0] tmp00_71_24;
	wire [WIDTH*2-1+0:0] tmp00_71_25;
	wire [WIDTH*2-1+0:0] tmp00_71_26;
	wire [WIDTH*2-1+0:0] tmp00_71_27;
	wire [WIDTH*2-1+0:0] tmp00_71_28;
	wire [WIDTH*2-1+0:0] tmp00_71_29;
	wire [WIDTH*2-1+0:0] tmp00_71_30;
	wire [WIDTH*2-1+0:0] tmp00_71_31;
	wire [WIDTH*2-1+0:0] tmp00_71_32;
	wire [WIDTH*2-1+0:0] tmp00_71_33;
	wire [WIDTH*2-1+0:0] tmp00_71_34;
	wire [WIDTH*2-1+0:0] tmp00_71_35;
	wire [WIDTH*2-1+0:0] tmp00_71_36;
	wire [WIDTH*2-1+0:0] tmp00_71_37;
	wire [WIDTH*2-1+0:0] tmp00_71_38;
	wire [WIDTH*2-1+0:0] tmp00_71_39;
	wire [WIDTH*2-1+0:0] tmp00_71_40;
	wire [WIDTH*2-1+0:0] tmp00_71_41;
	wire [WIDTH*2-1+0:0] tmp00_71_42;
	wire [WIDTH*2-1+0:0] tmp00_71_43;
	wire [WIDTH*2-1+0:0] tmp00_71_44;
	wire [WIDTH*2-1+0:0] tmp00_71_45;
	wire [WIDTH*2-1+0:0] tmp00_71_46;
	wire [WIDTH*2-1+0:0] tmp00_71_47;
	wire [WIDTH*2-1+0:0] tmp00_71_48;
	wire [WIDTH*2-1+0:0] tmp00_71_49;
	wire [WIDTH*2-1+0:0] tmp00_71_50;
	wire [WIDTH*2-1+0:0] tmp00_71_51;
	wire [WIDTH*2-1+0:0] tmp00_71_52;
	wire [WIDTH*2-1+0:0] tmp00_71_53;
	wire [WIDTH*2-1+0:0] tmp00_71_54;
	wire [WIDTH*2-1+0:0] tmp00_71_55;
	wire [WIDTH*2-1+0:0] tmp00_71_56;
	wire [WIDTH*2-1+0:0] tmp00_71_57;
	wire [WIDTH*2-1+0:0] tmp00_71_58;
	wire [WIDTH*2-1+0:0] tmp00_71_59;
	wire [WIDTH*2-1+0:0] tmp00_71_60;
	wire [WIDTH*2-1+0:0] tmp00_71_61;
	wire [WIDTH*2-1+0:0] tmp00_71_62;
	wire [WIDTH*2-1+0:0] tmp00_71_63;
	wire [WIDTH*2-1+0:0] tmp00_71_64;
	wire [WIDTH*2-1+0:0] tmp00_71_65;
	wire [WIDTH*2-1+0:0] tmp00_71_66;
	wire [WIDTH*2-1+0:0] tmp00_71_67;
	wire [WIDTH*2-1+0:0] tmp00_71_68;
	wire [WIDTH*2-1+0:0] tmp00_71_69;
	wire [WIDTH*2-1+0:0] tmp00_71_70;
	wire [WIDTH*2-1+0:0] tmp00_71_71;
	wire [WIDTH*2-1+0:0] tmp00_71_72;
	wire [WIDTH*2-1+0:0] tmp00_71_73;
	wire [WIDTH*2-1+0:0] tmp00_71_74;
	wire [WIDTH*2-1+0:0] tmp00_71_75;
	wire [WIDTH*2-1+0:0] tmp00_71_76;
	wire [WIDTH*2-1+0:0] tmp00_71_77;
	wire [WIDTH*2-1+0:0] tmp00_71_78;
	wire [WIDTH*2-1+0:0] tmp00_71_79;
	wire [WIDTH*2-1+0:0] tmp00_71_80;
	wire [WIDTH*2-1+0:0] tmp00_71_81;
	wire [WIDTH*2-1+0:0] tmp00_71_82;
	wire [WIDTH*2-1+0:0] tmp00_71_83;
	wire [WIDTH*2-1+0:0] tmp00_72_0;
	wire [WIDTH*2-1+0:0] tmp00_72_1;
	wire [WIDTH*2-1+0:0] tmp00_72_2;
	wire [WIDTH*2-1+0:0] tmp00_72_3;
	wire [WIDTH*2-1+0:0] tmp00_72_4;
	wire [WIDTH*2-1+0:0] tmp00_72_5;
	wire [WIDTH*2-1+0:0] tmp00_72_6;
	wire [WIDTH*2-1+0:0] tmp00_72_7;
	wire [WIDTH*2-1+0:0] tmp00_72_8;
	wire [WIDTH*2-1+0:0] tmp00_72_9;
	wire [WIDTH*2-1+0:0] tmp00_72_10;
	wire [WIDTH*2-1+0:0] tmp00_72_11;
	wire [WIDTH*2-1+0:0] tmp00_72_12;
	wire [WIDTH*2-1+0:0] tmp00_72_13;
	wire [WIDTH*2-1+0:0] tmp00_72_14;
	wire [WIDTH*2-1+0:0] tmp00_72_15;
	wire [WIDTH*2-1+0:0] tmp00_72_16;
	wire [WIDTH*2-1+0:0] tmp00_72_17;
	wire [WIDTH*2-1+0:0] tmp00_72_18;
	wire [WIDTH*2-1+0:0] tmp00_72_19;
	wire [WIDTH*2-1+0:0] tmp00_72_20;
	wire [WIDTH*2-1+0:0] tmp00_72_21;
	wire [WIDTH*2-1+0:0] tmp00_72_22;
	wire [WIDTH*2-1+0:0] tmp00_72_23;
	wire [WIDTH*2-1+0:0] tmp00_72_24;
	wire [WIDTH*2-1+0:0] tmp00_72_25;
	wire [WIDTH*2-1+0:0] tmp00_72_26;
	wire [WIDTH*2-1+0:0] tmp00_72_27;
	wire [WIDTH*2-1+0:0] tmp00_72_28;
	wire [WIDTH*2-1+0:0] tmp00_72_29;
	wire [WIDTH*2-1+0:0] tmp00_72_30;
	wire [WIDTH*2-1+0:0] tmp00_72_31;
	wire [WIDTH*2-1+0:0] tmp00_72_32;
	wire [WIDTH*2-1+0:0] tmp00_72_33;
	wire [WIDTH*2-1+0:0] tmp00_72_34;
	wire [WIDTH*2-1+0:0] tmp00_72_35;
	wire [WIDTH*2-1+0:0] tmp00_72_36;
	wire [WIDTH*2-1+0:0] tmp00_72_37;
	wire [WIDTH*2-1+0:0] tmp00_72_38;
	wire [WIDTH*2-1+0:0] tmp00_72_39;
	wire [WIDTH*2-1+0:0] tmp00_72_40;
	wire [WIDTH*2-1+0:0] tmp00_72_41;
	wire [WIDTH*2-1+0:0] tmp00_72_42;
	wire [WIDTH*2-1+0:0] tmp00_72_43;
	wire [WIDTH*2-1+0:0] tmp00_72_44;
	wire [WIDTH*2-1+0:0] tmp00_72_45;
	wire [WIDTH*2-1+0:0] tmp00_72_46;
	wire [WIDTH*2-1+0:0] tmp00_72_47;
	wire [WIDTH*2-1+0:0] tmp00_72_48;
	wire [WIDTH*2-1+0:0] tmp00_72_49;
	wire [WIDTH*2-1+0:0] tmp00_72_50;
	wire [WIDTH*2-1+0:0] tmp00_72_51;
	wire [WIDTH*2-1+0:0] tmp00_72_52;
	wire [WIDTH*2-1+0:0] tmp00_72_53;
	wire [WIDTH*2-1+0:0] tmp00_72_54;
	wire [WIDTH*2-1+0:0] tmp00_72_55;
	wire [WIDTH*2-1+0:0] tmp00_72_56;
	wire [WIDTH*2-1+0:0] tmp00_72_57;
	wire [WIDTH*2-1+0:0] tmp00_72_58;
	wire [WIDTH*2-1+0:0] tmp00_72_59;
	wire [WIDTH*2-1+0:0] tmp00_72_60;
	wire [WIDTH*2-1+0:0] tmp00_72_61;
	wire [WIDTH*2-1+0:0] tmp00_72_62;
	wire [WIDTH*2-1+0:0] tmp00_72_63;
	wire [WIDTH*2-1+0:0] tmp00_72_64;
	wire [WIDTH*2-1+0:0] tmp00_72_65;
	wire [WIDTH*2-1+0:0] tmp00_72_66;
	wire [WIDTH*2-1+0:0] tmp00_72_67;
	wire [WIDTH*2-1+0:0] tmp00_72_68;
	wire [WIDTH*2-1+0:0] tmp00_72_69;
	wire [WIDTH*2-1+0:0] tmp00_72_70;
	wire [WIDTH*2-1+0:0] tmp00_72_71;
	wire [WIDTH*2-1+0:0] tmp00_72_72;
	wire [WIDTH*2-1+0:0] tmp00_72_73;
	wire [WIDTH*2-1+0:0] tmp00_72_74;
	wire [WIDTH*2-1+0:0] tmp00_72_75;
	wire [WIDTH*2-1+0:0] tmp00_72_76;
	wire [WIDTH*2-1+0:0] tmp00_72_77;
	wire [WIDTH*2-1+0:0] tmp00_72_78;
	wire [WIDTH*2-1+0:0] tmp00_72_79;
	wire [WIDTH*2-1+0:0] tmp00_72_80;
	wire [WIDTH*2-1+0:0] tmp00_72_81;
	wire [WIDTH*2-1+0:0] tmp00_72_82;
	wire [WIDTH*2-1+0:0] tmp00_72_83;
	wire [WIDTH*2-1+0:0] tmp00_73_0;
	wire [WIDTH*2-1+0:0] tmp00_73_1;
	wire [WIDTH*2-1+0:0] tmp00_73_2;
	wire [WIDTH*2-1+0:0] tmp00_73_3;
	wire [WIDTH*2-1+0:0] tmp00_73_4;
	wire [WIDTH*2-1+0:0] tmp00_73_5;
	wire [WIDTH*2-1+0:0] tmp00_73_6;
	wire [WIDTH*2-1+0:0] tmp00_73_7;
	wire [WIDTH*2-1+0:0] tmp00_73_8;
	wire [WIDTH*2-1+0:0] tmp00_73_9;
	wire [WIDTH*2-1+0:0] tmp00_73_10;
	wire [WIDTH*2-1+0:0] tmp00_73_11;
	wire [WIDTH*2-1+0:0] tmp00_73_12;
	wire [WIDTH*2-1+0:0] tmp00_73_13;
	wire [WIDTH*2-1+0:0] tmp00_73_14;
	wire [WIDTH*2-1+0:0] tmp00_73_15;
	wire [WIDTH*2-1+0:0] tmp00_73_16;
	wire [WIDTH*2-1+0:0] tmp00_73_17;
	wire [WIDTH*2-1+0:0] tmp00_73_18;
	wire [WIDTH*2-1+0:0] tmp00_73_19;
	wire [WIDTH*2-1+0:0] tmp00_73_20;
	wire [WIDTH*2-1+0:0] tmp00_73_21;
	wire [WIDTH*2-1+0:0] tmp00_73_22;
	wire [WIDTH*2-1+0:0] tmp00_73_23;
	wire [WIDTH*2-1+0:0] tmp00_73_24;
	wire [WIDTH*2-1+0:0] tmp00_73_25;
	wire [WIDTH*2-1+0:0] tmp00_73_26;
	wire [WIDTH*2-1+0:0] tmp00_73_27;
	wire [WIDTH*2-1+0:0] tmp00_73_28;
	wire [WIDTH*2-1+0:0] tmp00_73_29;
	wire [WIDTH*2-1+0:0] tmp00_73_30;
	wire [WIDTH*2-1+0:0] tmp00_73_31;
	wire [WIDTH*2-1+0:0] tmp00_73_32;
	wire [WIDTH*2-1+0:0] tmp00_73_33;
	wire [WIDTH*2-1+0:0] tmp00_73_34;
	wire [WIDTH*2-1+0:0] tmp00_73_35;
	wire [WIDTH*2-1+0:0] tmp00_73_36;
	wire [WIDTH*2-1+0:0] tmp00_73_37;
	wire [WIDTH*2-1+0:0] tmp00_73_38;
	wire [WIDTH*2-1+0:0] tmp00_73_39;
	wire [WIDTH*2-1+0:0] tmp00_73_40;
	wire [WIDTH*2-1+0:0] tmp00_73_41;
	wire [WIDTH*2-1+0:0] tmp00_73_42;
	wire [WIDTH*2-1+0:0] tmp00_73_43;
	wire [WIDTH*2-1+0:0] tmp00_73_44;
	wire [WIDTH*2-1+0:0] tmp00_73_45;
	wire [WIDTH*2-1+0:0] tmp00_73_46;
	wire [WIDTH*2-1+0:0] tmp00_73_47;
	wire [WIDTH*2-1+0:0] tmp00_73_48;
	wire [WIDTH*2-1+0:0] tmp00_73_49;
	wire [WIDTH*2-1+0:0] tmp00_73_50;
	wire [WIDTH*2-1+0:0] tmp00_73_51;
	wire [WIDTH*2-1+0:0] tmp00_73_52;
	wire [WIDTH*2-1+0:0] tmp00_73_53;
	wire [WIDTH*2-1+0:0] tmp00_73_54;
	wire [WIDTH*2-1+0:0] tmp00_73_55;
	wire [WIDTH*2-1+0:0] tmp00_73_56;
	wire [WIDTH*2-1+0:0] tmp00_73_57;
	wire [WIDTH*2-1+0:0] tmp00_73_58;
	wire [WIDTH*2-1+0:0] tmp00_73_59;
	wire [WIDTH*2-1+0:0] tmp00_73_60;
	wire [WIDTH*2-1+0:0] tmp00_73_61;
	wire [WIDTH*2-1+0:0] tmp00_73_62;
	wire [WIDTH*2-1+0:0] tmp00_73_63;
	wire [WIDTH*2-1+0:0] tmp00_73_64;
	wire [WIDTH*2-1+0:0] tmp00_73_65;
	wire [WIDTH*2-1+0:0] tmp00_73_66;
	wire [WIDTH*2-1+0:0] tmp00_73_67;
	wire [WIDTH*2-1+0:0] tmp00_73_68;
	wire [WIDTH*2-1+0:0] tmp00_73_69;
	wire [WIDTH*2-1+0:0] tmp00_73_70;
	wire [WIDTH*2-1+0:0] tmp00_73_71;
	wire [WIDTH*2-1+0:0] tmp00_73_72;
	wire [WIDTH*2-1+0:0] tmp00_73_73;
	wire [WIDTH*2-1+0:0] tmp00_73_74;
	wire [WIDTH*2-1+0:0] tmp00_73_75;
	wire [WIDTH*2-1+0:0] tmp00_73_76;
	wire [WIDTH*2-1+0:0] tmp00_73_77;
	wire [WIDTH*2-1+0:0] tmp00_73_78;
	wire [WIDTH*2-1+0:0] tmp00_73_79;
	wire [WIDTH*2-1+0:0] tmp00_73_80;
	wire [WIDTH*2-1+0:0] tmp00_73_81;
	wire [WIDTH*2-1+0:0] tmp00_73_82;
	wire [WIDTH*2-1+0:0] tmp00_73_83;
	wire [WIDTH*2-1+0:0] tmp00_74_0;
	wire [WIDTH*2-1+0:0] tmp00_74_1;
	wire [WIDTH*2-1+0:0] tmp00_74_2;
	wire [WIDTH*2-1+0:0] tmp00_74_3;
	wire [WIDTH*2-1+0:0] tmp00_74_4;
	wire [WIDTH*2-1+0:0] tmp00_74_5;
	wire [WIDTH*2-1+0:0] tmp00_74_6;
	wire [WIDTH*2-1+0:0] tmp00_74_7;
	wire [WIDTH*2-1+0:0] tmp00_74_8;
	wire [WIDTH*2-1+0:0] tmp00_74_9;
	wire [WIDTH*2-1+0:0] tmp00_74_10;
	wire [WIDTH*2-1+0:0] tmp00_74_11;
	wire [WIDTH*2-1+0:0] tmp00_74_12;
	wire [WIDTH*2-1+0:0] tmp00_74_13;
	wire [WIDTH*2-1+0:0] tmp00_74_14;
	wire [WIDTH*2-1+0:0] tmp00_74_15;
	wire [WIDTH*2-1+0:0] tmp00_74_16;
	wire [WIDTH*2-1+0:0] tmp00_74_17;
	wire [WIDTH*2-1+0:0] tmp00_74_18;
	wire [WIDTH*2-1+0:0] tmp00_74_19;
	wire [WIDTH*2-1+0:0] tmp00_74_20;
	wire [WIDTH*2-1+0:0] tmp00_74_21;
	wire [WIDTH*2-1+0:0] tmp00_74_22;
	wire [WIDTH*2-1+0:0] tmp00_74_23;
	wire [WIDTH*2-1+0:0] tmp00_74_24;
	wire [WIDTH*2-1+0:0] tmp00_74_25;
	wire [WIDTH*2-1+0:0] tmp00_74_26;
	wire [WIDTH*2-1+0:0] tmp00_74_27;
	wire [WIDTH*2-1+0:0] tmp00_74_28;
	wire [WIDTH*2-1+0:0] tmp00_74_29;
	wire [WIDTH*2-1+0:0] tmp00_74_30;
	wire [WIDTH*2-1+0:0] tmp00_74_31;
	wire [WIDTH*2-1+0:0] tmp00_74_32;
	wire [WIDTH*2-1+0:0] tmp00_74_33;
	wire [WIDTH*2-1+0:0] tmp00_74_34;
	wire [WIDTH*2-1+0:0] tmp00_74_35;
	wire [WIDTH*2-1+0:0] tmp00_74_36;
	wire [WIDTH*2-1+0:0] tmp00_74_37;
	wire [WIDTH*2-1+0:0] tmp00_74_38;
	wire [WIDTH*2-1+0:0] tmp00_74_39;
	wire [WIDTH*2-1+0:0] tmp00_74_40;
	wire [WIDTH*2-1+0:0] tmp00_74_41;
	wire [WIDTH*2-1+0:0] tmp00_74_42;
	wire [WIDTH*2-1+0:0] tmp00_74_43;
	wire [WIDTH*2-1+0:0] tmp00_74_44;
	wire [WIDTH*2-1+0:0] tmp00_74_45;
	wire [WIDTH*2-1+0:0] tmp00_74_46;
	wire [WIDTH*2-1+0:0] tmp00_74_47;
	wire [WIDTH*2-1+0:0] tmp00_74_48;
	wire [WIDTH*2-1+0:0] tmp00_74_49;
	wire [WIDTH*2-1+0:0] tmp00_74_50;
	wire [WIDTH*2-1+0:0] tmp00_74_51;
	wire [WIDTH*2-1+0:0] tmp00_74_52;
	wire [WIDTH*2-1+0:0] tmp00_74_53;
	wire [WIDTH*2-1+0:0] tmp00_74_54;
	wire [WIDTH*2-1+0:0] tmp00_74_55;
	wire [WIDTH*2-1+0:0] tmp00_74_56;
	wire [WIDTH*2-1+0:0] tmp00_74_57;
	wire [WIDTH*2-1+0:0] tmp00_74_58;
	wire [WIDTH*2-1+0:0] tmp00_74_59;
	wire [WIDTH*2-1+0:0] tmp00_74_60;
	wire [WIDTH*2-1+0:0] tmp00_74_61;
	wire [WIDTH*2-1+0:0] tmp00_74_62;
	wire [WIDTH*2-1+0:0] tmp00_74_63;
	wire [WIDTH*2-1+0:0] tmp00_74_64;
	wire [WIDTH*2-1+0:0] tmp00_74_65;
	wire [WIDTH*2-1+0:0] tmp00_74_66;
	wire [WIDTH*2-1+0:0] tmp00_74_67;
	wire [WIDTH*2-1+0:0] tmp00_74_68;
	wire [WIDTH*2-1+0:0] tmp00_74_69;
	wire [WIDTH*2-1+0:0] tmp00_74_70;
	wire [WIDTH*2-1+0:0] tmp00_74_71;
	wire [WIDTH*2-1+0:0] tmp00_74_72;
	wire [WIDTH*2-1+0:0] tmp00_74_73;
	wire [WIDTH*2-1+0:0] tmp00_74_74;
	wire [WIDTH*2-1+0:0] tmp00_74_75;
	wire [WIDTH*2-1+0:0] tmp00_74_76;
	wire [WIDTH*2-1+0:0] tmp00_74_77;
	wire [WIDTH*2-1+0:0] tmp00_74_78;
	wire [WIDTH*2-1+0:0] tmp00_74_79;
	wire [WIDTH*2-1+0:0] tmp00_74_80;
	wire [WIDTH*2-1+0:0] tmp00_74_81;
	wire [WIDTH*2-1+0:0] tmp00_74_82;
	wire [WIDTH*2-1+0:0] tmp00_74_83;
	wire [WIDTH*2-1+0:0] tmp00_75_0;
	wire [WIDTH*2-1+0:0] tmp00_75_1;
	wire [WIDTH*2-1+0:0] tmp00_75_2;
	wire [WIDTH*2-1+0:0] tmp00_75_3;
	wire [WIDTH*2-1+0:0] tmp00_75_4;
	wire [WIDTH*2-1+0:0] tmp00_75_5;
	wire [WIDTH*2-1+0:0] tmp00_75_6;
	wire [WIDTH*2-1+0:0] tmp00_75_7;
	wire [WIDTH*2-1+0:0] tmp00_75_8;
	wire [WIDTH*2-1+0:0] tmp00_75_9;
	wire [WIDTH*2-1+0:0] tmp00_75_10;
	wire [WIDTH*2-1+0:0] tmp00_75_11;
	wire [WIDTH*2-1+0:0] tmp00_75_12;
	wire [WIDTH*2-1+0:0] tmp00_75_13;
	wire [WIDTH*2-1+0:0] tmp00_75_14;
	wire [WIDTH*2-1+0:0] tmp00_75_15;
	wire [WIDTH*2-1+0:0] tmp00_75_16;
	wire [WIDTH*2-1+0:0] tmp00_75_17;
	wire [WIDTH*2-1+0:0] tmp00_75_18;
	wire [WIDTH*2-1+0:0] tmp00_75_19;
	wire [WIDTH*2-1+0:0] tmp00_75_20;
	wire [WIDTH*2-1+0:0] tmp00_75_21;
	wire [WIDTH*2-1+0:0] tmp00_75_22;
	wire [WIDTH*2-1+0:0] tmp00_75_23;
	wire [WIDTH*2-1+0:0] tmp00_75_24;
	wire [WIDTH*2-1+0:0] tmp00_75_25;
	wire [WIDTH*2-1+0:0] tmp00_75_26;
	wire [WIDTH*2-1+0:0] tmp00_75_27;
	wire [WIDTH*2-1+0:0] tmp00_75_28;
	wire [WIDTH*2-1+0:0] tmp00_75_29;
	wire [WIDTH*2-1+0:0] tmp00_75_30;
	wire [WIDTH*2-1+0:0] tmp00_75_31;
	wire [WIDTH*2-1+0:0] tmp00_75_32;
	wire [WIDTH*2-1+0:0] tmp00_75_33;
	wire [WIDTH*2-1+0:0] tmp00_75_34;
	wire [WIDTH*2-1+0:0] tmp00_75_35;
	wire [WIDTH*2-1+0:0] tmp00_75_36;
	wire [WIDTH*2-1+0:0] tmp00_75_37;
	wire [WIDTH*2-1+0:0] tmp00_75_38;
	wire [WIDTH*2-1+0:0] tmp00_75_39;
	wire [WIDTH*2-1+0:0] tmp00_75_40;
	wire [WIDTH*2-1+0:0] tmp00_75_41;
	wire [WIDTH*2-1+0:0] tmp00_75_42;
	wire [WIDTH*2-1+0:0] tmp00_75_43;
	wire [WIDTH*2-1+0:0] tmp00_75_44;
	wire [WIDTH*2-1+0:0] tmp00_75_45;
	wire [WIDTH*2-1+0:0] tmp00_75_46;
	wire [WIDTH*2-1+0:0] tmp00_75_47;
	wire [WIDTH*2-1+0:0] tmp00_75_48;
	wire [WIDTH*2-1+0:0] tmp00_75_49;
	wire [WIDTH*2-1+0:0] tmp00_75_50;
	wire [WIDTH*2-1+0:0] tmp00_75_51;
	wire [WIDTH*2-1+0:0] tmp00_75_52;
	wire [WIDTH*2-1+0:0] tmp00_75_53;
	wire [WIDTH*2-1+0:0] tmp00_75_54;
	wire [WIDTH*2-1+0:0] tmp00_75_55;
	wire [WIDTH*2-1+0:0] tmp00_75_56;
	wire [WIDTH*2-1+0:0] tmp00_75_57;
	wire [WIDTH*2-1+0:0] tmp00_75_58;
	wire [WIDTH*2-1+0:0] tmp00_75_59;
	wire [WIDTH*2-1+0:0] tmp00_75_60;
	wire [WIDTH*2-1+0:0] tmp00_75_61;
	wire [WIDTH*2-1+0:0] tmp00_75_62;
	wire [WIDTH*2-1+0:0] tmp00_75_63;
	wire [WIDTH*2-1+0:0] tmp00_75_64;
	wire [WIDTH*2-1+0:0] tmp00_75_65;
	wire [WIDTH*2-1+0:0] tmp00_75_66;
	wire [WIDTH*2-1+0:0] tmp00_75_67;
	wire [WIDTH*2-1+0:0] tmp00_75_68;
	wire [WIDTH*2-1+0:0] tmp00_75_69;
	wire [WIDTH*2-1+0:0] tmp00_75_70;
	wire [WIDTH*2-1+0:0] tmp00_75_71;
	wire [WIDTH*2-1+0:0] tmp00_75_72;
	wire [WIDTH*2-1+0:0] tmp00_75_73;
	wire [WIDTH*2-1+0:0] tmp00_75_74;
	wire [WIDTH*2-1+0:0] tmp00_75_75;
	wire [WIDTH*2-1+0:0] tmp00_75_76;
	wire [WIDTH*2-1+0:0] tmp00_75_77;
	wire [WIDTH*2-1+0:0] tmp00_75_78;
	wire [WIDTH*2-1+0:0] tmp00_75_79;
	wire [WIDTH*2-1+0:0] tmp00_75_80;
	wire [WIDTH*2-1+0:0] tmp00_75_81;
	wire [WIDTH*2-1+0:0] tmp00_75_82;
	wire [WIDTH*2-1+0:0] tmp00_75_83;
	wire [WIDTH*2-1+0:0] tmp00_76_0;
	wire [WIDTH*2-1+0:0] tmp00_76_1;
	wire [WIDTH*2-1+0:0] tmp00_76_2;
	wire [WIDTH*2-1+0:0] tmp00_76_3;
	wire [WIDTH*2-1+0:0] tmp00_76_4;
	wire [WIDTH*2-1+0:0] tmp00_76_5;
	wire [WIDTH*2-1+0:0] tmp00_76_6;
	wire [WIDTH*2-1+0:0] tmp00_76_7;
	wire [WIDTH*2-1+0:0] tmp00_76_8;
	wire [WIDTH*2-1+0:0] tmp00_76_9;
	wire [WIDTH*2-1+0:0] tmp00_76_10;
	wire [WIDTH*2-1+0:0] tmp00_76_11;
	wire [WIDTH*2-1+0:0] tmp00_76_12;
	wire [WIDTH*2-1+0:0] tmp00_76_13;
	wire [WIDTH*2-1+0:0] tmp00_76_14;
	wire [WIDTH*2-1+0:0] tmp00_76_15;
	wire [WIDTH*2-1+0:0] tmp00_76_16;
	wire [WIDTH*2-1+0:0] tmp00_76_17;
	wire [WIDTH*2-1+0:0] tmp00_76_18;
	wire [WIDTH*2-1+0:0] tmp00_76_19;
	wire [WIDTH*2-1+0:0] tmp00_76_20;
	wire [WIDTH*2-1+0:0] tmp00_76_21;
	wire [WIDTH*2-1+0:0] tmp00_76_22;
	wire [WIDTH*2-1+0:0] tmp00_76_23;
	wire [WIDTH*2-1+0:0] tmp00_76_24;
	wire [WIDTH*2-1+0:0] tmp00_76_25;
	wire [WIDTH*2-1+0:0] tmp00_76_26;
	wire [WIDTH*2-1+0:0] tmp00_76_27;
	wire [WIDTH*2-1+0:0] tmp00_76_28;
	wire [WIDTH*2-1+0:0] tmp00_76_29;
	wire [WIDTH*2-1+0:0] tmp00_76_30;
	wire [WIDTH*2-1+0:0] tmp00_76_31;
	wire [WIDTH*2-1+0:0] tmp00_76_32;
	wire [WIDTH*2-1+0:0] tmp00_76_33;
	wire [WIDTH*2-1+0:0] tmp00_76_34;
	wire [WIDTH*2-1+0:0] tmp00_76_35;
	wire [WIDTH*2-1+0:0] tmp00_76_36;
	wire [WIDTH*2-1+0:0] tmp00_76_37;
	wire [WIDTH*2-1+0:0] tmp00_76_38;
	wire [WIDTH*2-1+0:0] tmp00_76_39;
	wire [WIDTH*2-1+0:0] tmp00_76_40;
	wire [WIDTH*2-1+0:0] tmp00_76_41;
	wire [WIDTH*2-1+0:0] tmp00_76_42;
	wire [WIDTH*2-1+0:0] tmp00_76_43;
	wire [WIDTH*2-1+0:0] tmp00_76_44;
	wire [WIDTH*2-1+0:0] tmp00_76_45;
	wire [WIDTH*2-1+0:0] tmp00_76_46;
	wire [WIDTH*2-1+0:0] tmp00_76_47;
	wire [WIDTH*2-1+0:0] tmp00_76_48;
	wire [WIDTH*2-1+0:0] tmp00_76_49;
	wire [WIDTH*2-1+0:0] tmp00_76_50;
	wire [WIDTH*2-1+0:0] tmp00_76_51;
	wire [WIDTH*2-1+0:0] tmp00_76_52;
	wire [WIDTH*2-1+0:0] tmp00_76_53;
	wire [WIDTH*2-1+0:0] tmp00_76_54;
	wire [WIDTH*2-1+0:0] tmp00_76_55;
	wire [WIDTH*2-1+0:0] tmp00_76_56;
	wire [WIDTH*2-1+0:0] tmp00_76_57;
	wire [WIDTH*2-1+0:0] tmp00_76_58;
	wire [WIDTH*2-1+0:0] tmp00_76_59;
	wire [WIDTH*2-1+0:0] tmp00_76_60;
	wire [WIDTH*2-1+0:0] tmp00_76_61;
	wire [WIDTH*2-1+0:0] tmp00_76_62;
	wire [WIDTH*2-1+0:0] tmp00_76_63;
	wire [WIDTH*2-1+0:0] tmp00_76_64;
	wire [WIDTH*2-1+0:0] tmp00_76_65;
	wire [WIDTH*2-1+0:0] tmp00_76_66;
	wire [WIDTH*2-1+0:0] tmp00_76_67;
	wire [WIDTH*2-1+0:0] tmp00_76_68;
	wire [WIDTH*2-1+0:0] tmp00_76_69;
	wire [WIDTH*2-1+0:0] tmp00_76_70;
	wire [WIDTH*2-1+0:0] tmp00_76_71;
	wire [WIDTH*2-1+0:0] tmp00_76_72;
	wire [WIDTH*2-1+0:0] tmp00_76_73;
	wire [WIDTH*2-1+0:0] tmp00_76_74;
	wire [WIDTH*2-1+0:0] tmp00_76_75;
	wire [WIDTH*2-1+0:0] tmp00_76_76;
	wire [WIDTH*2-1+0:0] tmp00_76_77;
	wire [WIDTH*2-1+0:0] tmp00_76_78;
	wire [WIDTH*2-1+0:0] tmp00_76_79;
	wire [WIDTH*2-1+0:0] tmp00_76_80;
	wire [WIDTH*2-1+0:0] tmp00_76_81;
	wire [WIDTH*2-1+0:0] tmp00_76_82;
	wire [WIDTH*2-1+0:0] tmp00_76_83;
	wire [WIDTH*2-1+0:0] tmp00_77_0;
	wire [WIDTH*2-1+0:0] tmp00_77_1;
	wire [WIDTH*2-1+0:0] tmp00_77_2;
	wire [WIDTH*2-1+0:0] tmp00_77_3;
	wire [WIDTH*2-1+0:0] tmp00_77_4;
	wire [WIDTH*2-1+0:0] tmp00_77_5;
	wire [WIDTH*2-1+0:0] tmp00_77_6;
	wire [WIDTH*2-1+0:0] tmp00_77_7;
	wire [WIDTH*2-1+0:0] tmp00_77_8;
	wire [WIDTH*2-1+0:0] tmp00_77_9;
	wire [WIDTH*2-1+0:0] tmp00_77_10;
	wire [WIDTH*2-1+0:0] tmp00_77_11;
	wire [WIDTH*2-1+0:0] tmp00_77_12;
	wire [WIDTH*2-1+0:0] tmp00_77_13;
	wire [WIDTH*2-1+0:0] tmp00_77_14;
	wire [WIDTH*2-1+0:0] tmp00_77_15;
	wire [WIDTH*2-1+0:0] tmp00_77_16;
	wire [WIDTH*2-1+0:0] tmp00_77_17;
	wire [WIDTH*2-1+0:0] tmp00_77_18;
	wire [WIDTH*2-1+0:0] tmp00_77_19;
	wire [WIDTH*2-1+0:0] tmp00_77_20;
	wire [WIDTH*2-1+0:0] tmp00_77_21;
	wire [WIDTH*2-1+0:0] tmp00_77_22;
	wire [WIDTH*2-1+0:0] tmp00_77_23;
	wire [WIDTH*2-1+0:0] tmp00_77_24;
	wire [WIDTH*2-1+0:0] tmp00_77_25;
	wire [WIDTH*2-1+0:0] tmp00_77_26;
	wire [WIDTH*2-1+0:0] tmp00_77_27;
	wire [WIDTH*2-1+0:0] tmp00_77_28;
	wire [WIDTH*2-1+0:0] tmp00_77_29;
	wire [WIDTH*2-1+0:0] tmp00_77_30;
	wire [WIDTH*2-1+0:0] tmp00_77_31;
	wire [WIDTH*2-1+0:0] tmp00_77_32;
	wire [WIDTH*2-1+0:0] tmp00_77_33;
	wire [WIDTH*2-1+0:0] tmp00_77_34;
	wire [WIDTH*2-1+0:0] tmp00_77_35;
	wire [WIDTH*2-1+0:0] tmp00_77_36;
	wire [WIDTH*2-1+0:0] tmp00_77_37;
	wire [WIDTH*2-1+0:0] tmp00_77_38;
	wire [WIDTH*2-1+0:0] tmp00_77_39;
	wire [WIDTH*2-1+0:0] tmp00_77_40;
	wire [WIDTH*2-1+0:0] tmp00_77_41;
	wire [WIDTH*2-1+0:0] tmp00_77_42;
	wire [WIDTH*2-1+0:0] tmp00_77_43;
	wire [WIDTH*2-1+0:0] tmp00_77_44;
	wire [WIDTH*2-1+0:0] tmp00_77_45;
	wire [WIDTH*2-1+0:0] tmp00_77_46;
	wire [WIDTH*2-1+0:0] tmp00_77_47;
	wire [WIDTH*2-1+0:0] tmp00_77_48;
	wire [WIDTH*2-1+0:0] tmp00_77_49;
	wire [WIDTH*2-1+0:0] tmp00_77_50;
	wire [WIDTH*2-1+0:0] tmp00_77_51;
	wire [WIDTH*2-1+0:0] tmp00_77_52;
	wire [WIDTH*2-1+0:0] tmp00_77_53;
	wire [WIDTH*2-1+0:0] tmp00_77_54;
	wire [WIDTH*2-1+0:0] tmp00_77_55;
	wire [WIDTH*2-1+0:0] tmp00_77_56;
	wire [WIDTH*2-1+0:0] tmp00_77_57;
	wire [WIDTH*2-1+0:0] tmp00_77_58;
	wire [WIDTH*2-1+0:0] tmp00_77_59;
	wire [WIDTH*2-1+0:0] tmp00_77_60;
	wire [WIDTH*2-1+0:0] tmp00_77_61;
	wire [WIDTH*2-1+0:0] tmp00_77_62;
	wire [WIDTH*2-1+0:0] tmp00_77_63;
	wire [WIDTH*2-1+0:0] tmp00_77_64;
	wire [WIDTH*2-1+0:0] tmp00_77_65;
	wire [WIDTH*2-1+0:0] tmp00_77_66;
	wire [WIDTH*2-1+0:0] tmp00_77_67;
	wire [WIDTH*2-1+0:0] tmp00_77_68;
	wire [WIDTH*2-1+0:0] tmp00_77_69;
	wire [WIDTH*2-1+0:0] tmp00_77_70;
	wire [WIDTH*2-1+0:0] tmp00_77_71;
	wire [WIDTH*2-1+0:0] tmp00_77_72;
	wire [WIDTH*2-1+0:0] tmp00_77_73;
	wire [WIDTH*2-1+0:0] tmp00_77_74;
	wire [WIDTH*2-1+0:0] tmp00_77_75;
	wire [WIDTH*2-1+0:0] tmp00_77_76;
	wire [WIDTH*2-1+0:0] tmp00_77_77;
	wire [WIDTH*2-1+0:0] tmp00_77_78;
	wire [WIDTH*2-1+0:0] tmp00_77_79;
	wire [WIDTH*2-1+0:0] tmp00_77_80;
	wire [WIDTH*2-1+0:0] tmp00_77_81;
	wire [WIDTH*2-1+0:0] tmp00_77_82;
	wire [WIDTH*2-1+0:0] tmp00_77_83;
	wire [WIDTH*2-1+0:0] tmp00_78_0;
	wire [WIDTH*2-1+0:0] tmp00_78_1;
	wire [WIDTH*2-1+0:0] tmp00_78_2;
	wire [WIDTH*2-1+0:0] tmp00_78_3;
	wire [WIDTH*2-1+0:0] tmp00_78_4;
	wire [WIDTH*2-1+0:0] tmp00_78_5;
	wire [WIDTH*2-1+0:0] tmp00_78_6;
	wire [WIDTH*2-1+0:0] tmp00_78_7;
	wire [WIDTH*2-1+0:0] tmp00_78_8;
	wire [WIDTH*2-1+0:0] tmp00_78_9;
	wire [WIDTH*2-1+0:0] tmp00_78_10;
	wire [WIDTH*2-1+0:0] tmp00_78_11;
	wire [WIDTH*2-1+0:0] tmp00_78_12;
	wire [WIDTH*2-1+0:0] tmp00_78_13;
	wire [WIDTH*2-1+0:0] tmp00_78_14;
	wire [WIDTH*2-1+0:0] tmp00_78_15;
	wire [WIDTH*2-1+0:0] tmp00_78_16;
	wire [WIDTH*2-1+0:0] tmp00_78_17;
	wire [WIDTH*2-1+0:0] tmp00_78_18;
	wire [WIDTH*2-1+0:0] tmp00_78_19;
	wire [WIDTH*2-1+0:0] tmp00_78_20;
	wire [WIDTH*2-1+0:0] tmp00_78_21;
	wire [WIDTH*2-1+0:0] tmp00_78_22;
	wire [WIDTH*2-1+0:0] tmp00_78_23;
	wire [WIDTH*2-1+0:0] tmp00_78_24;
	wire [WIDTH*2-1+0:0] tmp00_78_25;
	wire [WIDTH*2-1+0:0] tmp00_78_26;
	wire [WIDTH*2-1+0:0] tmp00_78_27;
	wire [WIDTH*2-1+0:0] tmp00_78_28;
	wire [WIDTH*2-1+0:0] tmp00_78_29;
	wire [WIDTH*2-1+0:0] tmp00_78_30;
	wire [WIDTH*2-1+0:0] tmp00_78_31;
	wire [WIDTH*2-1+0:0] tmp00_78_32;
	wire [WIDTH*2-1+0:0] tmp00_78_33;
	wire [WIDTH*2-1+0:0] tmp00_78_34;
	wire [WIDTH*2-1+0:0] tmp00_78_35;
	wire [WIDTH*2-1+0:0] tmp00_78_36;
	wire [WIDTH*2-1+0:0] tmp00_78_37;
	wire [WIDTH*2-1+0:0] tmp00_78_38;
	wire [WIDTH*2-1+0:0] tmp00_78_39;
	wire [WIDTH*2-1+0:0] tmp00_78_40;
	wire [WIDTH*2-1+0:0] tmp00_78_41;
	wire [WIDTH*2-1+0:0] tmp00_78_42;
	wire [WIDTH*2-1+0:0] tmp00_78_43;
	wire [WIDTH*2-1+0:0] tmp00_78_44;
	wire [WIDTH*2-1+0:0] tmp00_78_45;
	wire [WIDTH*2-1+0:0] tmp00_78_46;
	wire [WIDTH*2-1+0:0] tmp00_78_47;
	wire [WIDTH*2-1+0:0] tmp00_78_48;
	wire [WIDTH*2-1+0:0] tmp00_78_49;
	wire [WIDTH*2-1+0:0] tmp00_78_50;
	wire [WIDTH*2-1+0:0] tmp00_78_51;
	wire [WIDTH*2-1+0:0] tmp00_78_52;
	wire [WIDTH*2-1+0:0] tmp00_78_53;
	wire [WIDTH*2-1+0:0] tmp00_78_54;
	wire [WIDTH*2-1+0:0] tmp00_78_55;
	wire [WIDTH*2-1+0:0] tmp00_78_56;
	wire [WIDTH*2-1+0:0] tmp00_78_57;
	wire [WIDTH*2-1+0:0] tmp00_78_58;
	wire [WIDTH*2-1+0:0] tmp00_78_59;
	wire [WIDTH*2-1+0:0] tmp00_78_60;
	wire [WIDTH*2-1+0:0] tmp00_78_61;
	wire [WIDTH*2-1+0:0] tmp00_78_62;
	wire [WIDTH*2-1+0:0] tmp00_78_63;
	wire [WIDTH*2-1+0:0] tmp00_78_64;
	wire [WIDTH*2-1+0:0] tmp00_78_65;
	wire [WIDTH*2-1+0:0] tmp00_78_66;
	wire [WIDTH*2-1+0:0] tmp00_78_67;
	wire [WIDTH*2-1+0:0] tmp00_78_68;
	wire [WIDTH*2-1+0:0] tmp00_78_69;
	wire [WIDTH*2-1+0:0] tmp00_78_70;
	wire [WIDTH*2-1+0:0] tmp00_78_71;
	wire [WIDTH*2-1+0:0] tmp00_78_72;
	wire [WIDTH*2-1+0:0] tmp00_78_73;
	wire [WIDTH*2-1+0:0] tmp00_78_74;
	wire [WIDTH*2-1+0:0] tmp00_78_75;
	wire [WIDTH*2-1+0:0] tmp00_78_76;
	wire [WIDTH*2-1+0:0] tmp00_78_77;
	wire [WIDTH*2-1+0:0] tmp00_78_78;
	wire [WIDTH*2-1+0:0] tmp00_78_79;
	wire [WIDTH*2-1+0:0] tmp00_78_80;
	wire [WIDTH*2-1+0:0] tmp00_78_81;
	wire [WIDTH*2-1+0:0] tmp00_78_82;
	wire [WIDTH*2-1+0:0] tmp00_78_83;
	wire [WIDTH*2-1+0:0] tmp00_79_0;
	wire [WIDTH*2-1+0:0] tmp00_79_1;
	wire [WIDTH*2-1+0:0] tmp00_79_2;
	wire [WIDTH*2-1+0:0] tmp00_79_3;
	wire [WIDTH*2-1+0:0] tmp00_79_4;
	wire [WIDTH*2-1+0:0] tmp00_79_5;
	wire [WIDTH*2-1+0:0] tmp00_79_6;
	wire [WIDTH*2-1+0:0] tmp00_79_7;
	wire [WIDTH*2-1+0:0] tmp00_79_8;
	wire [WIDTH*2-1+0:0] tmp00_79_9;
	wire [WIDTH*2-1+0:0] tmp00_79_10;
	wire [WIDTH*2-1+0:0] tmp00_79_11;
	wire [WIDTH*2-1+0:0] tmp00_79_12;
	wire [WIDTH*2-1+0:0] tmp00_79_13;
	wire [WIDTH*2-1+0:0] tmp00_79_14;
	wire [WIDTH*2-1+0:0] tmp00_79_15;
	wire [WIDTH*2-1+0:0] tmp00_79_16;
	wire [WIDTH*2-1+0:0] tmp00_79_17;
	wire [WIDTH*2-1+0:0] tmp00_79_18;
	wire [WIDTH*2-1+0:0] tmp00_79_19;
	wire [WIDTH*2-1+0:0] tmp00_79_20;
	wire [WIDTH*2-1+0:0] tmp00_79_21;
	wire [WIDTH*2-1+0:0] tmp00_79_22;
	wire [WIDTH*2-1+0:0] tmp00_79_23;
	wire [WIDTH*2-1+0:0] tmp00_79_24;
	wire [WIDTH*2-1+0:0] tmp00_79_25;
	wire [WIDTH*2-1+0:0] tmp00_79_26;
	wire [WIDTH*2-1+0:0] tmp00_79_27;
	wire [WIDTH*2-1+0:0] tmp00_79_28;
	wire [WIDTH*2-1+0:0] tmp00_79_29;
	wire [WIDTH*2-1+0:0] tmp00_79_30;
	wire [WIDTH*2-1+0:0] tmp00_79_31;
	wire [WIDTH*2-1+0:0] tmp00_79_32;
	wire [WIDTH*2-1+0:0] tmp00_79_33;
	wire [WIDTH*2-1+0:0] tmp00_79_34;
	wire [WIDTH*2-1+0:0] tmp00_79_35;
	wire [WIDTH*2-1+0:0] tmp00_79_36;
	wire [WIDTH*2-1+0:0] tmp00_79_37;
	wire [WIDTH*2-1+0:0] tmp00_79_38;
	wire [WIDTH*2-1+0:0] tmp00_79_39;
	wire [WIDTH*2-1+0:0] tmp00_79_40;
	wire [WIDTH*2-1+0:0] tmp00_79_41;
	wire [WIDTH*2-1+0:0] tmp00_79_42;
	wire [WIDTH*2-1+0:0] tmp00_79_43;
	wire [WIDTH*2-1+0:0] tmp00_79_44;
	wire [WIDTH*2-1+0:0] tmp00_79_45;
	wire [WIDTH*2-1+0:0] tmp00_79_46;
	wire [WIDTH*2-1+0:0] tmp00_79_47;
	wire [WIDTH*2-1+0:0] tmp00_79_48;
	wire [WIDTH*2-1+0:0] tmp00_79_49;
	wire [WIDTH*2-1+0:0] tmp00_79_50;
	wire [WIDTH*2-1+0:0] tmp00_79_51;
	wire [WIDTH*2-1+0:0] tmp00_79_52;
	wire [WIDTH*2-1+0:0] tmp00_79_53;
	wire [WIDTH*2-1+0:0] tmp00_79_54;
	wire [WIDTH*2-1+0:0] tmp00_79_55;
	wire [WIDTH*2-1+0:0] tmp00_79_56;
	wire [WIDTH*2-1+0:0] tmp00_79_57;
	wire [WIDTH*2-1+0:0] tmp00_79_58;
	wire [WIDTH*2-1+0:0] tmp00_79_59;
	wire [WIDTH*2-1+0:0] tmp00_79_60;
	wire [WIDTH*2-1+0:0] tmp00_79_61;
	wire [WIDTH*2-1+0:0] tmp00_79_62;
	wire [WIDTH*2-1+0:0] tmp00_79_63;
	wire [WIDTH*2-1+0:0] tmp00_79_64;
	wire [WIDTH*2-1+0:0] tmp00_79_65;
	wire [WIDTH*2-1+0:0] tmp00_79_66;
	wire [WIDTH*2-1+0:0] tmp00_79_67;
	wire [WIDTH*2-1+0:0] tmp00_79_68;
	wire [WIDTH*2-1+0:0] tmp00_79_69;
	wire [WIDTH*2-1+0:0] tmp00_79_70;
	wire [WIDTH*2-1+0:0] tmp00_79_71;
	wire [WIDTH*2-1+0:0] tmp00_79_72;
	wire [WIDTH*2-1+0:0] tmp00_79_73;
	wire [WIDTH*2-1+0:0] tmp00_79_74;
	wire [WIDTH*2-1+0:0] tmp00_79_75;
	wire [WIDTH*2-1+0:0] tmp00_79_76;
	wire [WIDTH*2-1+0:0] tmp00_79_77;
	wire [WIDTH*2-1+0:0] tmp00_79_78;
	wire [WIDTH*2-1+0:0] tmp00_79_79;
	wire [WIDTH*2-1+0:0] tmp00_79_80;
	wire [WIDTH*2-1+0:0] tmp00_79_81;
	wire [WIDTH*2-1+0:0] tmp00_79_82;
	wire [WIDTH*2-1+0:0] tmp00_79_83;
	wire [WIDTH*2-1+0:0] tmp00_80_0;
	wire [WIDTH*2-1+0:0] tmp00_80_1;
	wire [WIDTH*2-1+0:0] tmp00_80_2;
	wire [WIDTH*2-1+0:0] tmp00_80_3;
	wire [WIDTH*2-1+0:0] tmp00_80_4;
	wire [WIDTH*2-1+0:0] tmp00_80_5;
	wire [WIDTH*2-1+0:0] tmp00_80_6;
	wire [WIDTH*2-1+0:0] tmp00_80_7;
	wire [WIDTH*2-1+0:0] tmp00_80_8;
	wire [WIDTH*2-1+0:0] tmp00_80_9;
	wire [WIDTH*2-1+0:0] tmp00_80_10;
	wire [WIDTH*2-1+0:0] tmp00_80_11;
	wire [WIDTH*2-1+0:0] tmp00_80_12;
	wire [WIDTH*2-1+0:0] tmp00_80_13;
	wire [WIDTH*2-1+0:0] tmp00_80_14;
	wire [WIDTH*2-1+0:0] tmp00_80_15;
	wire [WIDTH*2-1+0:0] tmp00_80_16;
	wire [WIDTH*2-1+0:0] tmp00_80_17;
	wire [WIDTH*2-1+0:0] tmp00_80_18;
	wire [WIDTH*2-1+0:0] tmp00_80_19;
	wire [WIDTH*2-1+0:0] tmp00_80_20;
	wire [WIDTH*2-1+0:0] tmp00_80_21;
	wire [WIDTH*2-1+0:0] tmp00_80_22;
	wire [WIDTH*2-1+0:0] tmp00_80_23;
	wire [WIDTH*2-1+0:0] tmp00_80_24;
	wire [WIDTH*2-1+0:0] tmp00_80_25;
	wire [WIDTH*2-1+0:0] tmp00_80_26;
	wire [WIDTH*2-1+0:0] tmp00_80_27;
	wire [WIDTH*2-1+0:0] tmp00_80_28;
	wire [WIDTH*2-1+0:0] tmp00_80_29;
	wire [WIDTH*2-1+0:0] tmp00_80_30;
	wire [WIDTH*2-1+0:0] tmp00_80_31;
	wire [WIDTH*2-1+0:0] tmp00_80_32;
	wire [WIDTH*2-1+0:0] tmp00_80_33;
	wire [WIDTH*2-1+0:0] tmp00_80_34;
	wire [WIDTH*2-1+0:0] tmp00_80_35;
	wire [WIDTH*2-1+0:0] tmp00_80_36;
	wire [WIDTH*2-1+0:0] tmp00_80_37;
	wire [WIDTH*2-1+0:0] tmp00_80_38;
	wire [WIDTH*2-1+0:0] tmp00_80_39;
	wire [WIDTH*2-1+0:0] tmp00_80_40;
	wire [WIDTH*2-1+0:0] tmp00_80_41;
	wire [WIDTH*2-1+0:0] tmp00_80_42;
	wire [WIDTH*2-1+0:0] tmp00_80_43;
	wire [WIDTH*2-1+0:0] tmp00_80_44;
	wire [WIDTH*2-1+0:0] tmp00_80_45;
	wire [WIDTH*2-1+0:0] tmp00_80_46;
	wire [WIDTH*2-1+0:0] tmp00_80_47;
	wire [WIDTH*2-1+0:0] tmp00_80_48;
	wire [WIDTH*2-1+0:0] tmp00_80_49;
	wire [WIDTH*2-1+0:0] tmp00_80_50;
	wire [WIDTH*2-1+0:0] tmp00_80_51;
	wire [WIDTH*2-1+0:0] tmp00_80_52;
	wire [WIDTH*2-1+0:0] tmp00_80_53;
	wire [WIDTH*2-1+0:0] tmp00_80_54;
	wire [WIDTH*2-1+0:0] tmp00_80_55;
	wire [WIDTH*2-1+0:0] tmp00_80_56;
	wire [WIDTH*2-1+0:0] tmp00_80_57;
	wire [WIDTH*2-1+0:0] tmp00_80_58;
	wire [WIDTH*2-1+0:0] tmp00_80_59;
	wire [WIDTH*2-1+0:0] tmp00_80_60;
	wire [WIDTH*2-1+0:0] tmp00_80_61;
	wire [WIDTH*2-1+0:0] tmp00_80_62;
	wire [WIDTH*2-1+0:0] tmp00_80_63;
	wire [WIDTH*2-1+0:0] tmp00_80_64;
	wire [WIDTH*2-1+0:0] tmp00_80_65;
	wire [WIDTH*2-1+0:0] tmp00_80_66;
	wire [WIDTH*2-1+0:0] tmp00_80_67;
	wire [WIDTH*2-1+0:0] tmp00_80_68;
	wire [WIDTH*2-1+0:0] tmp00_80_69;
	wire [WIDTH*2-1+0:0] tmp00_80_70;
	wire [WIDTH*2-1+0:0] tmp00_80_71;
	wire [WIDTH*2-1+0:0] tmp00_80_72;
	wire [WIDTH*2-1+0:0] tmp00_80_73;
	wire [WIDTH*2-1+0:0] tmp00_80_74;
	wire [WIDTH*2-1+0:0] tmp00_80_75;
	wire [WIDTH*2-1+0:0] tmp00_80_76;
	wire [WIDTH*2-1+0:0] tmp00_80_77;
	wire [WIDTH*2-1+0:0] tmp00_80_78;
	wire [WIDTH*2-1+0:0] tmp00_80_79;
	wire [WIDTH*2-1+0:0] tmp00_80_80;
	wire [WIDTH*2-1+0:0] tmp00_80_81;
	wire [WIDTH*2-1+0:0] tmp00_80_82;
	wire [WIDTH*2-1+0:0] tmp00_80_83;
	wire [WIDTH*2-1+0:0] tmp00_81_0;
	wire [WIDTH*2-1+0:0] tmp00_81_1;
	wire [WIDTH*2-1+0:0] tmp00_81_2;
	wire [WIDTH*2-1+0:0] tmp00_81_3;
	wire [WIDTH*2-1+0:0] tmp00_81_4;
	wire [WIDTH*2-1+0:0] tmp00_81_5;
	wire [WIDTH*2-1+0:0] tmp00_81_6;
	wire [WIDTH*2-1+0:0] tmp00_81_7;
	wire [WIDTH*2-1+0:0] tmp00_81_8;
	wire [WIDTH*2-1+0:0] tmp00_81_9;
	wire [WIDTH*2-1+0:0] tmp00_81_10;
	wire [WIDTH*2-1+0:0] tmp00_81_11;
	wire [WIDTH*2-1+0:0] tmp00_81_12;
	wire [WIDTH*2-1+0:0] tmp00_81_13;
	wire [WIDTH*2-1+0:0] tmp00_81_14;
	wire [WIDTH*2-1+0:0] tmp00_81_15;
	wire [WIDTH*2-1+0:0] tmp00_81_16;
	wire [WIDTH*2-1+0:0] tmp00_81_17;
	wire [WIDTH*2-1+0:0] tmp00_81_18;
	wire [WIDTH*2-1+0:0] tmp00_81_19;
	wire [WIDTH*2-1+0:0] tmp00_81_20;
	wire [WIDTH*2-1+0:0] tmp00_81_21;
	wire [WIDTH*2-1+0:0] tmp00_81_22;
	wire [WIDTH*2-1+0:0] tmp00_81_23;
	wire [WIDTH*2-1+0:0] tmp00_81_24;
	wire [WIDTH*2-1+0:0] tmp00_81_25;
	wire [WIDTH*2-1+0:0] tmp00_81_26;
	wire [WIDTH*2-1+0:0] tmp00_81_27;
	wire [WIDTH*2-1+0:0] tmp00_81_28;
	wire [WIDTH*2-1+0:0] tmp00_81_29;
	wire [WIDTH*2-1+0:0] tmp00_81_30;
	wire [WIDTH*2-1+0:0] tmp00_81_31;
	wire [WIDTH*2-1+0:0] tmp00_81_32;
	wire [WIDTH*2-1+0:0] tmp00_81_33;
	wire [WIDTH*2-1+0:0] tmp00_81_34;
	wire [WIDTH*2-1+0:0] tmp00_81_35;
	wire [WIDTH*2-1+0:0] tmp00_81_36;
	wire [WIDTH*2-1+0:0] tmp00_81_37;
	wire [WIDTH*2-1+0:0] tmp00_81_38;
	wire [WIDTH*2-1+0:0] tmp00_81_39;
	wire [WIDTH*2-1+0:0] tmp00_81_40;
	wire [WIDTH*2-1+0:0] tmp00_81_41;
	wire [WIDTH*2-1+0:0] tmp00_81_42;
	wire [WIDTH*2-1+0:0] tmp00_81_43;
	wire [WIDTH*2-1+0:0] tmp00_81_44;
	wire [WIDTH*2-1+0:0] tmp00_81_45;
	wire [WIDTH*2-1+0:0] tmp00_81_46;
	wire [WIDTH*2-1+0:0] tmp00_81_47;
	wire [WIDTH*2-1+0:0] tmp00_81_48;
	wire [WIDTH*2-1+0:0] tmp00_81_49;
	wire [WIDTH*2-1+0:0] tmp00_81_50;
	wire [WIDTH*2-1+0:0] tmp00_81_51;
	wire [WIDTH*2-1+0:0] tmp00_81_52;
	wire [WIDTH*2-1+0:0] tmp00_81_53;
	wire [WIDTH*2-1+0:0] tmp00_81_54;
	wire [WIDTH*2-1+0:0] tmp00_81_55;
	wire [WIDTH*2-1+0:0] tmp00_81_56;
	wire [WIDTH*2-1+0:0] tmp00_81_57;
	wire [WIDTH*2-1+0:0] tmp00_81_58;
	wire [WIDTH*2-1+0:0] tmp00_81_59;
	wire [WIDTH*2-1+0:0] tmp00_81_60;
	wire [WIDTH*2-1+0:0] tmp00_81_61;
	wire [WIDTH*2-1+0:0] tmp00_81_62;
	wire [WIDTH*2-1+0:0] tmp00_81_63;
	wire [WIDTH*2-1+0:0] tmp00_81_64;
	wire [WIDTH*2-1+0:0] tmp00_81_65;
	wire [WIDTH*2-1+0:0] tmp00_81_66;
	wire [WIDTH*2-1+0:0] tmp00_81_67;
	wire [WIDTH*2-1+0:0] tmp00_81_68;
	wire [WIDTH*2-1+0:0] tmp00_81_69;
	wire [WIDTH*2-1+0:0] tmp00_81_70;
	wire [WIDTH*2-1+0:0] tmp00_81_71;
	wire [WIDTH*2-1+0:0] tmp00_81_72;
	wire [WIDTH*2-1+0:0] tmp00_81_73;
	wire [WIDTH*2-1+0:0] tmp00_81_74;
	wire [WIDTH*2-1+0:0] tmp00_81_75;
	wire [WIDTH*2-1+0:0] tmp00_81_76;
	wire [WIDTH*2-1+0:0] tmp00_81_77;
	wire [WIDTH*2-1+0:0] tmp00_81_78;
	wire [WIDTH*2-1+0:0] tmp00_81_79;
	wire [WIDTH*2-1+0:0] tmp00_81_80;
	wire [WIDTH*2-1+0:0] tmp00_81_81;
	wire [WIDTH*2-1+0:0] tmp00_81_82;
	wire [WIDTH*2-1+0:0] tmp00_81_83;
	wire [WIDTH*2-1+0:0] tmp00_82_0;
	wire [WIDTH*2-1+0:0] tmp00_82_1;
	wire [WIDTH*2-1+0:0] tmp00_82_2;
	wire [WIDTH*2-1+0:0] tmp00_82_3;
	wire [WIDTH*2-1+0:0] tmp00_82_4;
	wire [WIDTH*2-1+0:0] tmp00_82_5;
	wire [WIDTH*2-1+0:0] tmp00_82_6;
	wire [WIDTH*2-1+0:0] tmp00_82_7;
	wire [WIDTH*2-1+0:0] tmp00_82_8;
	wire [WIDTH*2-1+0:0] tmp00_82_9;
	wire [WIDTH*2-1+0:0] tmp00_82_10;
	wire [WIDTH*2-1+0:0] tmp00_82_11;
	wire [WIDTH*2-1+0:0] tmp00_82_12;
	wire [WIDTH*2-1+0:0] tmp00_82_13;
	wire [WIDTH*2-1+0:0] tmp00_82_14;
	wire [WIDTH*2-1+0:0] tmp00_82_15;
	wire [WIDTH*2-1+0:0] tmp00_82_16;
	wire [WIDTH*2-1+0:0] tmp00_82_17;
	wire [WIDTH*2-1+0:0] tmp00_82_18;
	wire [WIDTH*2-1+0:0] tmp00_82_19;
	wire [WIDTH*2-1+0:0] tmp00_82_20;
	wire [WIDTH*2-1+0:0] tmp00_82_21;
	wire [WIDTH*2-1+0:0] tmp00_82_22;
	wire [WIDTH*2-1+0:0] tmp00_82_23;
	wire [WIDTH*2-1+0:0] tmp00_82_24;
	wire [WIDTH*2-1+0:0] tmp00_82_25;
	wire [WIDTH*2-1+0:0] tmp00_82_26;
	wire [WIDTH*2-1+0:0] tmp00_82_27;
	wire [WIDTH*2-1+0:0] tmp00_82_28;
	wire [WIDTH*2-1+0:0] tmp00_82_29;
	wire [WIDTH*2-1+0:0] tmp00_82_30;
	wire [WIDTH*2-1+0:0] tmp00_82_31;
	wire [WIDTH*2-1+0:0] tmp00_82_32;
	wire [WIDTH*2-1+0:0] tmp00_82_33;
	wire [WIDTH*2-1+0:0] tmp00_82_34;
	wire [WIDTH*2-1+0:0] tmp00_82_35;
	wire [WIDTH*2-1+0:0] tmp00_82_36;
	wire [WIDTH*2-1+0:0] tmp00_82_37;
	wire [WIDTH*2-1+0:0] tmp00_82_38;
	wire [WIDTH*2-1+0:0] tmp00_82_39;
	wire [WIDTH*2-1+0:0] tmp00_82_40;
	wire [WIDTH*2-1+0:0] tmp00_82_41;
	wire [WIDTH*2-1+0:0] tmp00_82_42;
	wire [WIDTH*2-1+0:0] tmp00_82_43;
	wire [WIDTH*2-1+0:0] tmp00_82_44;
	wire [WIDTH*2-1+0:0] tmp00_82_45;
	wire [WIDTH*2-1+0:0] tmp00_82_46;
	wire [WIDTH*2-1+0:0] tmp00_82_47;
	wire [WIDTH*2-1+0:0] tmp00_82_48;
	wire [WIDTH*2-1+0:0] tmp00_82_49;
	wire [WIDTH*2-1+0:0] tmp00_82_50;
	wire [WIDTH*2-1+0:0] tmp00_82_51;
	wire [WIDTH*2-1+0:0] tmp00_82_52;
	wire [WIDTH*2-1+0:0] tmp00_82_53;
	wire [WIDTH*2-1+0:0] tmp00_82_54;
	wire [WIDTH*2-1+0:0] tmp00_82_55;
	wire [WIDTH*2-1+0:0] tmp00_82_56;
	wire [WIDTH*2-1+0:0] tmp00_82_57;
	wire [WIDTH*2-1+0:0] tmp00_82_58;
	wire [WIDTH*2-1+0:0] tmp00_82_59;
	wire [WIDTH*2-1+0:0] tmp00_82_60;
	wire [WIDTH*2-1+0:0] tmp00_82_61;
	wire [WIDTH*2-1+0:0] tmp00_82_62;
	wire [WIDTH*2-1+0:0] tmp00_82_63;
	wire [WIDTH*2-1+0:0] tmp00_82_64;
	wire [WIDTH*2-1+0:0] tmp00_82_65;
	wire [WIDTH*2-1+0:0] tmp00_82_66;
	wire [WIDTH*2-1+0:0] tmp00_82_67;
	wire [WIDTH*2-1+0:0] tmp00_82_68;
	wire [WIDTH*2-1+0:0] tmp00_82_69;
	wire [WIDTH*2-1+0:0] tmp00_82_70;
	wire [WIDTH*2-1+0:0] tmp00_82_71;
	wire [WIDTH*2-1+0:0] tmp00_82_72;
	wire [WIDTH*2-1+0:0] tmp00_82_73;
	wire [WIDTH*2-1+0:0] tmp00_82_74;
	wire [WIDTH*2-1+0:0] tmp00_82_75;
	wire [WIDTH*2-1+0:0] tmp00_82_76;
	wire [WIDTH*2-1+0:0] tmp00_82_77;
	wire [WIDTH*2-1+0:0] tmp00_82_78;
	wire [WIDTH*2-1+0:0] tmp00_82_79;
	wire [WIDTH*2-1+0:0] tmp00_82_80;
	wire [WIDTH*2-1+0:0] tmp00_82_81;
	wire [WIDTH*2-1+0:0] tmp00_82_82;
	wire [WIDTH*2-1+0:0] tmp00_82_83;
	wire [WIDTH*2-1+0:0] tmp00_83_0;
	wire [WIDTH*2-1+0:0] tmp00_83_1;
	wire [WIDTH*2-1+0:0] tmp00_83_2;
	wire [WIDTH*2-1+0:0] tmp00_83_3;
	wire [WIDTH*2-1+0:0] tmp00_83_4;
	wire [WIDTH*2-1+0:0] tmp00_83_5;
	wire [WIDTH*2-1+0:0] tmp00_83_6;
	wire [WIDTH*2-1+0:0] tmp00_83_7;
	wire [WIDTH*2-1+0:0] tmp00_83_8;
	wire [WIDTH*2-1+0:0] tmp00_83_9;
	wire [WIDTH*2-1+0:0] tmp00_83_10;
	wire [WIDTH*2-1+0:0] tmp00_83_11;
	wire [WIDTH*2-1+0:0] tmp00_83_12;
	wire [WIDTH*2-1+0:0] tmp00_83_13;
	wire [WIDTH*2-1+0:0] tmp00_83_14;
	wire [WIDTH*2-1+0:0] tmp00_83_15;
	wire [WIDTH*2-1+0:0] tmp00_83_16;
	wire [WIDTH*2-1+0:0] tmp00_83_17;
	wire [WIDTH*2-1+0:0] tmp00_83_18;
	wire [WIDTH*2-1+0:0] tmp00_83_19;
	wire [WIDTH*2-1+0:0] tmp00_83_20;
	wire [WIDTH*2-1+0:0] tmp00_83_21;
	wire [WIDTH*2-1+0:0] tmp00_83_22;
	wire [WIDTH*2-1+0:0] tmp00_83_23;
	wire [WIDTH*2-1+0:0] tmp00_83_24;
	wire [WIDTH*2-1+0:0] tmp00_83_25;
	wire [WIDTH*2-1+0:0] tmp00_83_26;
	wire [WIDTH*2-1+0:0] tmp00_83_27;
	wire [WIDTH*2-1+0:0] tmp00_83_28;
	wire [WIDTH*2-1+0:0] tmp00_83_29;
	wire [WIDTH*2-1+0:0] tmp00_83_30;
	wire [WIDTH*2-1+0:0] tmp00_83_31;
	wire [WIDTH*2-1+0:0] tmp00_83_32;
	wire [WIDTH*2-1+0:0] tmp00_83_33;
	wire [WIDTH*2-1+0:0] tmp00_83_34;
	wire [WIDTH*2-1+0:0] tmp00_83_35;
	wire [WIDTH*2-1+0:0] tmp00_83_36;
	wire [WIDTH*2-1+0:0] tmp00_83_37;
	wire [WIDTH*2-1+0:0] tmp00_83_38;
	wire [WIDTH*2-1+0:0] tmp00_83_39;
	wire [WIDTH*2-1+0:0] tmp00_83_40;
	wire [WIDTH*2-1+0:0] tmp00_83_41;
	wire [WIDTH*2-1+0:0] tmp00_83_42;
	wire [WIDTH*2-1+0:0] tmp00_83_43;
	wire [WIDTH*2-1+0:0] tmp00_83_44;
	wire [WIDTH*2-1+0:0] tmp00_83_45;
	wire [WIDTH*2-1+0:0] tmp00_83_46;
	wire [WIDTH*2-1+0:0] tmp00_83_47;
	wire [WIDTH*2-1+0:0] tmp00_83_48;
	wire [WIDTH*2-1+0:0] tmp00_83_49;
	wire [WIDTH*2-1+0:0] tmp00_83_50;
	wire [WIDTH*2-1+0:0] tmp00_83_51;
	wire [WIDTH*2-1+0:0] tmp00_83_52;
	wire [WIDTH*2-1+0:0] tmp00_83_53;
	wire [WIDTH*2-1+0:0] tmp00_83_54;
	wire [WIDTH*2-1+0:0] tmp00_83_55;
	wire [WIDTH*2-1+0:0] tmp00_83_56;
	wire [WIDTH*2-1+0:0] tmp00_83_57;
	wire [WIDTH*2-1+0:0] tmp00_83_58;
	wire [WIDTH*2-1+0:0] tmp00_83_59;
	wire [WIDTH*2-1+0:0] tmp00_83_60;
	wire [WIDTH*2-1+0:0] tmp00_83_61;
	wire [WIDTH*2-1+0:0] tmp00_83_62;
	wire [WIDTH*2-1+0:0] tmp00_83_63;
	wire [WIDTH*2-1+0:0] tmp00_83_64;
	wire [WIDTH*2-1+0:0] tmp00_83_65;
	wire [WIDTH*2-1+0:0] tmp00_83_66;
	wire [WIDTH*2-1+0:0] tmp00_83_67;
	wire [WIDTH*2-1+0:0] tmp00_83_68;
	wire [WIDTH*2-1+0:0] tmp00_83_69;
	wire [WIDTH*2-1+0:0] tmp00_83_70;
	wire [WIDTH*2-1+0:0] tmp00_83_71;
	wire [WIDTH*2-1+0:0] tmp00_83_72;
	wire [WIDTH*2-1+0:0] tmp00_83_73;
	wire [WIDTH*2-1+0:0] tmp00_83_74;
	wire [WIDTH*2-1+0:0] tmp00_83_75;
	wire [WIDTH*2-1+0:0] tmp00_83_76;
	wire [WIDTH*2-1+0:0] tmp00_83_77;
	wire [WIDTH*2-1+0:0] tmp00_83_78;
	wire [WIDTH*2-1+0:0] tmp00_83_79;
	wire [WIDTH*2-1+0:0] tmp00_83_80;
	wire [WIDTH*2-1+0:0] tmp00_83_81;
	wire [WIDTH*2-1+0:0] tmp00_83_82;
	wire [WIDTH*2-1+0:0] tmp00_83_83;
	wire [WIDTH*2-1+0:0] tmp00_84_0;
	wire [WIDTH*2-1+0:0] tmp00_84_1;
	wire [WIDTH*2-1+0:0] tmp00_84_2;
	wire [WIDTH*2-1+0:0] tmp00_84_3;
	wire [WIDTH*2-1+0:0] tmp00_84_4;
	wire [WIDTH*2-1+0:0] tmp00_84_5;
	wire [WIDTH*2-1+0:0] tmp00_84_6;
	wire [WIDTH*2-1+0:0] tmp00_84_7;
	wire [WIDTH*2-1+0:0] tmp00_84_8;
	wire [WIDTH*2-1+0:0] tmp00_84_9;
	wire [WIDTH*2-1+0:0] tmp00_84_10;
	wire [WIDTH*2-1+0:0] tmp00_84_11;
	wire [WIDTH*2-1+0:0] tmp00_84_12;
	wire [WIDTH*2-1+0:0] tmp00_84_13;
	wire [WIDTH*2-1+0:0] tmp00_84_14;
	wire [WIDTH*2-1+0:0] tmp00_84_15;
	wire [WIDTH*2-1+0:0] tmp00_84_16;
	wire [WIDTH*2-1+0:0] tmp00_84_17;
	wire [WIDTH*2-1+0:0] tmp00_84_18;
	wire [WIDTH*2-1+0:0] tmp00_84_19;
	wire [WIDTH*2-1+0:0] tmp00_84_20;
	wire [WIDTH*2-1+0:0] tmp00_84_21;
	wire [WIDTH*2-1+0:0] tmp00_84_22;
	wire [WIDTH*2-1+0:0] tmp00_84_23;
	wire [WIDTH*2-1+0:0] tmp00_84_24;
	wire [WIDTH*2-1+0:0] tmp00_84_25;
	wire [WIDTH*2-1+0:0] tmp00_84_26;
	wire [WIDTH*2-1+0:0] tmp00_84_27;
	wire [WIDTH*2-1+0:0] tmp00_84_28;
	wire [WIDTH*2-1+0:0] tmp00_84_29;
	wire [WIDTH*2-1+0:0] tmp00_84_30;
	wire [WIDTH*2-1+0:0] tmp00_84_31;
	wire [WIDTH*2-1+0:0] tmp00_84_32;
	wire [WIDTH*2-1+0:0] tmp00_84_33;
	wire [WIDTH*2-1+0:0] tmp00_84_34;
	wire [WIDTH*2-1+0:0] tmp00_84_35;
	wire [WIDTH*2-1+0:0] tmp00_84_36;
	wire [WIDTH*2-1+0:0] tmp00_84_37;
	wire [WIDTH*2-1+0:0] tmp00_84_38;
	wire [WIDTH*2-1+0:0] tmp00_84_39;
	wire [WIDTH*2-1+0:0] tmp00_84_40;
	wire [WIDTH*2-1+0:0] tmp00_84_41;
	wire [WIDTH*2-1+0:0] tmp00_84_42;
	wire [WIDTH*2-1+0:0] tmp00_84_43;
	wire [WIDTH*2-1+0:0] tmp00_84_44;
	wire [WIDTH*2-1+0:0] tmp00_84_45;
	wire [WIDTH*2-1+0:0] tmp00_84_46;
	wire [WIDTH*2-1+0:0] tmp00_84_47;
	wire [WIDTH*2-1+0:0] tmp00_84_48;
	wire [WIDTH*2-1+0:0] tmp00_84_49;
	wire [WIDTH*2-1+0:0] tmp00_84_50;
	wire [WIDTH*2-1+0:0] tmp00_84_51;
	wire [WIDTH*2-1+0:0] tmp00_84_52;
	wire [WIDTH*2-1+0:0] tmp00_84_53;
	wire [WIDTH*2-1+0:0] tmp00_84_54;
	wire [WIDTH*2-1+0:0] tmp00_84_55;
	wire [WIDTH*2-1+0:0] tmp00_84_56;
	wire [WIDTH*2-1+0:0] tmp00_84_57;
	wire [WIDTH*2-1+0:0] tmp00_84_58;
	wire [WIDTH*2-1+0:0] tmp00_84_59;
	wire [WIDTH*2-1+0:0] tmp00_84_60;
	wire [WIDTH*2-1+0:0] tmp00_84_61;
	wire [WIDTH*2-1+0:0] tmp00_84_62;
	wire [WIDTH*2-1+0:0] tmp00_84_63;
	wire [WIDTH*2-1+0:0] tmp00_84_64;
	wire [WIDTH*2-1+0:0] tmp00_84_65;
	wire [WIDTH*2-1+0:0] tmp00_84_66;
	wire [WIDTH*2-1+0:0] tmp00_84_67;
	wire [WIDTH*2-1+0:0] tmp00_84_68;
	wire [WIDTH*2-1+0:0] tmp00_84_69;
	wire [WIDTH*2-1+0:0] tmp00_84_70;
	wire [WIDTH*2-1+0:0] tmp00_84_71;
	wire [WIDTH*2-1+0:0] tmp00_84_72;
	wire [WIDTH*2-1+0:0] tmp00_84_73;
	wire [WIDTH*2-1+0:0] tmp00_84_74;
	wire [WIDTH*2-1+0:0] tmp00_84_75;
	wire [WIDTH*2-1+0:0] tmp00_84_76;
	wire [WIDTH*2-1+0:0] tmp00_84_77;
	wire [WIDTH*2-1+0:0] tmp00_84_78;
	wire [WIDTH*2-1+0:0] tmp00_84_79;
	wire [WIDTH*2-1+0:0] tmp00_84_80;
	wire [WIDTH*2-1+0:0] tmp00_84_81;
	wire [WIDTH*2-1+0:0] tmp00_84_82;
	wire [WIDTH*2-1+0:0] tmp00_84_83;
	wire [WIDTH*2-1+0:0] tmp00_85_0;
	wire [WIDTH*2-1+0:0] tmp00_85_1;
	wire [WIDTH*2-1+0:0] tmp00_85_2;
	wire [WIDTH*2-1+0:0] tmp00_85_3;
	wire [WIDTH*2-1+0:0] tmp00_85_4;
	wire [WIDTH*2-1+0:0] tmp00_85_5;
	wire [WIDTH*2-1+0:0] tmp00_85_6;
	wire [WIDTH*2-1+0:0] tmp00_85_7;
	wire [WIDTH*2-1+0:0] tmp00_85_8;
	wire [WIDTH*2-1+0:0] tmp00_85_9;
	wire [WIDTH*2-1+0:0] tmp00_85_10;
	wire [WIDTH*2-1+0:0] tmp00_85_11;
	wire [WIDTH*2-1+0:0] tmp00_85_12;
	wire [WIDTH*2-1+0:0] tmp00_85_13;
	wire [WIDTH*2-1+0:0] tmp00_85_14;
	wire [WIDTH*2-1+0:0] tmp00_85_15;
	wire [WIDTH*2-1+0:0] tmp00_85_16;
	wire [WIDTH*2-1+0:0] tmp00_85_17;
	wire [WIDTH*2-1+0:0] tmp00_85_18;
	wire [WIDTH*2-1+0:0] tmp00_85_19;
	wire [WIDTH*2-1+0:0] tmp00_85_20;
	wire [WIDTH*2-1+0:0] tmp00_85_21;
	wire [WIDTH*2-1+0:0] tmp00_85_22;
	wire [WIDTH*2-1+0:0] tmp00_85_23;
	wire [WIDTH*2-1+0:0] tmp00_85_24;
	wire [WIDTH*2-1+0:0] tmp00_85_25;
	wire [WIDTH*2-1+0:0] tmp00_85_26;
	wire [WIDTH*2-1+0:0] tmp00_85_27;
	wire [WIDTH*2-1+0:0] tmp00_85_28;
	wire [WIDTH*2-1+0:0] tmp00_85_29;
	wire [WIDTH*2-1+0:0] tmp00_85_30;
	wire [WIDTH*2-1+0:0] tmp00_85_31;
	wire [WIDTH*2-1+0:0] tmp00_85_32;
	wire [WIDTH*2-1+0:0] tmp00_85_33;
	wire [WIDTH*2-1+0:0] tmp00_85_34;
	wire [WIDTH*2-1+0:0] tmp00_85_35;
	wire [WIDTH*2-1+0:0] tmp00_85_36;
	wire [WIDTH*2-1+0:0] tmp00_85_37;
	wire [WIDTH*2-1+0:0] tmp00_85_38;
	wire [WIDTH*2-1+0:0] tmp00_85_39;
	wire [WIDTH*2-1+0:0] tmp00_85_40;
	wire [WIDTH*2-1+0:0] tmp00_85_41;
	wire [WIDTH*2-1+0:0] tmp00_85_42;
	wire [WIDTH*2-1+0:0] tmp00_85_43;
	wire [WIDTH*2-1+0:0] tmp00_85_44;
	wire [WIDTH*2-1+0:0] tmp00_85_45;
	wire [WIDTH*2-1+0:0] tmp00_85_46;
	wire [WIDTH*2-1+0:0] tmp00_85_47;
	wire [WIDTH*2-1+0:0] tmp00_85_48;
	wire [WIDTH*2-1+0:0] tmp00_85_49;
	wire [WIDTH*2-1+0:0] tmp00_85_50;
	wire [WIDTH*2-1+0:0] tmp00_85_51;
	wire [WIDTH*2-1+0:0] tmp00_85_52;
	wire [WIDTH*2-1+0:0] tmp00_85_53;
	wire [WIDTH*2-1+0:0] tmp00_85_54;
	wire [WIDTH*2-1+0:0] tmp00_85_55;
	wire [WIDTH*2-1+0:0] tmp00_85_56;
	wire [WIDTH*2-1+0:0] tmp00_85_57;
	wire [WIDTH*2-1+0:0] tmp00_85_58;
	wire [WIDTH*2-1+0:0] tmp00_85_59;
	wire [WIDTH*2-1+0:0] tmp00_85_60;
	wire [WIDTH*2-1+0:0] tmp00_85_61;
	wire [WIDTH*2-1+0:0] tmp00_85_62;
	wire [WIDTH*2-1+0:0] tmp00_85_63;
	wire [WIDTH*2-1+0:0] tmp00_85_64;
	wire [WIDTH*2-1+0:0] tmp00_85_65;
	wire [WIDTH*2-1+0:0] tmp00_85_66;
	wire [WIDTH*2-1+0:0] tmp00_85_67;
	wire [WIDTH*2-1+0:0] tmp00_85_68;
	wire [WIDTH*2-1+0:0] tmp00_85_69;
	wire [WIDTH*2-1+0:0] tmp00_85_70;
	wire [WIDTH*2-1+0:0] tmp00_85_71;
	wire [WIDTH*2-1+0:0] tmp00_85_72;
	wire [WIDTH*2-1+0:0] tmp00_85_73;
	wire [WIDTH*2-1+0:0] tmp00_85_74;
	wire [WIDTH*2-1+0:0] tmp00_85_75;
	wire [WIDTH*2-1+0:0] tmp00_85_76;
	wire [WIDTH*2-1+0:0] tmp00_85_77;
	wire [WIDTH*2-1+0:0] tmp00_85_78;
	wire [WIDTH*2-1+0:0] tmp00_85_79;
	wire [WIDTH*2-1+0:0] tmp00_85_80;
	wire [WIDTH*2-1+0:0] tmp00_85_81;
	wire [WIDTH*2-1+0:0] tmp00_85_82;
	wire [WIDTH*2-1+0:0] tmp00_85_83;
	wire [WIDTH*2-1+0:0] tmp00_86_0;
	wire [WIDTH*2-1+0:0] tmp00_86_1;
	wire [WIDTH*2-1+0:0] tmp00_86_2;
	wire [WIDTH*2-1+0:0] tmp00_86_3;
	wire [WIDTH*2-1+0:0] tmp00_86_4;
	wire [WIDTH*2-1+0:0] tmp00_86_5;
	wire [WIDTH*2-1+0:0] tmp00_86_6;
	wire [WIDTH*2-1+0:0] tmp00_86_7;
	wire [WIDTH*2-1+0:0] tmp00_86_8;
	wire [WIDTH*2-1+0:0] tmp00_86_9;
	wire [WIDTH*2-1+0:0] tmp00_86_10;
	wire [WIDTH*2-1+0:0] tmp00_86_11;
	wire [WIDTH*2-1+0:0] tmp00_86_12;
	wire [WIDTH*2-1+0:0] tmp00_86_13;
	wire [WIDTH*2-1+0:0] tmp00_86_14;
	wire [WIDTH*2-1+0:0] tmp00_86_15;
	wire [WIDTH*2-1+0:0] tmp00_86_16;
	wire [WIDTH*2-1+0:0] tmp00_86_17;
	wire [WIDTH*2-1+0:0] tmp00_86_18;
	wire [WIDTH*2-1+0:0] tmp00_86_19;
	wire [WIDTH*2-1+0:0] tmp00_86_20;
	wire [WIDTH*2-1+0:0] tmp00_86_21;
	wire [WIDTH*2-1+0:0] tmp00_86_22;
	wire [WIDTH*2-1+0:0] tmp00_86_23;
	wire [WIDTH*2-1+0:0] tmp00_86_24;
	wire [WIDTH*2-1+0:0] tmp00_86_25;
	wire [WIDTH*2-1+0:0] tmp00_86_26;
	wire [WIDTH*2-1+0:0] tmp00_86_27;
	wire [WIDTH*2-1+0:0] tmp00_86_28;
	wire [WIDTH*2-1+0:0] tmp00_86_29;
	wire [WIDTH*2-1+0:0] tmp00_86_30;
	wire [WIDTH*2-1+0:0] tmp00_86_31;
	wire [WIDTH*2-1+0:0] tmp00_86_32;
	wire [WIDTH*2-1+0:0] tmp00_86_33;
	wire [WIDTH*2-1+0:0] tmp00_86_34;
	wire [WIDTH*2-1+0:0] tmp00_86_35;
	wire [WIDTH*2-1+0:0] tmp00_86_36;
	wire [WIDTH*2-1+0:0] tmp00_86_37;
	wire [WIDTH*2-1+0:0] tmp00_86_38;
	wire [WIDTH*2-1+0:0] tmp00_86_39;
	wire [WIDTH*2-1+0:0] tmp00_86_40;
	wire [WIDTH*2-1+0:0] tmp00_86_41;
	wire [WIDTH*2-1+0:0] tmp00_86_42;
	wire [WIDTH*2-1+0:0] tmp00_86_43;
	wire [WIDTH*2-1+0:0] tmp00_86_44;
	wire [WIDTH*2-1+0:0] tmp00_86_45;
	wire [WIDTH*2-1+0:0] tmp00_86_46;
	wire [WIDTH*2-1+0:0] tmp00_86_47;
	wire [WIDTH*2-1+0:0] tmp00_86_48;
	wire [WIDTH*2-1+0:0] tmp00_86_49;
	wire [WIDTH*2-1+0:0] tmp00_86_50;
	wire [WIDTH*2-1+0:0] tmp00_86_51;
	wire [WIDTH*2-1+0:0] tmp00_86_52;
	wire [WIDTH*2-1+0:0] tmp00_86_53;
	wire [WIDTH*2-1+0:0] tmp00_86_54;
	wire [WIDTH*2-1+0:0] tmp00_86_55;
	wire [WIDTH*2-1+0:0] tmp00_86_56;
	wire [WIDTH*2-1+0:0] tmp00_86_57;
	wire [WIDTH*2-1+0:0] tmp00_86_58;
	wire [WIDTH*2-1+0:0] tmp00_86_59;
	wire [WIDTH*2-1+0:0] tmp00_86_60;
	wire [WIDTH*2-1+0:0] tmp00_86_61;
	wire [WIDTH*2-1+0:0] tmp00_86_62;
	wire [WIDTH*2-1+0:0] tmp00_86_63;
	wire [WIDTH*2-1+0:0] tmp00_86_64;
	wire [WIDTH*2-1+0:0] tmp00_86_65;
	wire [WIDTH*2-1+0:0] tmp00_86_66;
	wire [WIDTH*2-1+0:0] tmp00_86_67;
	wire [WIDTH*2-1+0:0] tmp00_86_68;
	wire [WIDTH*2-1+0:0] tmp00_86_69;
	wire [WIDTH*2-1+0:0] tmp00_86_70;
	wire [WIDTH*2-1+0:0] tmp00_86_71;
	wire [WIDTH*2-1+0:0] tmp00_86_72;
	wire [WIDTH*2-1+0:0] tmp00_86_73;
	wire [WIDTH*2-1+0:0] tmp00_86_74;
	wire [WIDTH*2-1+0:0] tmp00_86_75;
	wire [WIDTH*2-1+0:0] tmp00_86_76;
	wire [WIDTH*2-1+0:0] tmp00_86_77;
	wire [WIDTH*2-1+0:0] tmp00_86_78;
	wire [WIDTH*2-1+0:0] tmp00_86_79;
	wire [WIDTH*2-1+0:0] tmp00_86_80;
	wire [WIDTH*2-1+0:0] tmp00_86_81;
	wire [WIDTH*2-1+0:0] tmp00_86_82;
	wire [WIDTH*2-1+0:0] tmp00_86_83;
	wire [WIDTH*2-1+0:0] tmp00_87_0;
	wire [WIDTH*2-1+0:0] tmp00_87_1;
	wire [WIDTH*2-1+0:0] tmp00_87_2;
	wire [WIDTH*2-1+0:0] tmp00_87_3;
	wire [WIDTH*2-1+0:0] tmp00_87_4;
	wire [WIDTH*2-1+0:0] tmp00_87_5;
	wire [WIDTH*2-1+0:0] tmp00_87_6;
	wire [WIDTH*2-1+0:0] tmp00_87_7;
	wire [WIDTH*2-1+0:0] tmp00_87_8;
	wire [WIDTH*2-1+0:0] tmp00_87_9;
	wire [WIDTH*2-1+0:0] tmp00_87_10;
	wire [WIDTH*2-1+0:0] tmp00_87_11;
	wire [WIDTH*2-1+0:0] tmp00_87_12;
	wire [WIDTH*2-1+0:0] tmp00_87_13;
	wire [WIDTH*2-1+0:0] tmp00_87_14;
	wire [WIDTH*2-1+0:0] tmp00_87_15;
	wire [WIDTH*2-1+0:0] tmp00_87_16;
	wire [WIDTH*2-1+0:0] tmp00_87_17;
	wire [WIDTH*2-1+0:0] tmp00_87_18;
	wire [WIDTH*2-1+0:0] tmp00_87_19;
	wire [WIDTH*2-1+0:0] tmp00_87_20;
	wire [WIDTH*2-1+0:0] tmp00_87_21;
	wire [WIDTH*2-1+0:0] tmp00_87_22;
	wire [WIDTH*2-1+0:0] tmp00_87_23;
	wire [WIDTH*2-1+0:0] tmp00_87_24;
	wire [WIDTH*2-1+0:0] tmp00_87_25;
	wire [WIDTH*2-1+0:0] tmp00_87_26;
	wire [WIDTH*2-1+0:0] tmp00_87_27;
	wire [WIDTH*2-1+0:0] tmp00_87_28;
	wire [WIDTH*2-1+0:0] tmp00_87_29;
	wire [WIDTH*2-1+0:0] tmp00_87_30;
	wire [WIDTH*2-1+0:0] tmp00_87_31;
	wire [WIDTH*2-1+0:0] tmp00_87_32;
	wire [WIDTH*2-1+0:0] tmp00_87_33;
	wire [WIDTH*2-1+0:0] tmp00_87_34;
	wire [WIDTH*2-1+0:0] tmp00_87_35;
	wire [WIDTH*2-1+0:0] tmp00_87_36;
	wire [WIDTH*2-1+0:0] tmp00_87_37;
	wire [WIDTH*2-1+0:0] tmp00_87_38;
	wire [WIDTH*2-1+0:0] tmp00_87_39;
	wire [WIDTH*2-1+0:0] tmp00_87_40;
	wire [WIDTH*2-1+0:0] tmp00_87_41;
	wire [WIDTH*2-1+0:0] tmp00_87_42;
	wire [WIDTH*2-1+0:0] tmp00_87_43;
	wire [WIDTH*2-1+0:0] tmp00_87_44;
	wire [WIDTH*2-1+0:0] tmp00_87_45;
	wire [WIDTH*2-1+0:0] tmp00_87_46;
	wire [WIDTH*2-1+0:0] tmp00_87_47;
	wire [WIDTH*2-1+0:0] tmp00_87_48;
	wire [WIDTH*2-1+0:0] tmp00_87_49;
	wire [WIDTH*2-1+0:0] tmp00_87_50;
	wire [WIDTH*2-1+0:0] tmp00_87_51;
	wire [WIDTH*2-1+0:0] tmp00_87_52;
	wire [WIDTH*2-1+0:0] tmp00_87_53;
	wire [WIDTH*2-1+0:0] tmp00_87_54;
	wire [WIDTH*2-1+0:0] tmp00_87_55;
	wire [WIDTH*2-1+0:0] tmp00_87_56;
	wire [WIDTH*2-1+0:0] tmp00_87_57;
	wire [WIDTH*2-1+0:0] tmp00_87_58;
	wire [WIDTH*2-1+0:0] tmp00_87_59;
	wire [WIDTH*2-1+0:0] tmp00_87_60;
	wire [WIDTH*2-1+0:0] tmp00_87_61;
	wire [WIDTH*2-1+0:0] tmp00_87_62;
	wire [WIDTH*2-1+0:0] tmp00_87_63;
	wire [WIDTH*2-1+0:0] tmp00_87_64;
	wire [WIDTH*2-1+0:0] tmp00_87_65;
	wire [WIDTH*2-1+0:0] tmp00_87_66;
	wire [WIDTH*2-1+0:0] tmp00_87_67;
	wire [WIDTH*2-1+0:0] tmp00_87_68;
	wire [WIDTH*2-1+0:0] tmp00_87_69;
	wire [WIDTH*2-1+0:0] tmp00_87_70;
	wire [WIDTH*2-1+0:0] tmp00_87_71;
	wire [WIDTH*2-1+0:0] tmp00_87_72;
	wire [WIDTH*2-1+0:0] tmp00_87_73;
	wire [WIDTH*2-1+0:0] tmp00_87_74;
	wire [WIDTH*2-1+0:0] tmp00_87_75;
	wire [WIDTH*2-1+0:0] tmp00_87_76;
	wire [WIDTH*2-1+0:0] tmp00_87_77;
	wire [WIDTH*2-1+0:0] tmp00_87_78;
	wire [WIDTH*2-1+0:0] tmp00_87_79;
	wire [WIDTH*2-1+0:0] tmp00_87_80;
	wire [WIDTH*2-1+0:0] tmp00_87_81;
	wire [WIDTH*2-1+0:0] tmp00_87_82;
	wire [WIDTH*2-1+0:0] tmp00_87_83;
	wire [WIDTH*2-1+0:0] tmp00_88_0;
	wire [WIDTH*2-1+0:0] tmp00_88_1;
	wire [WIDTH*2-1+0:0] tmp00_88_2;
	wire [WIDTH*2-1+0:0] tmp00_88_3;
	wire [WIDTH*2-1+0:0] tmp00_88_4;
	wire [WIDTH*2-1+0:0] tmp00_88_5;
	wire [WIDTH*2-1+0:0] tmp00_88_6;
	wire [WIDTH*2-1+0:0] tmp00_88_7;
	wire [WIDTH*2-1+0:0] tmp00_88_8;
	wire [WIDTH*2-1+0:0] tmp00_88_9;
	wire [WIDTH*2-1+0:0] tmp00_88_10;
	wire [WIDTH*2-1+0:0] tmp00_88_11;
	wire [WIDTH*2-1+0:0] tmp00_88_12;
	wire [WIDTH*2-1+0:0] tmp00_88_13;
	wire [WIDTH*2-1+0:0] tmp00_88_14;
	wire [WIDTH*2-1+0:0] tmp00_88_15;
	wire [WIDTH*2-1+0:0] tmp00_88_16;
	wire [WIDTH*2-1+0:0] tmp00_88_17;
	wire [WIDTH*2-1+0:0] tmp00_88_18;
	wire [WIDTH*2-1+0:0] tmp00_88_19;
	wire [WIDTH*2-1+0:0] tmp00_88_20;
	wire [WIDTH*2-1+0:0] tmp00_88_21;
	wire [WIDTH*2-1+0:0] tmp00_88_22;
	wire [WIDTH*2-1+0:0] tmp00_88_23;
	wire [WIDTH*2-1+0:0] tmp00_88_24;
	wire [WIDTH*2-1+0:0] tmp00_88_25;
	wire [WIDTH*2-1+0:0] tmp00_88_26;
	wire [WIDTH*2-1+0:0] tmp00_88_27;
	wire [WIDTH*2-1+0:0] tmp00_88_28;
	wire [WIDTH*2-1+0:0] tmp00_88_29;
	wire [WIDTH*2-1+0:0] tmp00_88_30;
	wire [WIDTH*2-1+0:0] tmp00_88_31;
	wire [WIDTH*2-1+0:0] tmp00_88_32;
	wire [WIDTH*2-1+0:0] tmp00_88_33;
	wire [WIDTH*2-1+0:0] tmp00_88_34;
	wire [WIDTH*2-1+0:0] tmp00_88_35;
	wire [WIDTH*2-1+0:0] tmp00_88_36;
	wire [WIDTH*2-1+0:0] tmp00_88_37;
	wire [WIDTH*2-1+0:0] tmp00_88_38;
	wire [WIDTH*2-1+0:0] tmp00_88_39;
	wire [WIDTH*2-1+0:0] tmp00_88_40;
	wire [WIDTH*2-1+0:0] tmp00_88_41;
	wire [WIDTH*2-1+0:0] tmp00_88_42;
	wire [WIDTH*2-1+0:0] tmp00_88_43;
	wire [WIDTH*2-1+0:0] tmp00_88_44;
	wire [WIDTH*2-1+0:0] tmp00_88_45;
	wire [WIDTH*2-1+0:0] tmp00_88_46;
	wire [WIDTH*2-1+0:0] tmp00_88_47;
	wire [WIDTH*2-1+0:0] tmp00_88_48;
	wire [WIDTH*2-1+0:0] tmp00_88_49;
	wire [WIDTH*2-1+0:0] tmp00_88_50;
	wire [WIDTH*2-1+0:0] tmp00_88_51;
	wire [WIDTH*2-1+0:0] tmp00_88_52;
	wire [WIDTH*2-1+0:0] tmp00_88_53;
	wire [WIDTH*2-1+0:0] tmp00_88_54;
	wire [WIDTH*2-1+0:0] tmp00_88_55;
	wire [WIDTH*2-1+0:0] tmp00_88_56;
	wire [WIDTH*2-1+0:0] tmp00_88_57;
	wire [WIDTH*2-1+0:0] tmp00_88_58;
	wire [WIDTH*2-1+0:0] tmp00_88_59;
	wire [WIDTH*2-1+0:0] tmp00_88_60;
	wire [WIDTH*2-1+0:0] tmp00_88_61;
	wire [WIDTH*2-1+0:0] tmp00_88_62;
	wire [WIDTH*2-1+0:0] tmp00_88_63;
	wire [WIDTH*2-1+0:0] tmp00_88_64;
	wire [WIDTH*2-1+0:0] tmp00_88_65;
	wire [WIDTH*2-1+0:0] tmp00_88_66;
	wire [WIDTH*2-1+0:0] tmp00_88_67;
	wire [WIDTH*2-1+0:0] tmp00_88_68;
	wire [WIDTH*2-1+0:0] tmp00_88_69;
	wire [WIDTH*2-1+0:0] tmp00_88_70;
	wire [WIDTH*2-1+0:0] tmp00_88_71;
	wire [WIDTH*2-1+0:0] tmp00_88_72;
	wire [WIDTH*2-1+0:0] tmp00_88_73;
	wire [WIDTH*2-1+0:0] tmp00_88_74;
	wire [WIDTH*2-1+0:0] tmp00_88_75;
	wire [WIDTH*2-1+0:0] tmp00_88_76;
	wire [WIDTH*2-1+0:0] tmp00_88_77;
	wire [WIDTH*2-1+0:0] tmp00_88_78;
	wire [WIDTH*2-1+0:0] tmp00_88_79;
	wire [WIDTH*2-1+0:0] tmp00_88_80;
	wire [WIDTH*2-1+0:0] tmp00_88_81;
	wire [WIDTH*2-1+0:0] tmp00_88_82;
	wire [WIDTH*2-1+0:0] tmp00_88_83;
	wire [WIDTH*2-1+0:0] tmp00_89_0;
	wire [WIDTH*2-1+0:0] tmp00_89_1;
	wire [WIDTH*2-1+0:0] tmp00_89_2;
	wire [WIDTH*2-1+0:0] tmp00_89_3;
	wire [WIDTH*2-1+0:0] tmp00_89_4;
	wire [WIDTH*2-1+0:0] tmp00_89_5;
	wire [WIDTH*2-1+0:0] tmp00_89_6;
	wire [WIDTH*2-1+0:0] tmp00_89_7;
	wire [WIDTH*2-1+0:0] tmp00_89_8;
	wire [WIDTH*2-1+0:0] tmp00_89_9;
	wire [WIDTH*2-1+0:0] tmp00_89_10;
	wire [WIDTH*2-1+0:0] tmp00_89_11;
	wire [WIDTH*2-1+0:0] tmp00_89_12;
	wire [WIDTH*2-1+0:0] tmp00_89_13;
	wire [WIDTH*2-1+0:0] tmp00_89_14;
	wire [WIDTH*2-1+0:0] tmp00_89_15;
	wire [WIDTH*2-1+0:0] tmp00_89_16;
	wire [WIDTH*2-1+0:0] tmp00_89_17;
	wire [WIDTH*2-1+0:0] tmp00_89_18;
	wire [WIDTH*2-1+0:0] tmp00_89_19;
	wire [WIDTH*2-1+0:0] tmp00_89_20;
	wire [WIDTH*2-1+0:0] tmp00_89_21;
	wire [WIDTH*2-1+0:0] tmp00_89_22;
	wire [WIDTH*2-1+0:0] tmp00_89_23;
	wire [WIDTH*2-1+0:0] tmp00_89_24;
	wire [WIDTH*2-1+0:0] tmp00_89_25;
	wire [WIDTH*2-1+0:0] tmp00_89_26;
	wire [WIDTH*2-1+0:0] tmp00_89_27;
	wire [WIDTH*2-1+0:0] tmp00_89_28;
	wire [WIDTH*2-1+0:0] tmp00_89_29;
	wire [WIDTH*2-1+0:0] tmp00_89_30;
	wire [WIDTH*2-1+0:0] tmp00_89_31;
	wire [WIDTH*2-1+0:0] tmp00_89_32;
	wire [WIDTH*2-1+0:0] tmp00_89_33;
	wire [WIDTH*2-1+0:0] tmp00_89_34;
	wire [WIDTH*2-1+0:0] tmp00_89_35;
	wire [WIDTH*2-1+0:0] tmp00_89_36;
	wire [WIDTH*2-1+0:0] tmp00_89_37;
	wire [WIDTH*2-1+0:0] tmp00_89_38;
	wire [WIDTH*2-1+0:0] tmp00_89_39;
	wire [WIDTH*2-1+0:0] tmp00_89_40;
	wire [WIDTH*2-1+0:0] tmp00_89_41;
	wire [WIDTH*2-1+0:0] tmp00_89_42;
	wire [WIDTH*2-1+0:0] tmp00_89_43;
	wire [WIDTH*2-1+0:0] tmp00_89_44;
	wire [WIDTH*2-1+0:0] tmp00_89_45;
	wire [WIDTH*2-1+0:0] tmp00_89_46;
	wire [WIDTH*2-1+0:0] tmp00_89_47;
	wire [WIDTH*2-1+0:0] tmp00_89_48;
	wire [WIDTH*2-1+0:0] tmp00_89_49;
	wire [WIDTH*2-1+0:0] tmp00_89_50;
	wire [WIDTH*2-1+0:0] tmp00_89_51;
	wire [WIDTH*2-1+0:0] tmp00_89_52;
	wire [WIDTH*2-1+0:0] tmp00_89_53;
	wire [WIDTH*2-1+0:0] tmp00_89_54;
	wire [WIDTH*2-1+0:0] tmp00_89_55;
	wire [WIDTH*2-1+0:0] tmp00_89_56;
	wire [WIDTH*2-1+0:0] tmp00_89_57;
	wire [WIDTH*2-1+0:0] tmp00_89_58;
	wire [WIDTH*2-1+0:0] tmp00_89_59;
	wire [WIDTH*2-1+0:0] tmp00_89_60;
	wire [WIDTH*2-1+0:0] tmp00_89_61;
	wire [WIDTH*2-1+0:0] tmp00_89_62;
	wire [WIDTH*2-1+0:0] tmp00_89_63;
	wire [WIDTH*2-1+0:0] tmp00_89_64;
	wire [WIDTH*2-1+0:0] tmp00_89_65;
	wire [WIDTH*2-1+0:0] tmp00_89_66;
	wire [WIDTH*2-1+0:0] tmp00_89_67;
	wire [WIDTH*2-1+0:0] tmp00_89_68;
	wire [WIDTH*2-1+0:0] tmp00_89_69;
	wire [WIDTH*2-1+0:0] tmp00_89_70;
	wire [WIDTH*2-1+0:0] tmp00_89_71;
	wire [WIDTH*2-1+0:0] tmp00_89_72;
	wire [WIDTH*2-1+0:0] tmp00_89_73;
	wire [WIDTH*2-1+0:0] tmp00_89_74;
	wire [WIDTH*2-1+0:0] tmp00_89_75;
	wire [WIDTH*2-1+0:0] tmp00_89_76;
	wire [WIDTH*2-1+0:0] tmp00_89_77;
	wire [WIDTH*2-1+0:0] tmp00_89_78;
	wire [WIDTH*2-1+0:0] tmp00_89_79;
	wire [WIDTH*2-1+0:0] tmp00_89_80;
	wire [WIDTH*2-1+0:0] tmp00_89_81;
	wire [WIDTH*2-1+0:0] tmp00_89_82;
	wire [WIDTH*2-1+0:0] tmp00_89_83;
	wire [WIDTH*2-1+0:0] tmp00_90_0;
	wire [WIDTH*2-1+0:0] tmp00_90_1;
	wire [WIDTH*2-1+0:0] tmp00_90_2;
	wire [WIDTH*2-1+0:0] tmp00_90_3;
	wire [WIDTH*2-1+0:0] tmp00_90_4;
	wire [WIDTH*2-1+0:0] tmp00_90_5;
	wire [WIDTH*2-1+0:0] tmp00_90_6;
	wire [WIDTH*2-1+0:0] tmp00_90_7;
	wire [WIDTH*2-1+0:0] tmp00_90_8;
	wire [WIDTH*2-1+0:0] tmp00_90_9;
	wire [WIDTH*2-1+0:0] tmp00_90_10;
	wire [WIDTH*2-1+0:0] tmp00_90_11;
	wire [WIDTH*2-1+0:0] tmp00_90_12;
	wire [WIDTH*2-1+0:0] tmp00_90_13;
	wire [WIDTH*2-1+0:0] tmp00_90_14;
	wire [WIDTH*2-1+0:0] tmp00_90_15;
	wire [WIDTH*2-1+0:0] tmp00_90_16;
	wire [WIDTH*2-1+0:0] tmp00_90_17;
	wire [WIDTH*2-1+0:0] tmp00_90_18;
	wire [WIDTH*2-1+0:0] tmp00_90_19;
	wire [WIDTH*2-1+0:0] tmp00_90_20;
	wire [WIDTH*2-1+0:0] tmp00_90_21;
	wire [WIDTH*2-1+0:0] tmp00_90_22;
	wire [WIDTH*2-1+0:0] tmp00_90_23;
	wire [WIDTH*2-1+0:0] tmp00_90_24;
	wire [WIDTH*2-1+0:0] tmp00_90_25;
	wire [WIDTH*2-1+0:0] tmp00_90_26;
	wire [WIDTH*2-1+0:0] tmp00_90_27;
	wire [WIDTH*2-1+0:0] tmp00_90_28;
	wire [WIDTH*2-1+0:0] tmp00_90_29;
	wire [WIDTH*2-1+0:0] tmp00_90_30;
	wire [WIDTH*2-1+0:0] tmp00_90_31;
	wire [WIDTH*2-1+0:0] tmp00_90_32;
	wire [WIDTH*2-1+0:0] tmp00_90_33;
	wire [WIDTH*2-1+0:0] tmp00_90_34;
	wire [WIDTH*2-1+0:0] tmp00_90_35;
	wire [WIDTH*2-1+0:0] tmp00_90_36;
	wire [WIDTH*2-1+0:0] tmp00_90_37;
	wire [WIDTH*2-1+0:0] tmp00_90_38;
	wire [WIDTH*2-1+0:0] tmp00_90_39;
	wire [WIDTH*2-1+0:0] tmp00_90_40;
	wire [WIDTH*2-1+0:0] tmp00_90_41;
	wire [WIDTH*2-1+0:0] tmp00_90_42;
	wire [WIDTH*2-1+0:0] tmp00_90_43;
	wire [WIDTH*2-1+0:0] tmp00_90_44;
	wire [WIDTH*2-1+0:0] tmp00_90_45;
	wire [WIDTH*2-1+0:0] tmp00_90_46;
	wire [WIDTH*2-1+0:0] tmp00_90_47;
	wire [WIDTH*2-1+0:0] tmp00_90_48;
	wire [WIDTH*2-1+0:0] tmp00_90_49;
	wire [WIDTH*2-1+0:0] tmp00_90_50;
	wire [WIDTH*2-1+0:0] tmp00_90_51;
	wire [WIDTH*2-1+0:0] tmp00_90_52;
	wire [WIDTH*2-1+0:0] tmp00_90_53;
	wire [WIDTH*2-1+0:0] tmp00_90_54;
	wire [WIDTH*2-1+0:0] tmp00_90_55;
	wire [WIDTH*2-1+0:0] tmp00_90_56;
	wire [WIDTH*2-1+0:0] tmp00_90_57;
	wire [WIDTH*2-1+0:0] tmp00_90_58;
	wire [WIDTH*2-1+0:0] tmp00_90_59;
	wire [WIDTH*2-1+0:0] tmp00_90_60;
	wire [WIDTH*2-1+0:0] tmp00_90_61;
	wire [WIDTH*2-1+0:0] tmp00_90_62;
	wire [WIDTH*2-1+0:0] tmp00_90_63;
	wire [WIDTH*2-1+0:0] tmp00_90_64;
	wire [WIDTH*2-1+0:0] tmp00_90_65;
	wire [WIDTH*2-1+0:0] tmp00_90_66;
	wire [WIDTH*2-1+0:0] tmp00_90_67;
	wire [WIDTH*2-1+0:0] tmp00_90_68;
	wire [WIDTH*2-1+0:0] tmp00_90_69;
	wire [WIDTH*2-1+0:0] tmp00_90_70;
	wire [WIDTH*2-1+0:0] tmp00_90_71;
	wire [WIDTH*2-1+0:0] tmp00_90_72;
	wire [WIDTH*2-1+0:0] tmp00_90_73;
	wire [WIDTH*2-1+0:0] tmp00_90_74;
	wire [WIDTH*2-1+0:0] tmp00_90_75;
	wire [WIDTH*2-1+0:0] tmp00_90_76;
	wire [WIDTH*2-1+0:0] tmp00_90_77;
	wire [WIDTH*2-1+0:0] tmp00_90_78;
	wire [WIDTH*2-1+0:0] tmp00_90_79;
	wire [WIDTH*2-1+0:0] tmp00_90_80;
	wire [WIDTH*2-1+0:0] tmp00_90_81;
	wire [WIDTH*2-1+0:0] tmp00_90_82;
	wire [WIDTH*2-1+0:0] tmp00_90_83;
	wire [WIDTH*2-1+0:0] tmp00_91_0;
	wire [WIDTH*2-1+0:0] tmp00_91_1;
	wire [WIDTH*2-1+0:0] tmp00_91_2;
	wire [WIDTH*2-1+0:0] tmp00_91_3;
	wire [WIDTH*2-1+0:0] tmp00_91_4;
	wire [WIDTH*2-1+0:0] tmp00_91_5;
	wire [WIDTH*2-1+0:0] tmp00_91_6;
	wire [WIDTH*2-1+0:0] tmp00_91_7;
	wire [WIDTH*2-1+0:0] tmp00_91_8;
	wire [WIDTH*2-1+0:0] tmp00_91_9;
	wire [WIDTH*2-1+0:0] tmp00_91_10;
	wire [WIDTH*2-1+0:0] tmp00_91_11;
	wire [WIDTH*2-1+0:0] tmp00_91_12;
	wire [WIDTH*2-1+0:0] tmp00_91_13;
	wire [WIDTH*2-1+0:0] tmp00_91_14;
	wire [WIDTH*2-1+0:0] tmp00_91_15;
	wire [WIDTH*2-1+0:0] tmp00_91_16;
	wire [WIDTH*2-1+0:0] tmp00_91_17;
	wire [WIDTH*2-1+0:0] tmp00_91_18;
	wire [WIDTH*2-1+0:0] tmp00_91_19;
	wire [WIDTH*2-1+0:0] tmp00_91_20;
	wire [WIDTH*2-1+0:0] tmp00_91_21;
	wire [WIDTH*2-1+0:0] tmp00_91_22;
	wire [WIDTH*2-1+0:0] tmp00_91_23;
	wire [WIDTH*2-1+0:0] tmp00_91_24;
	wire [WIDTH*2-1+0:0] tmp00_91_25;
	wire [WIDTH*2-1+0:0] tmp00_91_26;
	wire [WIDTH*2-1+0:0] tmp00_91_27;
	wire [WIDTH*2-1+0:0] tmp00_91_28;
	wire [WIDTH*2-1+0:0] tmp00_91_29;
	wire [WIDTH*2-1+0:0] tmp00_91_30;
	wire [WIDTH*2-1+0:0] tmp00_91_31;
	wire [WIDTH*2-1+0:0] tmp00_91_32;
	wire [WIDTH*2-1+0:0] tmp00_91_33;
	wire [WIDTH*2-1+0:0] tmp00_91_34;
	wire [WIDTH*2-1+0:0] tmp00_91_35;
	wire [WIDTH*2-1+0:0] tmp00_91_36;
	wire [WIDTH*2-1+0:0] tmp00_91_37;
	wire [WIDTH*2-1+0:0] tmp00_91_38;
	wire [WIDTH*2-1+0:0] tmp00_91_39;
	wire [WIDTH*2-1+0:0] tmp00_91_40;
	wire [WIDTH*2-1+0:0] tmp00_91_41;
	wire [WIDTH*2-1+0:0] tmp00_91_42;
	wire [WIDTH*2-1+0:0] tmp00_91_43;
	wire [WIDTH*2-1+0:0] tmp00_91_44;
	wire [WIDTH*2-1+0:0] tmp00_91_45;
	wire [WIDTH*2-1+0:0] tmp00_91_46;
	wire [WIDTH*2-1+0:0] tmp00_91_47;
	wire [WIDTH*2-1+0:0] tmp00_91_48;
	wire [WIDTH*2-1+0:0] tmp00_91_49;
	wire [WIDTH*2-1+0:0] tmp00_91_50;
	wire [WIDTH*2-1+0:0] tmp00_91_51;
	wire [WIDTH*2-1+0:0] tmp00_91_52;
	wire [WIDTH*2-1+0:0] tmp00_91_53;
	wire [WIDTH*2-1+0:0] tmp00_91_54;
	wire [WIDTH*2-1+0:0] tmp00_91_55;
	wire [WIDTH*2-1+0:0] tmp00_91_56;
	wire [WIDTH*2-1+0:0] tmp00_91_57;
	wire [WIDTH*2-1+0:0] tmp00_91_58;
	wire [WIDTH*2-1+0:0] tmp00_91_59;
	wire [WIDTH*2-1+0:0] tmp00_91_60;
	wire [WIDTH*2-1+0:0] tmp00_91_61;
	wire [WIDTH*2-1+0:0] tmp00_91_62;
	wire [WIDTH*2-1+0:0] tmp00_91_63;
	wire [WIDTH*2-1+0:0] tmp00_91_64;
	wire [WIDTH*2-1+0:0] tmp00_91_65;
	wire [WIDTH*2-1+0:0] tmp00_91_66;
	wire [WIDTH*2-1+0:0] tmp00_91_67;
	wire [WIDTH*2-1+0:0] tmp00_91_68;
	wire [WIDTH*2-1+0:0] tmp00_91_69;
	wire [WIDTH*2-1+0:0] tmp00_91_70;
	wire [WIDTH*2-1+0:0] tmp00_91_71;
	wire [WIDTH*2-1+0:0] tmp00_91_72;
	wire [WIDTH*2-1+0:0] tmp00_91_73;
	wire [WIDTH*2-1+0:0] tmp00_91_74;
	wire [WIDTH*2-1+0:0] tmp00_91_75;
	wire [WIDTH*2-1+0:0] tmp00_91_76;
	wire [WIDTH*2-1+0:0] tmp00_91_77;
	wire [WIDTH*2-1+0:0] tmp00_91_78;
	wire [WIDTH*2-1+0:0] tmp00_91_79;
	wire [WIDTH*2-1+0:0] tmp00_91_80;
	wire [WIDTH*2-1+0:0] tmp00_91_81;
	wire [WIDTH*2-1+0:0] tmp00_91_82;
	wire [WIDTH*2-1+0:0] tmp00_91_83;
	wire [WIDTH*2-1+0:0] tmp00_92_0;
	wire [WIDTH*2-1+0:0] tmp00_92_1;
	wire [WIDTH*2-1+0:0] tmp00_92_2;
	wire [WIDTH*2-1+0:0] tmp00_92_3;
	wire [WIDTH*2-1+0:0] tmp00_92_4;
	wire [WIDTH*2-1+0:0] tmp00_92_5;
	wire [WIDTH*2-1+0:0] tmp00_92_6;
	wire [WIDTH*2-1+0:0] tmp00_92_7;
	wire [WIDTH*2-1+0:0] tmp00_92_8;
	wire [WIDTH*2-1+0:0] tmp00_92_9;
	wire [WIDTH*2-1+0:0] tmp00_92_10;
	wire [WIDTH*2-1+0:0] tmp00_92_11;
	wire [WIDTH*2-1+0:0] tmp00_92_12;
	wire [WIDTH*2-1+0:0] tmp00_92_13;
	wire [WIDTH*2-1+0:0] tmp00_92_14;
	wire [WIDTH*2-1+0:0] tmp00_92_15;
	wire [WIDTH*2-1+0:0] tmp00_92_16;
	wire [WIDTH*2-1+0:0] tmp00_92_17;
	wire [WIDTH*2-1+0:0] tmp00_92_18;
	wire [WIDTH*2-1+0:0] tmp00_92_19;
	wire [WIDTH*2-1+0:0] tmp00_92_20;
	wire [WIDTH*2-1+0:0] tmp00_92_21;
	wire [WIDTH*2-1+0:0] tmp00_92_22;
	wire [WIDTH*2-1+0:0] tmp00_92_23;
	wire [WIDTH*2-1+0:0] tmp00_92_24;
	wire [WIDTH*2-1+0:0] tmp00_92_25;
	wire [WIDTH*2-1+0:0] tmp00_92_26;
	wire [WIDTH*2-1+0:0] tmp00_92_27;
	wire [WIDTH*2-1+0:0] tmp00_92_28;
	wire [WIDTH*2-1+0:0] tmp00_92_29;
	wire [WIDTH*2-1+0:0] tmp00_92_30;
	wire [WIDTH*2-1+0:0] tmp00_92_31;
	wire [WIDTH*2-1+0:0] tmp00_92_32;
	wire [WIDTH*2-1+0:0] tmp00_92_33;
	wire [WIDTH*2-1+0:0] tmp00_92_34;
	wire [WIDTH*2-1+0:0] tmp00_92_35;
	wire [WIDTH*2-1+0:0] tmp00_92_36;
	wire [WIDTH*2-1+0:0] tmp00_92_37;
	wire [WIDTH*2-1+0:0] tmp00_92_38;
	wire [WIDTH*2-1+0:0] tmp00_92_39;
	wire [WIDTH*2-1+0:0] tmp00_92_40;
	wire [WIDTH*2-1+0:0] tmp00_92_41;
	wire [WIDTH*2-1+0:0] tmp00_92_42;
	wire [WIDTH*2-1+0:0] tmp00_92_43;
	wire [WIDTH*2-1+0:0] tmp00_92_44;
	wire [WIDTH*2-1+0:0] tmp00_92_45;
	wire [WIDTH*2-1+0:0] tmp00_92_46;
	wire [WIDTH*2-1+0:0] tmp00_92_47;
	wire [WIDTH*2-1+0:0] tmp00_92_48;
	wire [WIDTH*2-1+0:0] tmp00_92_49;
	wire [WIDTH*2-1+0:0] tmp00_92_50;
	wire [WIDTH*2-1+0:0] tmp00_92_51;
	wire [WIDTH*2-1+0:0] tmp00_92_52;
	wire [WIDTH*2-1+0:0] tmp00_92_53;
	wire [WIDTH*2-1+0:0] tmp00_92_54;
	wire [WIDTH*2-1+0:0] tmp00_92_55;
	wire [WIDTH*2-1+0:0] tmp00_92_56;
	wire [WIDTH*2-1+0:0] tmp00_92_57;
	wire [WIDTH*2-1+0:0] tmp00_92_58;
	wire [WIDTH*2-1+0:0] tmp00_92_59;
	wire [WIDTH*2-1+0:0] tmp00_92_60;
	wire [WIDTH*2-1+0:0] tmp00_92_61;
	wire [WIDTH*2-1+0:0] tmp00_92_62;
	wire [WIDTH*2-1+0:0] tmp00_92_63;
	wire [WIDTH*2-1+0:0] tmp00_92_64;
	wire [WIDTH*2-1+0:0] tmp00_92_65;
	wire [WIDTH*2-1+0:0] tmp00_92_66;
	wire [WIDTH*2-1+0:0] tmp00_92_67;
	wire [WIDTH*2-1+0:0] tmp00_92_68;
	wire [WIDTH*2-1+0:0] tmp00_92_69;
	wire [WIDTH*2-1+0:0] tmp00_92_70;
	wire [WIDTH*2-1+0:0] tmp00_92_71;
	wire [WIDTH*2-1+0:0] tmp00_92_72;
	wire [WIDTH*2-1+0:0] tmp00_92_73;
	wire [WIDTH*2-1+0:0] tmp00_92_74;
	wire [WIDTH*2-1+0:0] tmp00_92_75;
	wire [WIDTH*2-1+0:0] tmp00_92_76;
	wire [WIDTH*2-1+0:0] tmp00_92_77;
	wire [WIDTH*2-1+0:0] tmp00_92_78;
	wire [WIDTH*2-1+0:0] tmp00_92_79;
	wire [WIDTH*2-1+0:0] tmp00_92_80;
	wire [WIDTH*2-1+0:0] tmp00_92_81;
	wire [WIDTH*2-1+0:0] tmp00_92_82;
	wire [WIDTH*2-1+0:0] tmp00_92_83;
	wire [WIDTH*2-1+0:0] tmp00_93_0;
	wire [WIDTH*2-1+0:0] tmp00_93_1;
	wire [WIDTH*2-1+0:0] tmp00_93_2;
	wire [WIDTH*2-1+0:0] tmp00_93_3;
	wire [WIDTH*2-1+0:0] tmp00_93_4;
	wire [WIDTH*2-1+0:0] tmp00_93_5;
	wire [WIDTH*2-1+0:0] tmp00_93_6;
	wire [WIDTH*2-1+0:0] tmp00_93_7;
	wire [WIDTH*2-1+0:0] tmp00_93_8;
	wire [WIDTH*2-1+0:0] tmp00_93_9;
	wire [WIDTH*2-1+0:0] tmp00_93_10;
	wire [WIDTH*2-1+0:0] tmp00_93_11;
	wire [WIDTH*2-1+0:0] tmp00_93_12;
	wire [WIDTH*2-1+0:0] tmp00_93_13;
	wire [WIDTH*2-1+0:0] tmp00_93_14;
	wire [WIDTH*2-1+0:0] tmp00_93_15;
	wire [WIDTH*2-1+0:0] tmp00_93_16;
	wire [WIDTH*2-1+0:0] tmp00_93_17;
	wire [WIDTH*2-1+0:0] tmp00_93_18;
	wire [WIDTH*2-1+0:0] tmp00_93_19;
	wire [WIDTH*2-1+0:0] tmp00_93_20;
	wire [WIDTH*2-1+0:0] tmp00_93_21;
	wire [WIDTH*2-1+0:0] tmp00_93_22;
	wire [WIDTH*2-1+0:0] tmp00_93_23;
	wire [WIDTH*2-1+0:0] tmp00_93_24;
	wire [WIDTH*2-1+0:0] tmp00_93_25;
	wire [WIDTH*2-1+0:0] tmp00_93_26;
	wire [WIDTH*2-1+0:0] tmp00_93_27;
	wire [WIDTH*2-1+0:0] tmp00_93_28;
	wire [WIDTH*2-1+0:0] tmp00_93_29;
	wire [WIDTH*2-1+0:0] tmp00_93_30;
	wire [WIDTH*2-1+0:0] tmp00_93_31;
	wire [WIDTH*2-1+0:0] tmp00_93_32;
	wire [WIDTH*2-1+0:0] tmp00_93_33;
	wire [WIDTH*2-1+0:0] tmp00_93_34;
	wire [WIDTH*2-1+0:0] tmp00_93_35;
	wire [WIDTH*2-1+0:0] tmp00_93_36;
	wire [WIDTH*2-1+0:0] tmp00_93_37;
	wire [WIDTH*2-1+0:0] tmp00_93_38;
	wire [WIDTH*2-1+0:0] tmp00_93_39;
	wire [WIDTH*2-1+0:0] tmp00_93_40;
	wire [WIDTH*2-1+0:0] tmp00_93_41;
	wire [WIDTH*2-1+0:0] tmp00_93_42;
	wire [WIDTH*2-1+0:0] tmp00_93_43;
	wire [WIDTH*2-1+0:0] tmp00_93_44;
	wire [WIDTH*2-1+0:0] tmp00_93_45;
	wire [WIDTH*2-1+0:0] tmp00_93_46;
	wire [WIDTH*2-1+0:0] tmp00_93_47;
	wire [WIDTH*2-1+0:0] tmp00_93_48;
	wire [WIDTH*2-1+0:0] tmp00_93_49;
	wire [WIDTH*2-1+0:0] tmp00_93_50;
	wire [WIDTH*2-1+0:0] tmp00_93_51;
	wire [WIDTH*2-1+0:0] tmp00_93_52;
	wire [WIDTH*2-1+0:0] tmp00_93_53;
	wire [WIDTH*2-1+0:0] tmp00_93_54;
	wire [WIDTH*2-1+0:0] tmp00_93_55;
	wire [WIDTH*2-1+0:0] tmp00_93_56;
	wire [WIDTH*2-1+0:0] tmp00_93_57;
	wire [WIDTH*2-1+0:0] tmp00_93_58;
	wire [WIDTH*2-1+0:0] tmp00_93_59;
	wire [WIDTH*2-1+0:0] tmp00_93_60;
	wire [WIDTH*2-1+0:0] tmp00_93_61;
	wire [WIDTH*2-1+0:0] tmp00_93_62;
	wire [WIDTH*2-1+0:0] tmp00_93_63;
	wire [WIDTH*2-1+0:0] tmp00_93_64;
	wire [WIDTH*2-1+0:0] tmp00_93_65;
	wire [WIDTH*2-1+0:0] tmp00_93_66;
	wire [WIDTH*2-1+0:0] tmp00_93_67;
	wire [WIDTH*2-1+0:0] tmp00_93_68;
	wire [WIDTH*2-1+0:0] tmp00_93_69;
	wire [WIDTH*2-1+0:0] tmp00_93_70;
	wire [WIDTH*2-1+0:0] tmp00_93_71;
	wire [WIDTH*2-1+0:0] tmp00_93_72;
	wire [WIDTH*2-1+0:0] tmp00_93_73;
	wire [WIDTH*2-1+0:0] tmp00_93_74;
	wire [WIDTH*2-1+0:0] tmp00_93_75;
	wire [WIDTH*2-1+0:0] tmp00_93_76;
	wire [WIDTH*2-1+0:0] tmp00_93_77;
	wire [WIDTH*2-1+0:0] tmp00_93_78;
	wire [WIDTH*2-1+0:0] tmp00_93_79;
	wire [WIDTH*2-1+0:0] tmp00_93_80;
	wire [WIDTH*2-1+0:0] tmp00_93_81;
	wire [WIDTH*2-1+0:0] tmp00_93_82;
	wire [WIDTH*2-1+0:0] tmp00_93_83;
	wire [WIDTH*2-1+0:0] tmp00_94_0;
	wire [WIDTH*2-1+0:0] tmp00_94_1;
	wire [WIDTH*2-1+0:0] tmp00_94_2;
	wire [WIDTH*2-1+0:0] tmp00_94_3;
	wire [WIDTH*2-1+0:0] tmp00_94_4;
	wire [WIDTH*2-1+0:0] tmp00_94_5;
	wire [WIDTH*2-1+0:0] tmp00_94_6;
	wire [WIDTH*2-1+0:0] tmp00_94_7;
	wire [WIDTH*2-1+0:0] tmp00_94_8;
	wire [WIDTH*2-1+0:0] tmp00_94_9;
	wire [WIDTH*2-1+0:0] tmp00_94_10;
	wire [WIDTH*2-1+0:0] tmp00_94_11;
	wire [WIDTH*2-1+0:0] tmp00_94_12;
	wire [WIDTH*2-1+0:0] tmp00_94_13;
	wire [WIDTH*2-1+0:0] tmp00_94_14;
	wire [WIDTH*2-1+0:0] tmp00_94_15;
	wire [WIDTH*2-1+0:0] tmp00_94_16;
	wire [WIDTH*2-1+0:0] tmp00_94_17;
	wire [WIDTH*2-1+0:0] tmp00_94_18;
	wire [WIDTH*2-1+0:0] tmp00_94_19;
	wire [WIDTH*2-1+0:0] tmp00_94_20;
	wire [WIDTH*2-1+0:0] tmp00_94_21;
	wire [WIDTH*2-1+0:0] tmp00_94_22;
	wire [WIDTH*2-1+0:0] tmp00_94_23;
	wire [WIDTH*2-1+0:0] tmp00_94_24;
	wire [WIDTH*2-1+0:0] tmp00_94_25;
	wire [WIDTH*2-1+0:0] tmp00_94_26;
	wire [WIDTH*2-1+0:0] tmp00_94_27;
	wire [WIDTH*2-1+0:0] tmp00_94_28;
	wire [WIDTH*2-1+0:0] tmp00_94_29;
	wire [WIDTH*2-1+0:0] tmp00_94_30;
	wire [WIDTH*2-1+0:0] tmp00_94_31;
	wire [WIDTH*2-1+0:0] tmp00_94_32;
	wire [WIDTH*2-1+0:0] tmp00_94_33;
	wire [WIDTH*2-1+0:0] tmp00_94_34;
	wire [WIDTH*2-1+0:0] tmp00_94_35;
	wire [WIDTH*2-1+0:0] tmp00_94_36;
	wire [WIDTH*2-1+0:0] tmp00_94_37;
	wire [WIDTH*2-1+0:0] tmp00_94_38;
	wire [WIDTH*2-1+0:0] tmp00_94_39;
	wire [WIDTH*2-1+0:0] tmp00_94_40;
	wire [WIDTH*2-1+0:0] tmp00_94_41;
	wire [WIDTH*2-1+0:0] tmp00_94_42;
	wire [WIDTH*2-1+0:0] tmp00_94_43;
	wire [WIDTH*2-1+0:0] tmp00_94_44;
	wire [WIDTH*2-1+0:0] tmp00_94_45;
	wire [WIDTH*2-1+0:0] tmp00_94_46;
	wire [WIDTH*2-1+0:0] tmp00_94_47;
	wire [WIDTH*2-1+0:0] tmp00_94_48;
	wire [WIDTH*2-1+0:0] tmp00_94_49;
	wire [WIDTH*2-1+0:0] tmp00_94_50;
	wire [WIDTH*2-1+0:0] tmp00_94_51;
	wire [WIDTH*2-1+0:0] tmp00_94_52;
	wire [WIDTH*2-1+0:0] tmp00_94_53;
	wire [WIDTH*2-1+0:0] tmp00_94_54;
	wire [WIDTH*2-1+0:0] tmp00_94_55;
	wire [WIDTH*2-1+0:0] tmp00_94_56;
	wire [WIDTH*2-1+0:0] tmp00_94_57;
	wire [WIDTH*2-1+0:0] tmp00_94_58;
	wire [WIDTH*2-1+0:0] tmp00_94_59;
	wire [WIDTH*2-1+0:0] tmp00_94_60;
	wire [WIDTH*2-1+0:0] tmp00_94_61;
	wire [WIDTH*2-1+0:0] tmp00_94_62;
	wire [WIDTH*2-1+0:0] tmp00_94_63;
	wire [WIDTH*2-1+0:0] tmp00_94_64;
	wire [WIDTH*2-1+0:0] tmp00_94_65;
	wire [WIDTH*2-1+0:0] tmp00_94_66;
	wire [WIDTH*2-1+0:0] tmp00_94_67;
	wire [WIDTH*2-1+0:0] tmp00_94_68;
	wire [WIDTH*2-1+0:0] tmp00_94_69;
	wire [WIDTH*2-1+0:0] tmp00_94_70;
	wire [WIDTH*2-1+0:0] tmp00_94_71;
	wire [WIDTH*2-1+0:0] tmp00_94_72;
	wire [WIDTH*2-1+0:0] tmp00_94_73;
	wire [WIDTH*2-1+0:0] tmp00_94_74;
	wire [WIDTH*2-1+0:0] tmp00_94_75;
	wire [WIDTH*2-1+0:0] tmp00_94_76;
	wire [WIDTH*2-1+0:0] tmp00_94_77;
	wire [WIDTH*2-1+0:0] tmp00_94_78;
	wire [WIDTH*2-1+0:0] tmp00_94_79;
	wire [WIDTH*2-1+0:0] tmp00_94_80;
	wire [WIDTH*2-1+0:0] tmp00_94_81;
	wire [WIDTH*2-1+0:0] tmp00_94_82;
	wire [WIDTH*2-1+0:0] tmp00_94_83;
	wire [WIDTH*2-1+0:0] tmp00_95_0;
	wire [WIDTH*2-1+0:0] tmp00_95_1;
	wire [WIDTH*2-1+0:0] tmp00_95_2;
	wire [WIDTH*2-1+0:0] tmp00_95_3;
	wire [WIDTH*2-1+0:0] tmp00_95_4;
	wire [WIDTH*2-1+0:0] tmp00_95_5;
	wire [WIDTH*2-1+0:0] tmp00_95_6;
	wire [WIDTH*2-1+0:0] tmp00_95_7;
	wire [WIDTH*2-1+0:0] tmp00_95_8;
	wire [WIDTH*2-1+0:0] tmp00_95_9;
	wire [WIDTH*2-1+0:0] tmp00_95_10;
	wire [WIDTH*2-1+0:0] tmp00_95_11;
	wire [WIDTH*2-1+0:0] tmp00_95_12;
	wire [WIDTH*2-1+0:0] tmp00_95_13;
	wire [WIDTH*2-1+0:0] tmp00_95_14;
	wire [WIDTH*2-1+0:0] tmp00_95_15;
	wire [WIDTH*2-1+0:0] tmp00_95_16;
	wire [WIDTH*2-1+0:0] tmp00_95_17;
	wire [WIDTH*2-1+0:0] tmp00_95_18;
	wire [WIDTH*2-1+0:0] tmp00_95_19;
	wire [WIDTH*2-1+0:0] tmp00_95_20;
	wire [WIDTH*2-1+0:0] tmp00_95_21;
	wire [WIDTH*2-1+0:0] tmp00_95_22;
	wire [WIDTH*2-1+0:0] tmp00_95_23;
	wire [WIDTH*2-1+0:0] tmp00_95_24;
	wire [WIDTH*2-1+0:0] tmp00_95_25;
	wire [WIDTH*2-1+0:0] tmp00_95_26;
	wire [WIDTH*2-1+0:0] tmp00_95_27;
	wire [WIDTH*2-1+0:0] tmp00_95_28;
	wire [WIDTH*2-1+0:0] tmp00_95_29;
	wire [WIDTH*2-1+0:0] tmp00_95_30;
	wire [WIDTH*2-1+0:0] tmp00_95_31;
	wire [WIDTH*2-1+0:0] tmp00_95_32;
	wire [WIDTH*2-1+0:0] tmp00_95_33;
	wire [WIDTH*2-1+0:0] tmp00_95_34;
	wire [WIDTH*2-1+0:0] tmp00_95_35;
	wire [WIDTH*2-1+0:0] tmp00_95_36;
	wire [WIDTH*2-1+0:0] tmp00_95_37;
	wire [WIDTH*2-1+0:0] tmp00_95_38;
	wire [WIDTH*2-1+0:0] tmp00_95_39;
	wire [WIDTH*2-1+0:0] tmp00_95_40;
	wire [WIDTH*2-1+0:0] tmp00_95_41;
	wire [WIDTH*2-1+0:0] tmp00_95_42;
	wire [WIDTH*2-1+0:0] tmp00_95_43;
	wire [WIDTH*2-1+0:0] tmp00_95_44;
	wire [WIDTH*2-1+0:0] tmp00_95_45;
	wire [WIDTH*2-1+0:0] tmp00_95_46;
	wire [WIDTH*2-1+0:0] tmp00_95_47;
	wire [WIDTH*2-1+0:0] tmp00_95_48;
	wire [WIDTH*2-1+0:0] tmp00_95_49;
	wire [WIDTH*2-1+0:0] tmp00_95_50;
	wire [WIDTH*2-1+0:0] tmp00_95_51;
	wire [WIDTH*2-1+0:0] tmp00_95_52;
	wire [WIDTH*2-1+0:0] tmp00_95_53;
	wire [WIDTH*2-1+0:0] tmp00_95_54;
	wire [WIDTH*2-1+0:0] tmp00_95_55;
	wire [WIDTH*2-1+0:0] tmp00_95_56;
	wire [WIDTH*2-1+0:0] tmp00_95_57;
	wire [WIDTH*2-1+0:0] tmp00_95_58;
	wire [WIDTH*2-1+0:0] tmp00_95_59;
	wire [WIDTH*2-1+0:0] tmp00_95_60;
	wire [WIDTH*2-1+0:0] tmp00_95_61;
	wire [WIDTH*2-1+0:0] tmp00_95_62;
	wire [WIDTH*2-1+0:0] tmp00_95_63;
	wire [WIDTH*2-1+0:0] tmp00_95_64;
	wire [WIDTH*2-1+0:0] tmp00_95_65;
	wire [WIDTH*2-1+0:0] tmp00_95_66;
	wire [WIDTH*2-1+0:0] tmp00_95_67;
	wire [WIDTH*2-1+0:0] tmp00_95_68;
	wire [WIDTH*2-1+0:0] tmp00_95_69;
	wire [WIDTH*2-1+0:0] tmp00_95_70;
	wire [WIDTH*2-1+0:0] tmp00_95_71;
	wire [WIDTH*2-1+0:0] tmp00_95_72;
	wire [WIDTH*2-1+0:0] tmp00_95_73;
	wire [WIDTH*2-1+0:0] tmp00_95_74;
	wire [WIDTH*2-1+0:0] tmp00_95_75;
	wire [WIDTH*2-1+0:0] tmp00_95_76;
	wire [WIDTH*2-1+0:0] tmp00_95_77;
	wire [WIDTH*2-1+0:0] tmp00_95_78;
	wire [WIDTH*2-1+0:0] tmp00_95_79;
	wire [WIDTH*2-1+0:0] tmp00_95_80;
	wire [WIDTH*2-1+0:0] tmp00_95_81;
	wire [WIDTH*2-1+0:0] tmp00_95_82;
	wire [WIDTH*2-1+0:0] tmp00_95_83;
	wire [WIDTH*2-1+0:0] tmp00_96_0;
	wire [WIDTH*2-1+0:0] tmp00_96_1;
	wire [WIDTH*2-1+0:0] tmp00_96_2;
	wire [WIDTH*2-1+0:0] tmp00_96_3;
	wire [WIDTH*2-1+0:0] tmp00_96_4;
	wire [WIDTH*2-1+0:0] tmp00_96_5;
	wire [WIDTH*2-1+0:0] tmp00_96_6;
	wire [WIDTH*2-1+0:0] tmp00_96_7;
	wire [WIDTH*2-1+0:0] tmp00_96_8;
	wire [WIDTH*2-1+0:0] tmp00_96_9;
	wire [WIDTH*2-1+0:0] tmp00_96_10;
	wire [WIDTH*2-1+0:0] tmp00_96_11;
	wire [WIDTH*2-1+0:0] tmp00_96_12;
	wire [WIDTH*2-1+0:0] tmp00_96_13;
	wire [WIDTH*2-1+0:0] tmp00_96_14;
	wire [WIDTH*2-1+0:0] tmp00_96_15;
	wire [WIDTH*2-1+0:0] tmp00_96_16;
	wire [WIDTH*2-1+0:0] tmp00_96_17;
	wire [WIDTH*2-1+0:0] tmp00_96_18;
	wire [WIDTH*2-1+0:0] tmp00_96_19;
	wire [WIDTH*2-1+0:0] tmp00_96_20;
	wire [WIDTH*2-1+0:0] tmp00_96_21;
	wire [WIDTH*2-1+0:0] tmp00_96_22;
	wire [WIDTH*2-1+0:0] tmp00_96_23;
	wire [WIDTH*2-1+0:0] tmp00_96_24;
	wire [WIDTH*2-1+0:0] tmp00_96_25;
	wire [WIDTH*2-1+0:0] tmp00_96_26;
	wire [WIDTH*2-1+0:0] tmp00_96_27;
	wire [WIDTH*2-1+0:0] tmp00_96_28;
	wire [WIDTH*2-1+0:0] tmp00_96_29;
	wire [WIDTH*2-1+0:0] tmp00_96_30;
	wire [WIDTH*2-1+0:0] tmp00_96_31;
	wire [WIDTH*2-1+0:0] tmp00_96_32;
	wire [WIDTH*2-1+0:0] tmp00_96_33;
	wire [WIDTH*2-1+0:0] tmp00_96_34;
	wire [WIDTH*2-1+0:0] tmp00_96_35;
	wire [WIDTH*2-1+0:0] tmp00_96_36;
	wire [WIDTH*2-1+0:0] tmp00_96_37;
	wire [WIDTH*2-1+0:0] tmp00_96_38;
	wire [WIDTH*2-1+0:0] tmp00_96_39;
	wire [WIDTH*2-1+0:0] tmp00_96_40;
	wire [WIDTH*2-1+0:0] tmp00_96_41;
	wire [WIDTH*2-1+0:0] tmp00_96_42;
	wire [WIDTH*2-1+0:0] tmp00_96_43;
	wire [WIDTH*2-1+0:0] tmp00_96_44;
	wire [WIDTH*2-1+0:0] tmp00_96_45;
	wire [WIDTH*2-1+0:0] tmp00_96_46;
	wire [WIDTH*2-1+0:0] tmp00_96_47;
	wire [WIDTH*2-1+0:0] tmp00_96_48;
	wire [WIDTH*2-1+0:0] tmp00_96_49;
	wire [WIDTH*2-1+0:0] tmp00_96_50;
	wire [WIDTH*2-1+0:0] tmp00_96_51;
	wire [WIDTH*2-1+0:0] tmp00_96_52;
	wire [WIDTH*2-1+0:0] tmp00_96_53;
	wire [WIDTH*2-1+0:0] tmp00_96_54;
	wire [WIDTH*2-1+0:0] tmp00_96_55;
	wire [WIDTH*2-1+0:0] tmp00_96_56;
	wire [WIDTH*2-1+0:0] tmp00_96_57;
	wire [WIDTH*2-1+0:0] tmp00_96_58;
	wire [WIDTH*2-1+0:0] tmp00_96_59;
	wire [WIDTH*2-1+0:0] tmp00_96_60;
	wire [WIDTH*2-1+0:0] tmp00_96_61;
	wire [WIDTH*2-1+0:0] tmp00_96_62;
	wire [WIDTH*2-1+0:0] tmp00_96_63;
	wire [WIDTH*2-1+0:0] tmp00_96_64;
	wire [WIDTH*2-1+0:0] tmp00_96_65;
	wire [WIDTH*2-1+0:0] tmp00_96_66;
	wire [WIDTH*2-1+0:0] tmp00_96_67;
	wire [WIDTH*2-1+0:0] tmp00_96_68;
	wire [WIDTH*2-1+0:0] tmp00_96_69;
	wire [WIDTH*2-1+0:0] tmp00_96_70;
	wire [WIDTH*2-1+0:0] tmp00_96_71;
	wire [WIDTH*2-1+0:0] tmp00_96_72;
	wire [WIDTH*2-1+0:0] tmp00_96_73;
	wire [WIDTH*2-1+0:0] tmp00_96_74;
	wire [WIDTH*2-1+0:0] tmp00_96_75;
	wire [WIDTH*2-1+0:0] tmp00_96_76;
	wire [WIDTH*2-1+0:0] tmp00_96_77;
	wire [WIDTH*2-1+0:0] tmp00_96_78;
	wire [WIDTH*2-1+0:0] tmp00_96_79;
	wire [WIDTH*2-1+0:0] tmp00_96_80;
	wire [WIDTH*2-1+0:0] tmp00_96_81;
	wire [WIDTH*2-1+0:0] tmp00_96_82;
	wire [WIDTH*2-1+0:0] tmp00_96_83;
	wire [WIDTH*2-1+0:0] tmp00_97_0;
	wire [WIDTH*2-1+0:0] tmp00_97_1;
	wire [WIDTH*2-1+0:0] tmp00_97_2;
	wire [WIDTH*2-1+0:0] tmp00_97_3;
	wire [WIDTH*2-1+0:0] tmp00_97_4;
	wire [WIDTH*2-1+0:0] tmp00_97_5;
	wire [WIDTH*2-1+0:0] tmp00_97_6;
	wire [WIDTH*2-1+0:0] tmp00_97_7;
	wire [WIDTH*2-1+0:0] tmp00_97_8;
	wire [WIDTH*2-1+0:0] tmp00_97_9;
	wire [WIDTH*2-1+0:0] tmp00_97_10;
	wire [WIDTH*2-1+0:0] tmp00_97_11;
	wire [WIDTH*2-1+0:0] tmp00_97_12;
	wire [WIDTH*2-1+0:0] tmp00_97_13;
	wire [WIDTH*2-1+0:0] tmp00_97_14;
	wire [WIDTH*2-1+0:0] tmp00_97_15;
	wire [WIDTH*2-1+0:0] tmp00_97_16;
	wire [WIDTH*2-1+0:0] tmp00_97_17;
	wire [WIDTH*2-1+0:0] tmp00_97_18;
	wire [WIDTH*2-1+0:0] tmp00_97_19;
	wire [WIDTH*2-1+0:0] tmp00_97_20;
	wire [WIDTH*2-1+0:0] tmp00_97_21;
	wire [WIDTH*2-1+0:0] tmp00_97_22;
	wire [WIDTH*2-1+0:0] tmp00_97_23;
	wire [WIDTH*2-1+0:0] tmp00_97_24;
	wire [WIDTH*2-1+0:0] tmp00_97_25;
	wire [WIDTH*2-1+0:0] tmp00_97_26;
	wire [WIDTH*2-1+0:0] tmp00_97_27;
	wire [WIDTH*2-1+0:0] tmp00_97_28;
	wire [WIDTH*2-1+0:0] tmp00_97_29;
	wire [WIDTH*2-1+0:0] tmp00_97_30;
	wire [WIDTH*2-1+0:0] tmp00_97_31;
	wire [WIDTH*2-1+0:0] tmp00_97_32;
	wire [WIDTH*2-1+0:0] tmp00_97_33;
	wire [WIDTH*2-1+0:0] tmp00_97_34;
	wire [WIDTH*2-1+0:0] tmp00_97_35;
	wire [WIDTH*2-1+0:0] tmp00_97_36;
	wire [WIDTH*2-1+0:0] tmp00_97_37;
	wire [WIDTH*2-1+0:0] tmp00_97_38;
	wire [WIDTH*2-1+0:0] tmp00_97_39;
	wire [WIDTH*2-1+0:0] tmp00_97_40;
	wire [WIDTH*2-1+0:0] tmp00_97_41;
	wire [WIDTH*2-1+0:0] tmp00_97_42;
	wire [WIDTH*2-1+0:0] tmp00_97_43;
	wire [WIDTH*2-1+0:0] tmp00_97_44;
	wire [WIDTH*2-1+0:0] tmp00_97_45;
	wire [WIDTH*2-1+0:0] tmp00_97_46;
	wire [WIDTH*2-1+0:0] tmp00_97_47;
	wire [WIDTH*2-1+0:0] tmp00_97_48;
	wire [WIDTH*2-1+0:0] tmp00_97_49;
	wire [WIDTH*2-1+0:0] tmp00_97_50;
	wire [WIDTH*2-1+0:0] tmp00_97_51;
	wire [WIDTH*2-1+0:0] tmp00_97_52;
	wire [WIDTH*2-1+0:0] tmp00_97_53;
	wire [WIDTH*2-1+0:0] tmp00_97_54;
	wire [WIDTH*2-1+0:0] tmp00_97_55;
	wire [WIDTH*2-1+0:0] tmp00_97_56;
	wire [WIDTH*2-1+0:0] tmp00_97_57;
	wire [WIDTH*2-1+0:0] tmp00_97_58;
	wire [WIDTH*2-1+0:0] tmp00_97_59;
	wire [WIDTH*2-1+0:0] tmp00_97_60;
	wire [WIDTH*2-1+0:0] tmp00_97_61;
	wire [WIDTH*2-1+0:0] tmp00_97_62;
	wire [WIDTH*2-1+0:0] tmp00_97_63;
	wire [WIDTH*2-1+0:0] tmp00_97_64;
	wire [WIDTH*2-1+0:0] tmp00_97_65;
	wire [WIDTH*2-1+0:0] tmp00_97_66;
	wire [WIDTH*2-1+0:0] tmp00_97_67;
	wire [WIDTH*2-1+0:0] tmp00_97_68;
	wire [WIDTH*2-1+0:0] tmp00_97_69;
	wire [WIDTH*2-1+0:0] tmp00_97_70;
	wire [WIDTH*2-1+0:0] tmp00_97_71;
	wire [WIDTH*2-1+0:0] tmp00_97_72;
	wire [WIDTH*2-1+0:0] tmp00_97_73;
	wire [WIDTH*2-1+0:0] tmp00_97_74;
	wire [WIDTH*2-1+0:0] tmp00_97_75;
	wire [WIDTH*2-1+0:0] tmp00_97_76;
	wire [WIDTH*2-1+0:0] tmp00_97_77;
	wire [WIDTH*2-1+0:0] tmp00_97_78;
	wire [WIDTH*2-1+0:0] tmp00_97_79;
	wire [WIDTH*2-1+0:0] tmp00_97_80;
	wire [WIDTH*2-1+0:0] tmp00_97_81;
	wire [WIDTH*2-1+0:0] tmp00_97_82;
	wire [WIDTH*2-1+0:0] tmp00_97_83;
	wire [WIDTH*2-1+0:0] tmp00_98_0;
	wire [WIDTH*2-1+0:0] tmp00_98_1;
	wire [WIDTH*2-1+0:0] tmp00_98_2;
	wire [WIDTH*2-1+0:0] tmp00_98_3;
	wire [WIDTH*2-1+0:0] tmp00_98_4;
	wire [WIDTH*2-1+0:0] tmp00_98_5;
	wire [WIDTH*2-1+0:0] tmp00_98_6;
	wire [WIDTH*2-1+0:0] tmp00_98_7;
	wire [WIDTH*2-1+0:0] tmp00_98_8;
	wire [WIDTH*2-1+0:0] tmp00_98_9;
	wire [WIDTH*2-1+0:0] tmp00_98_10;
	wire [WIDTH*2-1+0:0] tmp00_98_11;
	wire [WIDTH*2-1+0:0] tmp00_98_12;
	wire [WIDTH*2-1+0:0] tmp00_98_13;
	wire [WIDTH*2-1+0:0] tmp00_98_14;
	wire [WIDTH*2-1+0:0] tmp00_98_15;
	wire [WIDTH*2-1+0:0] tmp00_98_16;
	wire [WIDTH*2-1+0:0] tmp00_98_17;
	wire [WIDTH*2-1+0:0] tmp00_98_18;
	wire [WIDTH*2-1+0:0] tmp00_98_19;
	wire [WIDTH*2-1+0:0] tmp00_98_20;
	wire [WIDTH*2-1+0:0] tmp00_98_21;
	wire [WIDTH*2-1+0:0] tmp00_98_22;
	wire [WIDTH*2-1+0:0] tmp00_98_23;
	wire [WIDTH*2-1+0:0] tmp00_98_24;
	wire [WIDTH*2-1+0:0] tmp00_98_25;
	wire [WIDTH*2-1+0:0] tmp00_98_26;
	wire [WIDTH*2-1+0:0] tmp00_98_27;
	wire [WIDTH*2-1+0:0] tmp00_98_28;
	wire [WIDTH*2-1+0:0] tmp00_98_29;
	wire [WIDTH*2-1+0:0] tmp00_98_30;
	wire [WIDTH*2-1+0:0] tmp00_98_31;
	wire [WIDTH*2-1+0:0] tmp00_98_32;
	wire [WIDTH*2-1+0:0] tmp00_98_33;
	wire [WIDTH*2-1+0:0] tmp00_98_34;
	wire [WIDTH*2-1+0:0] tmp00_98_35;
	wire [WIDTH*2-1+0:0] tmp00_98_36;
	wire [WIDTH*2-1+0:0] tmp00_98_37;
	wire [WIDTH*2-1+0:0] tmp00_98_38;
	wire [WIDTH*2-1+0:0] tmp00_98_39;
	wire [WIDTH*2-1+0:0] tmp00_98_40;
	wire [WIDTH*2-1+0:0] tmp00_98_41;
	wire [WIDTH*2-1+0:0] tmp00_98_42;
	wire [WIDTH*2-1+0:0] tmp00_98_43;
	wire [WIDTH*2-1+0:0] tmp00_98_44;
	wire [WIDTH*2-1+0:0] tmp00_98_45;
	wire [WIDTH*2-1+0:0] tmp00_98_46;
	wire [WIDTH*2-1+0:0] tmp00_98_47;
	wire [WIDTH*2-1+0:0] tmp00_98_48;
	wire [WIDTH*2-1+0:0] tmp00_98_49;
	wire [WIDTH*2-1+0:0] tmp00_98_50;
	wire [WIDTH*2-1+0:0] tmp00_98_51;
	wire [WIDTH*2-1+0:0] tmp00_98_52;
	wire [WIDTH*2-1+0:0] tmp00_98_53;
	wire [WIDTH*2-1+0:0] tmp00_98_54;
	wire [WIDTH*2-1+0:0] tmp00_98_55;
	wire [WIDTH*2-1+0:0] tmp00_98_56;
	wire [WIDTH*2-1+0:0] tmp00_98_57;
	wire [WIDTH*2-1+0:0] tmp00_98_58;
	wire [WIDTH*2-1+0:0] tmp00_98_59;
	wire [WIDTH*2-1+0:0] tmp00_98_60;
	wire [WIDTH*2-1+0:0] tmp00_98_61;
	wire [WIDTH*2-1+0:0] tmp00_98_62;
	wire [WIDTH*2-1+0:0] tmp00_98_63;
	wire [WIDTH*2-1+0:0] tmp00_98_64;
	wire [WIDTH*2-1+0:0] tmp00_98_65;
	wire [WIDTH*2-1+0:0] tmp00_98_66;
	wire [WIDTH*2-1+0:0] tmp00_98_67;
	wire [WIDTH*2-1+0:0] tmp00_98_68;
	wire [WIDTH*2-1+0:0] tmp00_98_69;
	wire [WIDTH*2-1+0:0] tmp00_98_70;
	wire [WIDTH*2-1+0:0] tmp00_98_71;
	wire [WIDTH*2-1+0:0] tmp00_98_72;
	wire [WIDTH*2-1+0:0] tmp00_98_73;
	wire [WIDTH*2-1+0:0] tmp00_98_74;
	wire [WIDTH*2-1+0:0] tmp00_98_75;
	wire [WIDTH*2-1+0:0] tmp00_98_76;
	wire [WIDTH*2-1+0:0] tmp00_98_77;
	wire [WIDTH*2-1+0:0] tmp00_98_78;
	wire [WIDTH*2-1+0:0] tmp00_98_79;
	wire [WIDTH*2-1+0:0] tmp00_98_80;
	wire [WIDTH*2-1+0:0] tmp00_98_81;
	wire [WIDTH*2-1+0:0] tmp00_98_82;
	wire [WIDTH*2-1+0:0] tmp00_98_83;
	wire [WIDTH*2-1+0:0] tmp00_99_0;
	wire [WIDTH*2-1+0:0] tmp00_99_1;
	wire [WIDTH*2-1+0:0] tmp00_99_2;
	wire [WIDTH*2-1+0:0] tmp00_99_3;
	wire [WIDTH*2-1+0:0] tmp00_99_4;
	wire [WIDTH*2-1+0:0] tmp00_99_5;
	wire [WIDTH*2-1+0:0] tmp00_99_6;
	wire [WIDTH*2-1+0:0] tmp00_99_7;
	wire [WIDTH*2-1+0:0] tmp00_99_8;
	wire [WIDTH*2-1+0:0] tmp00_99_9;
	wire [WIDTH*2-1+0:0] tmp00_99_10;
	wire [WIDTH*2-1+0:0] tmp00_99_11;
	wire [WIDTH*2-1+0:0] tmp00_99_12;
	wire [WIDTH*2-1+0:0] tmp00_99_13;
	wire [WIDTH*2-1+0:0] tmp00_99_14;
	wire [WIDTH*2-1+0:0] tmp00_99_15;
	wire [WIDTH*2-1+0:0] tmp00_99_16;
	wire [WIDTH*2-1+0:0] tmp00_99_17;
	wire [WIDTH*2-1+0:0] tmp00_99_18;
	wire [WIDTH*2-1+0:0] tmp00_99_19;
	wire [WIDTH*2-1+0:0] tmp00_99_20;
	wire [WIDTH*2-1+0:0] tmp00_99_21;
	wire [WIDTH*2-1+0:0] tmp00_99_22;
	wire [WIDTH*2-1+0:0] tmp00_99_23;
	wire [WIDTH*2-1+0:0] tmp00_99_24;
	wire [WIDTH*2-1+0:0] tmp00_99_25;
	wire [WIDTH*2-1+0:0] tmp00_99_26;
	wire [WIDTH*2-1+0:0] tmp00_99_27;
	wire [WIDTH*2-1+0:0] tmp00_99_28;
	wire [WIDTH*2-1+0:0] tmp00_99_29;
	wire [WIDTH*2-1+0:0] tmp00_99_30;
	wire [WIDTH*2-1+0:0] tmp00_99_31;
	wire [WIDTH*2-1+0:0] tmp00_99_32;
	wire [WIDTH*2-1+0:0] tmp00_99_33;
	wire [WIDTH*2-1+0:0] tmp00_99_34;
	wire [WIDTH*2-1+0:0] tmp00_99_35;
	wire [WIDTH*2-1+0:0] tmp00_99_36;
	wire [WIDTH*2-1+0:0] tmp00_99_37;
	wire [WIDTH*2-1+0:0] tmp00_99_38;
	wire [WIDTH*2-1+0:0] tmp00_99_39;
	wire [WIDTH*2-1+0:0] tmp00_99_40;
	wire [WIDTH*2-1+0:0] tmp00_99_41;
	wire [WIDTH*2-1+0:0] tmp00_99_42;
	wire [WIDTH*2-1+0:0] tmp00_99_43;
	wire [WIDTH*2-1+0:0] tmp00_99_44;
	wire [WIDTH*2-1+0:0] tmp00_99_45;
	wire [WIDTH*2-1+0:0] tmp00_99_46;
	wire [WIDTH*2-1+0:0] tmp00_99_47;
	wire [WIDTH*2-1+0:0] tmp00_99_48;
	wire [WIDTH*2-1+0:0] tmp00_99_49;
	wire [WIDTH*2-1+0:0] tmp00_99_50;
	wire [WIDTH*2-1+0:0] tmp00_99_51;
	wire [WIDTH*2-1+0:0] tmp00_99_52;
	wire [WIDTH*2-1+0:0] tmp00_99_53;
	wire [WIDTH*2-1+0:0] tmp00_99_54;
	wire [WIDTH*2-1+0:0] tmp00_99_55;
	wire [WIDTH*2-1+0:0] tmp00_99_56;
	wire [WIDTH*2-1+0:0] tmp00_99_57;
	wire [WIDTH*2-1+0:0] tmp00_99_58;
	wire [WIDTH*2-1+0:0] tmp00_99_59;
	wire [WIDTH*2-1+0:0] tmp00_99_60;
	wire [WIDTH*2-1+0:0] tmp00_99_61;
	wire [WIDTH*2-1+0:0] tmp00_99_62;
	wire [WIDTH*2-1+0:0] tmp00_99_63;
	wire [WIDTH*2-1+0:0] tmp00_99_64;
	wire [WIDTH*2-1+0:0] tmp00_99_65;
	wire [WIDTH*2-1+0:0] tmp00_99_66;
	wire [WIDTH*2-1+0:0] tmp00_99_67;
	wire [WIDTH*2-1+0:0] tmp00_99_68;
	wire [WIDTH*2-1+0:0] tmp00_99_69;
	wire [WIDTH*2-1+0:0] tmp00_99_70;
	wire [WIDTH*2-1+0:0] tmp00_99_71;
	wire [WIDTH*2-1+0:0] tmp00_99_72;
	wire [WIDTH*2-1+0:0] tmp00_99_73;
	wire [WIDTH*2-1+0:0] tmp00_99_74;
	wire [WIDTH*2-1+0:0] tmp00_99_75;
	wire [WIDTH*2-1+0:0] tmp00_99_76;
	wire [WIDTH*2-1+0:0] tmp00_99_77;
	wire [WIDTH*2-1+0:0] tmp00_99_78;
	wire [WIDTH*2-1+0:0] tmp00_99_79;
	wire [WIDTH*2-1+0:0] tmp00_99_80;
	wire [WIDTH*2-1+0:0] tmp00_99_81;
	wire [WIDTH*2-1+0:0] tmp00_99_82;
	wire [WIDTH*2-1+0:0] tmp00_99_83;
	wire [WIDTH*2-1+0:0] tmp00_100_0;
	wire [WIDTH*2-1+0:0] tmp00_100_1;
	wire [WIDTH*2-1+0:0] tmp00_100_2;
	wire [WIDTH*2-1+0:0] tmp00_100_3;
	wire [WIDTH*2-1+0:0] tmp00_100_4;
	wire [WIDTH*2-1+0:0] tmp00_100_5;
	wire [WIDTH*2-1+0:0] tmp00_100_6;
	wire [WIDTH*2-1+0:0] tmp00_100_7;
	wire [WIDTH*2-1+0:0] tmp00_100_8;
	wire [WIDTH*2-1+0:0] tmp00_100_9;
	wire [WIDTH*2-1+0:0] tmp00_100_10;
	wire [WIDTH*2-1+0:0] tmp00_100_11;
	wire [WIDTH*2-1+0:0] tmp00_100_12;
	wire [WIDTH*2-1+0:0] tmp00_100_13;
	wire [WIDTH*2-1+0:0] tmp00_100_14;
	wire [WIDTH*2-1+0:0] tmp00_100_15;
	wire [WIDTH*2-1+0:0] tmp00_100_16;
	wire [WIDTH*2-1+0:0] tmp00_100_17;
	wire [WIDTH*2-1+0:0] tmp00_100_18;
	wire [WIDTH*2-1+0:0] tmp00_100_19;
	wire [WIDTH*2-1+0:0] tmp00_100_20;
	wire [WIDTH*2-1+0:0] tmp00_100_21;
	wire [WIDTH*2-1+0:0] tmp00_100_22;
	wire [WIDTH*2-1+0:0] tmp00_100_23;
	wire [WIDTH*2-1+0:0] tmp00_100_24;
	wire [WIDTH*2-1+0:0] tmp00_100_25;
	wire [WIDTH*2-1+0:0] tmp00_100_26;
	wire [WIDTH*2-1+0:0] tmp00_100_27;
	wire [WIDTH*2-1+0:0] tmp00_100_28;
	wire [WIDTH*2-1+0:0] tmp00_100_29;
	wire [WIDTH*2-1+0:0] tmp00_100_30;
	wire [WIDTH*2-1+0:0] tmp00_100_31;
	wire [WIDTH*2-1+0:0] tmp00_100_32;
	wire [WIDTH*2-1+0:0] tmp00_100_33;
	wire [WIDTH*2-1+0:0] tmp00_100_34;
	wire [WIDTH*2-1+0:0] tmp00_100_35;
	wire [WIDTH*2-1+0:0] tmp00_100_36;
	wire [WIDTH*2-1+0:0] tmp00_100_37;
	wire [WIDTH*2-1+0:0] tmp00_100_38;
	wire [WIDTH*2-1+0:0] tmp00_100_39;
	wire [WIDTH*2-1+0:0] tmp00_100_40;
	wire [WIDTH*2-1+0:0] tmp00_100_41;
	wire [WIDTH*2-1+0:0] tmp00_100_42;
	wire [WIDTH*2-1+0:0] tmp00_100_43;
	wire [WIDTH*2-1+0:0] tmp00_100_44;
	wire [WIDTH*2-1+0:0] tmp00_100_45;
	wire [WIDTH*2-1+0:0] tmp00_100_46;
	wire [WIDTH*2-1+0:0] tmp00_100_47;
	wire [WIDTH*2-1+0:0] tmp00_100_48;
	wire [WIDTH*2-1+0:0] tmp00_100_49;
	wire [WIDTH*2-1+0:0] tmp00_100_50;
	wire [WIDTH*2-1+0:0] tmp00_100_51;
	wire [WIDTH*2-1+0:0] tmp00_100_52;
	wire [WIDTH*2-1+0:0] tmp00_100_53;
	wire [WIDTH*2-1+0:0] tmp00_100_54;
	wire [WIDTH*2-1+0:0] tmp00_100_55;
	wire [WIDTH*2-1+0:0] tmp00_100_56;
	wire [WIDTH*2-1+0:0] tmp00_100_57;
	wire [WIDTH*2-1+0:0] tmp00_100_58;
	wire [WIDTH*2-1+0:0] tmp00_100_59;
	wire [WIDTH*2-1+0:0] tmp00_100_60;
	wire [WIDTH*2-1+0:0] tmp00_100_61;
	wire [WIDTH*2-1+0:0] tmp00_100_62;
	wire [WIDTH*2-1+0:0] tmp00_100_63;
	wire [WIDTH*2-1+0:0] tmp00_100_64;
	wire [WIDTH*2-1+0:0] tmp00_100_65;
	wire [WIDTH*2-1+0:0] tmp00_100_66;
	wire [WIDTH*2-1+0:0] tmp00_100_67;
	wire [WIDTH*2-1+0:0] tmp00_100_68;
	wire [WIDTH*2-1+0:0] tmp00_100_69;
	wire [WIDTH*2-1+0:0] tmp00_100_70;
	wire [WIDTH*2-1+0:0] tmp00_100_71;
	wire [WIDTH*2-1+0:0] tmp00_100_72;
	wire [WIDTH*2-1+0:0] tmp00_100_73;
	wire [WIDTH*2-1+0:0] tmp00_100_74;
	wire [WIDTH*2-1+0:0] tmp00_100_75;
	wire [WIDTH*2-1+0:0] tmp00_100_76;
	wire [WIDTH*2-1+0:0] tmp00_100_77;
	wire [WIDTH*2-1+0:0] tmp00_100_78;
	wire [WIDTH*2-1+0:0] tmp00_100_79;
	wire [WIDTH*2-1+0:0] tmp00_100_80;
	wire [WIDTH*2-1+0:0] tmp00_100_81;
	wire [WIDTH*2-1+0:0] tmp00_100_82;
	wire [WIDTH*2-1+0:0] tmp00_100_83;
	wire [WIDTH*2-1+0:0] tmp00_101_0;
	wire [WIDTH*2-1+0:0] tmp00_101_1;
	wire [WIDTH*2-1+0:0] tmp00_101_2;
	wire [WIDTH*2-1+0:0] tmp00_101_3;
	wire [WIDTH*2-1+0:0] tmp00_101_4;
	wire [WIDTH*2-1+0:0] tmp00_101_5;
	wire [WIDTH*2-1+0:0] tmp00_101_6;
	wire [WIDTH*2-1+0:0] tmp00_101_7;
	wire [WIDTH*2-1+0:0] tmp00_101_8;
	wire [WIDTH*2-1+0:0] tmp00_101_9;
	wire [WIDTH*2-1+0:0] tmp00_101_10;
	wire [WIDTH*2-1+0:0] tmp00_101_11;
	wire [WIDTH*2-1+0:0] tmp00_101_12;
	wire [WIDTH*2-1+0:0] tmp00_101_13;
	wire [WIDTH*2-1+0:0] tmp00_101_14;
	wire [WIDTH*2-1+0:0] tmp00_101_15;
	wire [WIDTH*2-1+0:0] tmp00_101_16;
	wire [WIDTH*2-1+0:0] tmp00_101_17;
	wire [WIDTH*2-1+0:0] tmp00_101_18;
	wire [WIDTH*2-1+0:0] tmp00_101_19;
	wire [WIDTH*2-1+0:0] tmp00_101_20;
	wire [WIDTH*2-1+0:0] tmp00_101_21;
	wire [WIDTH*2-1+0:0] tmp00_101_22;
	wire [WIDTH*2-1+0:0] tmp00_101_23;
	wire [WIDTH*2-1+0:0] tmp00_101_24;
	wire [WIDTH*2-1+0:0] tmp00_101_25;
	wire [WIDTH*2-1+0:0] tmp00_101_26;
	wire [WIDTH*2-1+0:0] tmp00_101_27;
	wire [WIDTH*2-1+0:0] tmp00_101_28;
	wire [WIDTH*2-1+0:0] tmp00_101_29;
	wire [WIDTH*2-1+0:0] tmp00_101_30;
	wire [WIDTH*2-1+0:0] tmp00_101_31;
	wire [WIDTH*2-1+0:0] tmp00_101_32;
	wire [WIDTH*2-1+0:0] tmp00_101_33;
	wire [WIDTH*2-1+0:0] tmp00_101_34;
	wire [WIDTH*2-1+0:0] tmp00_101_35;
	wire [WIDTH*2-1+0:0] tmp00_101_36;
	wire [WIDTH*2-1+0:0] tmp00_101_37;
	wire [WIDTH*2-1+0:0] tmp00_101_38;
	wire [WIDTH*2-1+0:0] tmp00_101_39;
	wire [WIDTH*2-1+0:0] tmp00_101_40;
	wire [WIDTH*2-1+0:0] tmp00_101_41;
	wire [WIDTH*2-1+0:0] tmp00_101_42;
	wire [WIDTH*2-1+0:0] tmp00_101_43;
	wire [WIDTH*2-1+0:0] tmp00_101_44;
	wire [WIDTH*2-1+0:0] tmp00_101_45;
	wire [WIDTH*2-1+0:0] tmp00_101_46;
	wire [WIDTH*2-1+0:0] tmp00_101_47;
	wire [WIDTH*2-1+0:0] tmp00_101_48;
	wire [WIDTH*2-1+0:0] tmp00_101_49;
	wire [WIDTH*2-1+0:0] tmp00_101_50;
	wire [WIDTH*2-1+0:0] tmp00_101_51;
	wire [WIDTH*2-1+0:0] tmp00_101_52;
	wire [WIDTH*2-1+0:0] tmp00_101_53;
	wire [WIDTH*2-1+0:0] tmp00_101_54;
	wire [WIDTH*2-1+0:0] tmp00_101_55;
	wire [WIDTH*2-1+0:0] tmp00_101_56;
	wire [WIDTH*2-1+0:0] tmp00_101_57;
	wire [WIDTH*2-1+0:0] tmp00_101_58;
	wire [WIDTH*2-1+0:0] tmp00_101_59;
	wire [WIDTH*2-1+0:0] tmp00_101_60;
	wire [WIDTH*2-1+0:0] tmp00_101_61;
	wire [WIDTH*2-1+0:0] tmp00_101_62;
	wire [WIDTH*2-1+0:0] tmp00_101_63;
	wire [WIDTH*2-1+0:0] tmp00_101_64;
	wire [WIDTH*2-1+0:0] tmp00_101_65;
	wire [WIDTH*2-1+0:0] tmp00_101_66;
	wire [WIDTH*2-1+0:0] tmp00_101_67;
	wire [WIDTH*2-1+0:0] tmp00_101_68;
	wire [WIDTH*2-1+0:0] tmp00_101_69;
	wire [WIDTH*2-1+0:0] tmp00_101_70;
	wire [WIDTH*2-1+0:0] tmp00_101_71;
	wire [WIDTH*2-1+0:0] tmp00_101_72;
	wire [WIDTH*2-1+0:0] tmp00_101_73;
	wire [WIDTH*2-1+0:0] tmp00_101_74;
	wire [WIDTH*2-1+0:0] tmp00_101_75;
	wire [WIDTH*2-1+0:0] tmp00_101_76;
	wire [WIDTH*2-1+0:0] tmp00_101_77;
	wire [WIDTH*2-1+0:0] tmp00_101_78;
	wire [WIDTH*2-1+0:0] tmp00_101_79;
	wire [WIDTH*2-1+0:0] tmp00_101_80;
	wire [WIDTH*2-1+0:0] tmp00_101_81;
	wire [WIDTH*2-1+0:0] tmp00_101_82;
	wire [WIDTH*2-1+0:0] tmp00_101_83;
	wire [WIDTH*2-1+0:0] tmp00_102_0;
	wire [WIDTH*2-1+0:0] tmp00_102_1;
	wire [WIDTH*2-1+0:0] tmp00_102_2;
	wire [WIDTH*2-1+0:0] tmp00_102_3;
	wire [WIDTH*2-1+0:0] tmp00_102_4;
	wire [WIDTH*2-1+0:0] tmp00_102_5;
	wire [WIDTH*2-1+0:0] tmp00_102_6;
	wire [WIDTH*2-1+0:0] tmp00_102_7;
	wire [WIDTH*2-1+0:0] tmp00_102_8;
	wire [WIDTH*2-1+0:0] tmp00_102_9;
	wire [WIDTH*2-1+0:0] tmp00_102_10;
	wire [WIDTH*2-1+0:0] tmp00_102_11;
	wire [WIDTH*2-1+0:0] tmp00_102_12;
	wire [WIDTH*2-1+0:0] tmp00_102_13;
	wire [WIDTH*2-1+0:0] tmp00_102_14;
	wire [WIDTH*2-1+0:0] tmp00_102_15;
	wire [WIDTH*2-1+0:0] tmp00_102_16;
	wire [WIDTH*2-1+0:0] tmp00_102_17;
	wire [WIDTH*2-1+0:0] tmp00_102_18;
	wire [WIDTH*2-1+0:0] tmp00_102_19;
	wire [WIDTH*2-1+0:0] tmp00_102_20;
	wire [WIDTH*2-1+0:0] tmp00_102_21;
	wire [WIDTH*2-1+0:0] tmp00_102_22;
	wire [WIDTH*2-1+0:0] tmp00_102_23;
	wire [WIDTH*2-1+0:0] tmp00_102_24;
	wire [WIDTH*2-1+0:0] tmp00_102_25;
	wire [WIDTH*2-1+0:0] tmp00_102_26;
	wire [WIDTH*2-1+0:0] tmp00_102_27;
	wire [WIDTH*2-1+0:0] tmp00_102_28;
	wire [WIDTH*2-1+0:0] tmp00_102_29;
	wire [WIDTH*2-1+0:0] tmp00_102_30;
	wire [WIDTH*2-1+0:0] tmp00_102_31;
	wire [WIDTH*2-1+0:0] tmp00_102_32;
	wire [WIDTH*2-1+0:0] tmp00_102_33;
	wire [WIDTH*2-1+0:0] tmp00_102_34;
	wire [WIDTH*2-1+0:0] tmp00_102_35;
	wire [WIDTH*2-1+0:0] tmp00_102_36;
	wire [WIDTH*2-1+0:0] tmp00_102_37;
	wire [WIDTH*2-1+0:0] tmp00_102_38;
	wire [WIDTH*2-1+0:0] tmp00_102_39;
	wire [WIDTH*2-1+0:0] tmp00_102_40;
	wire [WIDTH*2-1+0:0] tmp00_102_41;
	wire [WIDTH*2-1+0:0] tmp00_102_42;
	wire [WIDTH*2-1+0:0] tmp00_102_43;
	wire [WIDTH*2-1+0:0] tmp00_102_44;
	wire [WIDTH*2-1+0:0] tmp00_102_45;
	wire [WIDTH*2-1+0:0] tmp00_102_46;
	wire [WIDTH*2-1+0:0] tmp00_102_47;
	wire [WIDTH*2-1+0:0] tmp00_102_48;
	wire [WIDTH*2-1+0:0] tmp00_102_49;
	wire [WIDTH*2-1+0:0] tmp00_102_50;
	wire [WIDTH*2-1+0:0] tmp00_102_51;
	wire [WIDTH*2-1+0:0] tmp00_102_52;
	wire [WIDTH*2-1+0:0] tmp00_102_53;
	wire [WIDTH*2-1+0:0] tmp00_102_54;
	wire [WIDTH*2-1+0:0] tmp00_102_55;
	wire [WIDTH*2-1+0:0] tmp00_102_56;
	wire [WIDTH*2-1+0:0] tmp00_102_57;
	wire [WIDTH*2-1+0:0] tmp00_102_58;
	wire [WIDTH*2-1+0:0] tmp00_102_59;
	wire [WIDTH*2-1+0:0] tmp00_102_60;
	wire [WIDTH*2-1+0:0] tmp00_102_61;
	wire [WIDTH*2-1+0:0] tmp00_102_62;
	wire [WIDTH*2-1+0:0] tmp00_102_63;
	wire [WIDTH*2-1+0:0] tmp00_102_64;
	wire [WIDTH*2-1+0:0] tmp00_102_65;
	wire [WIDTH*2-1+0:0] tmp00_102_66;
	wire [WIDTH*2-1+0:0] tmp00_102_67;
	wire [WIDTH*2-1+0:0] tmp00_102_68;
	wire [WIDTH*2-1+0:0] tmp00_102_69;
	wire [WIDTH*2-1+0:0] tmp00_102_70;
	wire [WIDTH*2-1+0:0] tmp00_102_71;
	wire [WIDTH*2-1+0:0] tmp00_102_72;
	wire [WIDTH*2-1+0:0] tmp00_102_73;
	wire [WIDTH*2-1+0:0] tmp00_102_74;
	wire [WIDTH*2-1+0:0] tmp00_102_75;
	wire [WIDTH*2-1+0:0] tmp00_102_76;
	wire [WIDTH*2-1+0:0] tmp00_102_77;
	wire [WIDTH*2-1+0:0] tmp00_102_78;
	wire [WIDTH*2-1+0:0] tmp00_102_79;
	wire [WIDTH*2-1+0:0] tmp00_102_80;
	wire [WIDTH*2-1+0:0] tmp00_102_81;
	wire [WIDTH*2-1+0:0] tmp00_102_82;
	wire [WIDTH*2-1+0:0] tmp00_102_83;
	wire [WIDTH*2-1+0:0] tmp00_103_0;
	wire [WIDTH*2-1+0:0] tmp00_103_1;
	wire [WIDTH*2-1+0:0] tmp00_103_2;
	wire [WIDTH*2-1+0:0] tmp00_103_3;
	wire [WIDTH*2-1+0:0] tmp00_103_4;
	wire [WIDTH*2-1+0:0] tmp00_103_5;
	wire [WIDTH*2-1+0:0] tmp00_103_6;
	wire [WIDTH*2-1+0:0] tmp00_103_7;
	wire [WIDTH*2-1+0:0] tmp00_103_8;
	wire [WIDTH*2-1+0:0] tmp00_103_9;
	wire [WIDTH*2-1+0:0] tmp00_103_10;
	wire [WIDTH*2-1+0:0] tmp00_103_11;
	wire [WIDTH*2-1+0:0] tmp00_103_12;
	wire [WIDTH*2-1+0:0] tmp00_103_13;
	wire [WIDTH*2-1+0:0] tmp00_103_14;
	wire [WIDTH*2-1+0:0] tmp00_103_15;
	wire [WIDTH*2-1+0:0] tmp00_103_16;
	wire [WIDTH*2-1+0:0] tmp00_103_17;
	wire [WIDTH*2-1+0:0] tmp00_103_18;
	wire [WIDTH*2-1+0:0] tmp00_103_19;
	wire [WIDTH*2-1+0:0] tmp00_103_20;
	wire [WIDTH*2-1+0:0] tmp00_103_21;
	wire [WIDTH*2-1+0:0] tmp00_103_22;
	wire [WIDTH*2-1+0:0] tmp00_103_23;
	wire [WIDTH*2-1+0:0] tmp00_103_24;
	wire [WIDTH*2-1+0:0] tmp00_103_25;
	wire [WIDTH*2-1+0:0] tmp00_103_26;
	wire [WIDTH*2-1+0:0] tmp00_103_27;
	wire [WIDTH*2-1+0:0] tmp00_103_28;
	wire [WIDTH*2-1+0:0] tmp00_103_29;
	wire [WIDTH*2-1+0:0] tmp00_103_30;
	wire [WIDTH*2-1+0:0] tmp00_103_31;
	wire [WIDTH*2-1+0:0] tmp00_103_32;
	wire [WIDTH*2-1+0:0] tmp00_103_33;
	wire [WIDTH*2-1+0:0] tmp00_103_34;
	wire [WIDTH*2-1+0:0] tmp00_103_35;
	wire [WIDTH*2-1+0:0] tmp00_103_36;
	wire [WIDTH*2-1+0:0] tmp00_103_37;
	wire [WIDTH*2-1+0:0] tmp00_103_38;
	wire [WIDTH*2-1+0:0] tmp00_103_39;
	wire [WIDTH*2-1+0:0] tmp00_103_40;
	wire [WIDTH*2-1+0:0] tmp00_103_41;
	wire [WIDTH*2-1+0:0] tmp00_103_42;
	wire [WIDTH*2-1+0:0] tmp00_103_43;
	wire [WIDTH*2-1+0:0] tmp00_103_44;
	wire [WIDTH*2-1+0:0] tmp00_103_45;
	wire [WIDTH*2-1+0:0] tmp00_103_46;
	wire [WIDTH*2-1+0:0] tmp00_103_47;
	wire [WIDTH*2-1+0:0] tmp00_103_48;
	wire [WIDTH*2-1+0:0] tmp00_103_49;
	wire [WIDTH*2-1+0:0] tmp00_103_50;
	wire [WIDTH*2-1+0:0] tmp00_103_51;
	wire [WIDTH*2-1+0:0] tmp00_103_52;
	wire [WIDTH*2-1+0:0] tmp00_103_53;
	wire [WIDTH*2-1+0:0] tmp00_103_54;
	wire [WIDTH*2-1+0:0] tmp00_103_55;
	wire [WIDTH*2-1+0:0] tmp00_103_56;
	wire [WIDTH*2-1+0:0] tmp00_103_57;
	wire [WIDTH*2-1+0:0] tmp00_103_58;
	wire [WIDTH*2-1+0:0] tmp00_103_59;
	wire [WIDTH*2-1+0:0] tmp00_103_60;
	wire [WIDTH*2-1+0:0] tmp00_103_61;
	wire [WIDTH*2-1+0:0] tmp00_103_62;
	wire [WIDTH*2-1+0:0] tmp00_103_63;
	wire [WIDTH*2-1+0:0] tmp00_103_64;
	wire [WIDTH*2-1+0:0] tmp00_103_65;
	wire [WIDTH*2-1+0:0] tmp00_103_66;
	wire [WIDTH*2-1+0:0] tmp00_103_67;
	wire [WIDTH*2-1+0:0] tmp00_103_68;
	wire [WIDTH*2-1+0:0] tmp00_103_69;
	wire [WIDTH*2-1+0:0] tmp00_103_70;
	wire [WIDTH*2-1+0:0] tmp00_103_71;
	wire [WIDTH*2-1+0:0] tmp00_103_72;
	wire [WIDTH*2-1+0:0] tmp00_103_73;
	wire [WIDTH*2-1+0:0] tmp00_103_74;
	wire [WIDTH*2-1+0:0] tmp00_103_75;
	wire [WIDTH*2-1+0:0] tmp00_103_76;
	wire [WIDTH*2-1+0:0] tmp00_103_77;
	wire [WIDTH*2-1+0:0] tmp00_103_78;
	wire [WIDTH*2-1+0:0] tmp00_103_79;
	wire [WIDTH*2-1+0:0] tmp00_103_80;
	wire [WIDTH*2-1+0:0] tmp00_103_81;
	wire [WIDTH*2-1+0:0] tmp00_103_82;
	wire [WIDTH*2-1+0:0] tmp00_103_83;
	wire [WIDTH*2-1+0:0] tmp00_104_0;
	wire [WIDTH*2-1+0:0] tmp00_104_1;
	wire [WIDTH*2-1+0:0] tmp00_104_2;
	wire [WIDTH*2-1+0:0] tmp00_104_3;
	wire [WIDTH*2-1+0:0] tmp00_104_4;
	wire [WIDTH*2-1+0:0] tmp00_104_5;
	wire [WIDTH*2-1+0:0] tmp00_104_6;
	wire [WIDTH*2-1+0:0] tmp00_104_7;
	wire [WIDTH*2-1+0:0] tmp00_104_8;
	wire [WIDTH*2-1+0:0] tmp00_104_9;
	wire [WIDTH*2-1+0:0] tmp00_104_10;
	wire [WIDTH*2-1+0:0] tmp00_104_11;
	wire [WIDTH*2-1+0:0] tmp00_104_12;
	wire [WIDTH*2-1+0:0] tmp00_104_13;
	wire [WIDTH*2-1+0:0] tmp00_104_14;
	wire [WIDTH*2-1+0:0] tmp00_104_15;
	wire [WIDTH*2-1+0:0] tmp00_104_16;
	wire [WIDTH*2-1+0:0] tmp00_104_17;
	wire [WIDTH*2-1+0:0] tmp00_104_18;
	wire [WIDTH*2-1+0:0] tmp00_104_19;
	wire [WIDTH*2-1+0:0] tmp00_104_20;
	wire [WIDTH*2-1+0:0] tmp00_104_21;
	wire [WIDTH*2-1+0:0] tmp00_104_22;
	wire [WIDTH*2-1+0:0] tmp00_104_23;
	wire [WIDTH*2-1+0:0] tmp00_104_24;
	wire [WIDTH*2-1+0:0] tmp00_104_25;
	wire [WIDTH*2-1+0:0] tmp00_104_26;
	wire [WIDTH*2-1+0:0] tmp00_104_27;
	wire [WIDTH*2-1+0:0] tmp00_104_28;
	wire [WIDTH*2-1+0:0] tmp00_104_29;
	wire [WIDTH*2-1+0:0] tmp00_104_30;
	wire [WIDTH*2-1+0:0] tmp00_104_31;
	wire [WIDTH*2-1+0:0] tmp00_104_32;
	wire [WIDTH*2-1+0:0] tmp00_104_33;
	wire [WIDTH*2-1+0:0] tmp00_104_34;
	wire [WIDTH*2-1+0:0] tmp00_104_35;
	wire [WIDTH*2-1+0:0] tmp00_104_36;
	wire [WIDTH*2-1+0:0] tmp00_104_37;
	wire [WIDTH*2-1+0:0] tmp00_104_38;
	wire [WIDTH*2-1+0:0] tmp00_104_39;
	wire [WIDTH*2-1+0:0] tmp00_104_40;
	wire [WIDTH*2-1+0:0] tmp00_104_41;
	wire [WIDTH*2-1+0:0] tmp00_104_42;
	wire [WIDTH*2-1+0:0] tmp00_104_43;
	wire [WIDTH*2-1+0:0] tmp00_104_44;
	wire [WIDTH*2-1+0:0] tmp00_104_45;
	wire [WIDTH*2-1+0:0] tmp00_104_46;
	wire [WIDTH*2-1+0:0] tmp00_104_47;
	wire [WIDTH*2-1+0:0] tmp00_104_48;
	wire [WIDTH*2-1+0:0] tmp00_104_49;
	wire [WIDTH*2-1+0:0] tmp00_104_50;
	wire [WIDTH*2-1+0:0] tmp00_104_51;
	wire [WIDTH*2-1+0:0] tmp00_104_52;
	wire [WIDTH*2-1+0:0] tmp00_104_53;
	wire [WIDTH*2-1+0:0] tmp00_104_54;
	wire [WIDTH*2-1+0:0] tmp00_104_55;
	wire [WIDTH*2-1+0:0] tmp00_104_56;
	wire [WIDTH*2-1+0:0] tmp00_104_57;
	wire [WIDTH*2-1+0:0] tmp00_104_58;
	wire [WIDTH*2-1+0:0] tmp00_104_59;
	wire [WIDTH*2-1+0:0] tmp00_104_60;
	wire [WIDTH*2-1+0:0] tmp00_104_61;
	wire [WIDTH*2-1+0:0] tmp00_104_62;
	wire [WIDTH*2-1+0:0] tmp00_104_63;
	wire [WIDTH*2-1+0:0] tmp00_104_64;
	wire [WIDTH*2-1+0:0] tmp00_104_65;
	wire [WIDTH*2-1+0:0] tmp00_104_66;
	wire [WIDTH*2-1+0:0] tmp00_104_67;
	wire [WIDTH*2-1+0:0] tmp00_104_68;
	wire [WIDTH*2-1+0:0] tmp00_104_69;
	wire [WIDTH*2-1+0:0] tmp00_104_70;
	wire [WIDTH*2-1+0:0] tmp00_104_71;
	wire [WIDTH*2-1+0:0] tmp00_104_72;
	wire [WIDTH*2-1+0:0] tmp00_104_73;
	wire [WIDTH*2-1+0:0] tmp00_104_74;
	wire [WIDTH*2-1+0:0] tmp00_104_75;
	wire [WIDTH*2-1+0:0] tmp00_104_76;
	wire [WIDTH*2-1+0:0] tmp00_104_77;
	wire [WIDTH*2-1+0:0] tmp00_104_78;
	wire [WIDTH*2-1+0:0] tmp00_104_79;
	wire [WIDTH*2-1+0:0] tmp00_104_80;
	wire [WIDTH*2-1+0:0] tmp00_104_81;
	wire [WIDTH*2-1+0:0] tmp00_104_82;
	wire [WIDTH*2-1+0:0] tmp00_104_83;
	wire [WIDTH*2-1+0:0] tmp00_105_0;
	wire [WIDTH*2-1+0:0] tmp00_105_1;
	wire [WIDTH*2-1+0:0] tmp00_105_2;
	wire [WIDTH*2-1+0:0] tmp00_105_3;
	wire [WIDTH*2-1+0:0] tmp00_105_4;
	wire [WIDTH*2-1+0:0] tmp00_105_5;
	wire [WIDTH*2-1+0:0] tmp00_105_6;
	wire [WIDTH*2-1+0:0] tmp00_105_7;
	wire [WIDTH*2-1+0:0] tmp00_105_8;
	wire [WIDTH*2-1+0:0] tmp00_105_9;
	wire [WIDTH*2-1+0:0] tmp00_105_10;
	wire [WIDTH*2-1+0:0] tmp00_105_11;
	wire [WIDTH*2-1+0:0] tmp00_105_12;
	wire [WIDTH*2-1+0:0] tmp00_105_13;
	wire [WIDTH*2-1+0:0] tmp00_105_14;
	wire [WIDTH*2-1+0:0] tmp00_105_15;
	wire [WIDTH*2-1+0:0] tmp00_105_16;
	wire [WIDTH*2-1+0:0] tmp00_105_17;
	wire [WIDTH*2-1+0:0] tmp00_105_18;
	wire [WIDTH*2-1+0:0] tmp00_105_19;
	wire [WIDTH*2-1+0:0] tmp00_105_20;
	wire [WIDTH*2-1+0:0] tmp00_105_21;
	wire [WIDTH*2-1+0:0] tmp00_105_22;
	wire [WIDTH*2-1+0:0] tmp00_105_23;
	wire [WIDTH*2-1+0:0] tmp00_105_24;
	wire [WIDTH*2-1+0:0] tmp00_105_25;
	wire [WIDTH*2-1+0:0] tmp00_105_26;
	wire [WIDTH*2-1+0:0] tmp00_105_27;
	wire [WIDTH*2-1+0:0] tmp00_105_28;
	wire [WIDTH*2-1+0:0] tmp00_105_29;
	wire [WIDTH*2-1+0:0] tmp00_105_30;
	wire [WIDTH*2-1+0:0] tmp00_105_31;
	wire [WIDTH*2-1+0:0] tmp00_105_32;
	wire [WIDTH*2-1+0:0] tmp00_105_33;
	wire [WIDTH*2-1+0:0] tmp00_105_34;
	wire [WIDTH*2-1+0:0] tmp00_105_35;
	wire [WIDTH*2-1+0:0] tmp00_105_36;
	wire [WIDTH*2-1+0:0] tmp00_105_37;
	wire [WIDTH*2-1+0:0] tmp00_105_38;
	wire [WIDTH*2-1+0:0] tmp00_105_39;
	wire [WIDTH*2-1+0:0] tmp00_105_40;
	wire [WIDTH*2-1+0:0] tmp00_105_41;
	wire [WIDTH*2-1+0:0] tmp00_105_42;
	wire [WIDTH*2-1+0:0] tmp00_105_43;
	wire [WIDTH*2-1+0:0] tmp00_105_44;
	wire [WIDTH*2-1+0:0] tmp00_105_45;
	wire [WIDTH*2-1+0:0] tmp00_105_46;
	wire [WIDTH*2-1+0:0] tmp00_105_47;
	wire [WIDTH*2-1+0:0] tmp00_105_48;
	wire [WIDTH*2-1+0:0] tmp00_105_49;
	wire [WIDTH*2-1+0:0] tmp00_105_50;
	wire [WIDTH*2-1+0:0] tmp00_105_51;
	wire [WIDTH*2-1+0:0] tmp00_105_52;
	wire [WIDTH*2-1+0:0] tmp00_105_53;
	wire [WIDTH*2-1+0:0] tmp00_105_54;
	wire [WIDTH*2-1+0:0] tmp00_105_55;
	wire [WIDTH*2-1+0:0] tmp00_105_56;
	wire [WIDTH*2-1+0:0] tmp00_105_57;
	wire [WIDTH*2-1+0:0] tmp00_105_58;
	wire [WIDTH*2-1+0:0] tmp00_105_59;
	wire [WIDTH*2-1+0:0] tmp00_105_60;
	wire [WIDTH*2-1+0:0] tmp00_105_61;
	wire [WIDTH*2-1+0:0] tmp00_105_62;
	wire [WIDTH*2-1+0:0] tmp00_105_63;
	wire [WIDTH*2-1+0:0] tmp00_105_64;
	wire [WIDTH*2-1+0:0] tmp00_105_65;
	wire [WIDTH*2-1+0:0] tmp00_105_66;
	wire [WIDTH*2-1+0:0] tmp00_105_67;
	wire [WIDTH*2-1+0:0] tmp00_105_68;
	wire [WIDTH*2-1+0:0] tmp00_105_69;
	wire [WIDTH*2-1+0:0] tmp00_105_70;
	wire [WIDTH*2-1+0:0] tmp00_105_71;
	wire [WIDTH*2-1+0:0] tmp00_105_72;
	wire [WIDTH*2-1+0:0] tmp00_105_73;
	wire [WIDTH*2-1+0:0] tmp00_105_74;
	wire [WIDTH*2-1+0:0] tmp00_105_75;
	wire [WIDTH*2-1+0:0] tmp00_105_76;
	wire [WIDTH*2-1+0:0] tmp00_105_77;
	wire [WIDTH*2-1+0:0] tmp00_105_78;
	wire [WIDTH*2-1+0:0] tmp00_105_79;
	wire [WIDTH*2-1+0:0] tmp00_105_80;
	wire [WIDTH*2-1+0:0] tmp00_105_81;
	wire [WIDTH*2-1+0:0] tmp00_105_82;
	wire [WIDTH*2-1+0:0] tmp00_105_83;
	wire [WIDTH*2-1+0:0] tmp00_106_0;
	wire [WIDTH*2-1+0:0] tmp00_106_1;
	wire [WIDTH*2-1+0:0] tmp00_106_2;
	wire [WIDTH*2-1+0:0] tmp00_106_3;
	wire [WIDTH*2-1+0:0] tmp00_106_4;
	wire [WIDTH*2-1+0:0] tmp00_106_5;
	wire [WIDTH*2-1+0:0] tmp00_106_6;
	wire [WIDTH*2-1+0:0] tmp00_106_7;
	wire [WIDTH*2-1+0:0] tmp00_106_8;
	wire [WIDTH*2-1+0:0] tmp00_106_9;
	wire [WIDTH*2-1+0:0] tmp00_106_10;
	wire [WIDTH*2-1+0:0] tmp00_106_11;
	wire [WIDTH*2-1+0:0] tmp00_106_12;
	wire [WIDTH*2-1+0:0] tmp00_106_13;
	wire [WIDTH*2-1+0:0] tmp00_106_14;
	wire [WIDTH*2-1+0:0] tmp00_106_15;
	wire [WIDTH*2-1+0:0] tmp00_106_16;
	wire [WIDTH*2-1+0:0] tmp00_106_17;
	wire [WIDTH*2-1+0:0] tmp00_106_18;
	wire [WIDTH*2-1+0:0] tmp00_106_19;
	wire [WIDTH*2-1+0:0] tmp00_106_20;
	wire [WIDTH*2-1+0:0] tmp00_106_21;
	wire [WIDTH*2-1+0:0] tmp00_106_22;
	wire [WIDTH*2-1+0:0] tmp00_106_23;
	wire [WIDTH*2-1+0:0] tmp00_106_24;
	wire [WIDTH*2-1+0:0] tmp00_106_25;
	wire [WIDTH*2-1+0:0] tmp00_106_26;
	wire [WIDTH*2-1+0:0] tmp00_106_27;
	wire [WIDTH*2-1+0:0] tmp00_106_28;
	wire [WIDTH*2-1+0:0] tmp00_106_29;
	wire [WIDTH*2-1+0:0] tmp00_106_30;
	wire [WIDTH*2-1+0:0] tmp00_106_31;
	wire [WIDTH*2-1+0:0] tmp00_106_32;
	wire [WIDTH*2-1+0:0] tmp00_106_33;
	wire [WIDTH*2-1+0:0] tmp00_106_34;
	wire [WIDTH*2-1+0:0] tmp00_106_35;
	wire [WIDTH*2-1+0:0] tmp00_106_36;
	wire [WIDTH*2-1+0:0] tmp00_106_37;
	wire [WIDTH*2-1+0:0] tmp00_106_38;
	wire [WIDTH*2-1+0:0] tmp00_106_39;
	wire [WIDTH*2-1+0:0] tmp00_106_40;
	wire [WIDTH*2-1+0:0] tmp00_106_41;
	wire [WIDTH*2-1+0:0] tmp00_106_42;
	wire [WIDTH*2-1+0:0] tmp00_106_43;
	wire [WIDTH*2-1+0:0] tmp00_106_44;
	wire [WIDTH*2-1+0:0] tmp00_106_45;
	wire [WIDTH*2-1+0:0] tmp00_106_46;
	wire [WIDTH*2-1+0:0] tmp00_106_47;
	wire [WIDTH*2-1+0:0] tmp00_106_48;
	wire [WIDTH*2-1+0:0] tmp00_106_49;
	wire [WIDTH*2-1+0:0] tmp00_106_50;
	wire [WIDTH*2-1+0:0] tmp00_106_51;
	wire [WIDTH*2-1+0:0] tmp00_106_52;
	wire [WIDTH*2-1+0:0] tmp00_106_53;
	wire [WIDTH*2-1+0:0] tmp00_106_54;
	wire [WIDTH*2-1+0:0] tmp00_106_55;
	wire [WIDTH*2-1+0:0] tmp00_106_56;
	wire [WIDTH*2-1+0:0] tmp00_106_57;
	wire [WIDTH*2-1+0:0] tmp00_106_58;
	wire [WIDTH*2-1+0:0] tmp00_106_59;
	wire [WIDTH*2-1+0:0] tmp00_106_60;
	wire [WIDTH*2-1+0:0] tmp00_106_61;
	wire [WIDTH*2-1+0:0] tmp00_106_62;
	wire [WIDTH*2-1+0:0] tmp00_106_63;
	wire [WIDTH*2-1+0:0] tmp00_106_64;
	wire [WIDTH*2-1+0:0] tmp00_106_65;
	wire [WIDTH*2-1+0:0] tmp00_106_66;
	wire [WIDTH*2-1+0:0] tmp00_106_67;
	wire [WIDTH*2-1+0:0] tmp00_106_68;
	wire [WIDTH*2-1+0:0] tmp00_106_69;
	wire [WIDTH*2-1+0:0] tmp00_106_70;
	wire [WIDTH*2-1+0:0] tmp00_106_71;
	wire [WIDTH*2-1+0:0] tmp00_106_72;
	wire [WIDTH*2-1+0:0] tmp00_106_73;
	wire [WIDTH*2-1+0:0] tmp00_106_74;
	wire [WIDTH*2-1+0:0] tmp00_106_75;
	wire [WIDTH*2-1+0:0] tmp00_106_76;
	wire [WIDTH*2-1+0:0] tmp00_106_77;
	wire [WIDTH*2-1+0:0] tmp00_106_78;
	wire [WIDTH*2-1+0:0] tmp00_106_79;
	wire [WIDTH*2-1+0:0] tmp00_106_80;
	wire [WIDTH*2-1+0:0] tmp00_106_81;
	wire [WIDTH*2-1+0:0] tmp00_106_82;
	wire [WIDTH*2-1+0:0] tmp00_106_83;
	wire [WIDTH*2-1+0:0] tmp00_107_0;
	wire [WIDTH*2-1+0:0] tmp00_107_1;
	wire [WIDTH*2-1+0:0] tmp00_107_2;
	wire [WIDTH*2-1+0:0] tmp00_107_3;
	wire [WIDTH*2-1+0:0] tmp00_107_4;
	wire [WIDTH*2-1+0:0] tmp00_107_5;
	wire [WIDTH*2-1+0:0] tmp00_107_6;
	wire [WIDTH*2-1+0:0] tmp00_107_7;
	wire [WIDTH*2-1+0:0] tmp00_107_8;
	wire [WIDTH*2-1+0:0] tmp00_107_9;
	wire [WIDTH*2-1+0:0] tmp00_107_10;
	wire [WIDTH*2-1+0:0] tmp00_107_11;
	wire [WIDTH*2-1+0:0] tmp00_107_12;
	wire [WIDTH*2-1+0:0] tmp00_107_13;
	wire [WIDTH*2-1+0:0] tmp00_107_14;
	wire [WIDTH*2-1+0:0] tmp00_107_15;
	wire [WIDTH*2-1+0:0] tmp00_107_16;
	wire [WIDTH*2-1+0:0] tmp00_107_17;
	wire [WIDTH*2-1+0:0] tmp00_107_18;
	wire [WIDTH*2-1+0:0] tmp00_107_19;
	wire [WIDTH*2-1+0:0] tmp00_107_20;
	wire [WIDTH*2-1+0:0] tmp00_107_21;
	wire [WIDTH*2-1+0:0] tmp00_107_22;
	wire [WIDTH*2-1+0:0] tmp00_107_23;
	wire [WIDTH*2-1+0:0] tmp00_107_24;
	wire [WIDTH*2-1+0:0] tmp00_107_25;
	wire [WIDTH*2-1+0:0] tmp00_107_26;
	wire [WIDTH*2-1+0:0] tmp00_107_27;
	wire [WIDTH*2-1+0:0] tmp00_107_28;
	wire [WIDTH*2-1+0:0] tmp00_107_29;
	wire [WIDTH*2-1+0:0] tmp00_107_30;
	wire [WIDTH*2-1+0:0] tmp00_107_31;
	wire [WIDTH*2-1+0:0] tmp00_107_32;
	wire [WIDTH*2-1+0:0] tmp00_107_33;
	wire [WIDTH*2-1+0:0] tmp00_107_34;
	wire [WIDTH*2-1+0:0] tmp00_107_35;
	wire [WIDTH*2-1+0:0] tmp00_107_36;
	wire [WIDTH*2-1+0:0] tmp00_107_37;
	wire [WIDTH*2-1+0:0] tmp00_107_38;
	wire [WIDTH*2-1+0:0] tmp00_107_39;
	wire [WIDTH*2-1+0:0] tmp00_107_40;
	wire [WIDTH*2-1+0:0] tmp00_107_41;
	wire [WIDTH*2-1+0:0] tmp00_107_42;
	wire [WIDTH*2-1+0:0] tmp00_107_43;
	wire [WIDTH*2-1+0:0] tmp00_107_44;
	wire [WIDTH*2-1+0:0] tmp00_107_45;
	wire [WIDTH*2-1+0:0] tmp00_107_46;
	wire [WIDTH*2-1+0:0] tmp00_107_47;
	wire [WIDTH*2-1+0:0] tmp00_107_48;
	wire [WIDTH*2-1+0:0] tmp00_107_49;
	wire [WIDTH*2-1+0:0] tmp00_107_50;
	wire [WIDTH*2-1+0:0] tmp00_107_51;
	wire [WIDTH*2-1+0:0] tmp00_107_52;
	wire [WIDTH*2-1+0:0] tmp00_107_53;
	wire [WIDTH*2-1+0:0] tmp00_107_54;
	wire [WIDTH*2-1+0:0] tmp00_107_55;
	wire [WIDTH*2-1+0:0] tmp00_107_56;
	wire [WIDTH*2-1+0:0] tmp00_107_57;
	wire [WIDTH*2-1+0:0] tmp00_107_58;
	wire [WIDTH*2-1+0:0] tmp00_107_59;
	wire [WIDTH*2-1+0:0] tmp00_107_60;
	wire [WIDTH*2-1+0:0] tmp00_107_61;
	wire [WIDTH*2-1+0:0] tmp00_107_62;
	wire [WIDTH*2-1+0:0] tmp00_107_63;
	wire [WIDTH*2-1+0:0] tmp00_107_64;
	wire [WIDTH*2-1+0:0] tmp00_107_65;
	wire [WIDTH*2-1+0:0] tmp00_107_66;
	wire [WIDTH*2-1+0:0] tmp00_107_67;
	wire [WIDTH*2-1+0:0] tmp00_107_68;
	wire [WIDTH*2-1+0:0] tmp00_107_69;
	wire [WIDTH*2-1+0:0] tmp00_107_70;
	wire [WIDTH*2-1+0:0] tmp00_107_71;
	wire [WIDTH*2-1+0:0] tmp00_107_72;
	wire [WIDTH*2-1+0:0] tmp00_107_73;
	wire [WIDTH*2-1+0:0] tmp00_107_74;
	wire [WIDTH*2-1+0:0] tmp00_107_75;
	wire [WIDTH*2-1+0:0] tmp00_107_76;
	wire [WIDTH*2-1+0:0] tmp00_107_77;
	wire [WIDTH*2-1+0:0] tmp00_107_78;
	wire [WIDTH*2-1+0:0] tmp00_107_79;
	wire [WIDTH*2-1+0:0] tmp00_107_80;
	wire [WIDTH*2-1+0:0] tmp00_107_81;
	wire [WIDTH*2-1+0:0] tmp00_107_82;
	wire [WIDTH*2-1+0:0] tmp00_107_83;
	wire [WIDTH*2-1+0:0] tmp00_108_0;
	wire [WIDTH*2-1+0:0] tmp00_108_1;
	wire [WIDTH*2-1+0:0] tmp00_108_2;
	wire [WIDTH*2-1+0:0] tmp00_108_3;
	wire [WIDTH*2-1+0:0] tmp00_108_4;
	wire [WIDTH*2-1+0:0] tmp00_108_5;
	wire [WIDTH*2-1+0:0] tmp00_108_6;
	wire [WIDTH*2-1+0:0] tmp00_108_7;
	wire [WIDTH*2-1+0:0] tmp00_108_8;
	wire [WIDTH*2-1+0:0] tmp00_108_9;
	wire [WIDTH*2-1+0:0] tmp00_108_10;
	wire [WIDTH*2-1+0:0] tmp00_108_11;
	wire [WIDTH*2-1+0:0] tmp00_108_12;
	wire [WIDTH*2-1+0:0] tmp00_108_13;
	wire [WIDTH*2-1+0:0] tmp00_108_14;
	wire [WIDTH*2-1+0:0] tmp00_108_15;
	wire [WIDTH*2-1+0:0] tmp00_108_16;
	wire [WIDTH*2-1+0:0] tmp00_108_17;
	wire [WIDTH*2-1+0:0] tmp00_108_18;
	wire [WIDTH*2-1+0:0] tmp00_108_19;
	wire [WIDTH*2-1+0:0] tmp00_108_20;
	wire [WIDTH*2-1+0:0] tmp00_108_21;
	wire [WIDTH*2-1+0:0] tmp00_108_22;
	wire [WIDTH*2-1+0:0] tmp00_108_23;
	wire [WIDTH*2-1+0:0] tmp00_108_24;
	wire [WIDTH*2-1+0:0] tmp00_108_25;
	wire [WIDTH*2-1+0:0] tmp00_108_26;
	wire [WIDTH*2-1+0:0] tmp00_108_27;
	wire [WIDTH*2-1+0:0] tmp00_108_28;
	wire [WIDTH*2-1+0:0] tmp00_108_29;
	wire [WIDTH*2-1+0:0] tmp00_108_30;
	wire [WIDTH*2-1+0:0] tmp00_108_31;
	wire [WIDTH*2-1+0:0] tmp00_108_32;
	wire [WIDTH*2-1+0:0] tmp00_108_33;
	wire [WIDTH*2-1+0:0] tmp00_108_34;
	wire [WIDTH*2-1+0:0] tmp00_108_35;
	wire [WIDTH*2-1+0:0] tmp00_108_36;
	wire [WIDTH*2-1+0:0] tmp00_108_37;
	wire [WIDTH*2-1+0:0] tmp00_108_38;
	wire [WIDTH*2-1+0:0] tmp00_108_39;
	wire [WIDTH*2-1+0:0] tmp00_108_40;
	wire [WIDTH*2-1+0:0] tmp00_108_41;
	wire [WIDTH*2-1+0:0] tmp00_108_42;
	wire [WIDTH*2-1+0:0] tmp00_108_43;
	wire [WIDTH*2-1+0:0] tmp00_108_44;
	wire [WIDTH*2-1+0:0] tmp00_108_45;
	wire [WIDTH*2-1+0:0] tmp00_108_46;
	wire [WIDTH*2-1+0:0] tmp00_108_47;
	wire [WIDTH*2-1+0:0] tmp00_108_48;
	wire [WIDTH*2-1+0:0] tmp00_108_49;
	wire [WIDTH*2-1+0:0] tmp00_108_50;
	wire [WIDTH*2-1+0:0] tmp00_108_51;
	wire [WIDTH*2-1+0:0] tmp00_108_52;
	wire [WIDTH*2-1+0:0] tmp00_108_53;
	wire [WIDTH*2-1+0:0] tmp00_108_54;
	wire [WIDTH*2-1+0:0] tmp00_108_55;
	wire [WIDTH*2-1+0:0] tmp00_108_56;
	wire [WIDTH*2-1+0:0] tmp00_108_57;
	wire [WIDTH*2-1+0:0] tmp00_108_58;
	wire [WIDTH*2-1+0:0] tmp00_108_59;
	wire [WIDTH*2-1+0:0] tmp00_108_60;
	wire [WIDTH*2-1+0:0] tmp00_108_61;
	wire [WIDTH*2-1+0:0] tmp00_108_62;
	wire [WIDTH*2-1+0:0] tmp00_108_63;
	wire [WIDTH*2-1+0:0] tmp00_108_64;
	wire [WIDTH*2-1+0:0] tmp00_108_65;
	wire [WIDTH*2-1+0:0] tmp00_108_66;
	wire [WIDTH*2-1+0:0] tmp00_108_67;
	wire [WIDTH*2-1+0:0] tmp00_108_68;
	wire [WIDTH*2-1+0:0] tmp00_108_69;
	wire [WIDTH*2-1+0:0] tmp00_108_70;
	wire [WIDTH*2-1+0:0] tmp00_108_71;
	wire [WIDTH*2-1+0:0] tmp00_108_72;
	wire [WIDTH*2-1+0:0] tmp00_108_73;
	wire [WIDTH*2-1+0:0] tmp00_108_74;
	wire [WIDTH*2-1+0:0] tmp00_108_75;
	wire [WIDTH*2-1+0:0] tmp00_108_76;
	wire [WIDTH*2-1+0:0] tmp00_108_77;
	wire [WIDTH*2-1+0:0] tmp00_108_78;
	wire [WIDTH*2-1+0:0] tmp00_108_79;
	wire [WIDTH*2-1+0:0] tmp00_108_80;
	wire [WIDTH*2-1+0:0] tmp00_108_81;
	wire [WIDTH*2-1+0:0] tmp00_108_82;
	wire [WIDTH*2-1+0:0] tmp00_108_83;
	wire [WIDTH*2-1+0:0] tmp00_109_0;
	wire [WIDTH*2-1+0:0] tmp00_109_1;
	wire [WIDTH*2-1+0:0] tmp00_109_2;
	wire [WIDTH*2-1+0:0] tmp00_109_3;
	wire [WIDTH*2-1+0:0] tmp00_109_4;
	wire [WIDTH*2-1+0:0] tmp00_109_5;
	wire [WIDTH*2-1+0:0] tmp00_109_6;
	wire [WIDTH*2-1+0:0] tmp00_109_7;
	wire [WIDTH*2-1+0:0] tmp00_109_8;
	wire [WIDTH*2-1+0:0] tmp00_109_9;
	wire [WIDTH*2-1+0:0] tmp00_109_10;
	wire [WIDTH*2-1+0:0] tmp00_109_11;
	wire [WIDTH*2-1+0:0] tmp00_109_12;
	wire [WIDTH*2-1+0:0] tmp00_109_13;
	wire [WIDTH*2-1+0:0] tmp00_109_14;
	wire [WIDTH*2-1+0:0] tmp00_109_15;
	wire [WIDTH*2-1+0:0] tmp00_109_16;
	wire [WIDTH*2-1+0:0] tmp00_109_17;
	wire [WIDTH*2-1+0:0] tmp00_109_18;
	wire [WIDTH*2-1+0:0] tmp00_109_19;
	wire [WIDTH*2-1+0:0] tmp00_109_20;
	wire [WIDTH*2-1+0:0] tmp00_109_21;
	wire [WIDTH*2-1+0:0] tmp00_109_22;
	wire [WIDTH*2-1+0:0] tmp00_109_23;
	wire [WIDTH*2-1+0:0] tmp00_109_24;
	wire [WIDTH*2-1+0:0] tmp00_109_25;
	wire [WIDTH*2-1+0:0] tmp00_109_26;
	wire [WIDTH*2-1+0:0] tmp00_109_27;
	wire [WIDTH*2-1+0:0] tmp00_109_28;
	wire [WIDTH*2-1+0:0] tmp00_109_29;
	wire [WIDTH*2-1+0:0] tmp00_109_30;
	wire [WIDTH*2-1+0:0] tmp00_109_31;
	wire [WIDTH*2-1+0:0] tmp00_109_32;
	wire [WIDTH*2-1+0:0] tmp00_109_33;
	wire [WIDTH*2-1+0:0] tmp00_109_34;
	wire [WIDTH*2-1+0:0] tmp00_109_35;
	wire [WIDTH*2-1+0:0] tmp00_109_36;
	wire [WIDTH*2-1+0:0] tmp00_109_37;
	wire [WIDTH*2-1+0:0] tmp00_109_38;
	wire [WIDTH*2-1+0:0] tmp00_109_39;
	wire [WIDTH*2-1+0:0] tmp00_109_40;
	wire [WIDTH*2-1+0:0] tmp00_109_41;
	wire [WIDTH*2-1+0:0] tmp00_109_42;
	wire [WIDTH*2-1+0:0] tmp00_109_43;
	wire [WIDTH*2-1+0:0] tmp00_109_44;
	wire [WIDTH*2-1+0:0] tmp00_109_45;
	wire [WIDTH*2-1+0:0] tmp00_109_46;
	wire [WIDTH*2-1+0:0] tmp00_109_47;
	wire [WIDTH*2-1+0:0] tmp00_109_48;
	wire [WIDTH*2-1+0:0] tmp00_109_49;
	wire [WIDTH*2-1+0:0] tmp00_109_50;
	wire [WIDTH*2-1+0:0] tmp00_109_51;
	wire [WIDTH*2-1+0:0] tmp00_109_52;
	wire [WIDTH*2-1+0:0] tmp00_109_53;
	wire [WIDTH*2-1+0:0] tmp00_109_54;
	wire [WIDTH*2-1+0:0] tmp00_109_55;
	wire [WIDTH*2-1+0:0] tmp00_109_56;
	wire [WIDTH*2-1+0:0] tmp00_109_57;
	wire [WIDTH*2-1+0:0] tmp00_109_58;
	wire [WIDTH*2-1+0:0] tmp00_109_59;
	wire [WIDTH*2-1+0:0] tmp00_109_60;
	wire [WIDTH*2-1+0:0] tmp00_109_61;
	wire [WIDTH*2-1+0:0] tmp00_109_62;
	wire [WIDTH*2-1+0:0] tmp00_109_63;
	wire [WIDTH*2-1+0:0] tmp00_109_64;
	wire [WIDTH*2-1+0:0] tmp00_109_65;
	wire [WIDTH*2-1+0:0] tmp00_109_66;
	wire [WIDTH*2-1+0:0] tmp00_109_67;
	wire [WIDTH*2-1+0:0] tmp00_109_68;
	wire [WIDTH*2-1+0:0] tmp00_109_69;
	wire [WIDTH*2-1+0:0] tmp00_109_70;
	wire [WIDTH*2-1+0:0] tmp00_109_71;
	wire [WIDTH*2-1+0:0] tmp00_109_72;
	wire [WIDTH*2-1+0:0] tmp00_109_73;
	wire [WIDTH*2-1+0:0] tmp00_109_74;
	wire [WIDTH*2-1+0:0] tmp00_109_75;
	wire [WIDTH*2-1+0:0] tmp00_109_76;
	wire [WIDTH*2-1+0:0] tmp00_109_77;
	wire [WIDTH*2-1+0:0] tmp00_109_78;
	wire [WIDTH*2-1+0:0] tmp00_109_79;
	wire [WIDTH*2-1+0:0] tmp00_109_80;
	wire [WIDTH*2-1+0:0] tmp00_109_81;
	wire [WIDTH*2-1+0:0] tmp00_109_82;
	wire [WIDTH*2-1+0:0] tmp00_109_83;
	wire [WIDTH*2-1+0:0] tmp00_110_0;
	wire [WIDTH*2-1+0:0] tmp00_110_1;
	wire [WIDTH*2-1+0:0] tmp00_110_2;
	wire [WIDTH*2-1+0:0] tmp00_110_3;
	wire [WIDTH*2-1+0:0] tmp00_110_4;
	wire [WIDTH*2-1+0:0] tmp00_110_5;
	wire [WIDTH*2-1+0:0] tmp00_110_6;
	wire [WIDTH*2-1+0:0] tmp00_110_7;
	wire [WIDTH*2-1+0:0] tmp00_110_8;
	wire [WIDTH*2-1+0:0] tmp00_110_9;
	wire [WIDTH*2-1+0:0] tmp00_110_10;
	wire [WIDTH*2-1+0:0] tmp00_110_11;
	wire [WIDTH*2-1+0:0] tmp00_110_12;
	wire [WIDTH*2-1+0:0] tmp00_110_13;
	wire [WIDTH*2-1+0:0] tmp00_110_14;
	wire [WIDTH*2-1+0:0] tmp00_110_15;
	wire [WIDTH*2-1+0:0] tmp00_110_16;
	wire [WIDTH*2-1+0:0] tmp00_110_17;
	wire [WIDTH*2-1+0:0] tmp00_110_18;
	wire [WIDTH*2-1+0:0] tmp00_110_19;
	wire [WIDTH*2-1+0:0] tmp00_110_20;
	wire [WIDTH*2-1+0:0] tmp00_110_21;
	wire [WIDTH*2-1+0:0] tmp00_110_22;
	wire [WIDTH*2-1+0:0] tmp00_110_23;
	wire [WIDTH*2-1+0:0] tmp00_110_24;
	wire [WIDTH*2-1+0:0] tmp00_110_25;
	wire [WIDTH*2-1+0:0] tmp00_110_26;
	wire [WIDTH*2-1+0:0] tmp00_110_27;
	wire [WIDTH*2-1+0:0] tmp00_110_28;
	wire [WIDTH*2-1+0:0] tmp00_110_29;
	wire [WIDTH*2-1+0:0] tmp00_110_30;
	wire [WIDTH*2-1+0:0] tmp00_110_31;
	wire [WIDTH*2-1+0:0] tmp00_110_32;
	wire [WIDTH*2-1+0:0] tmp00_110_33;
	wire [WIDTH*2-1+0:0] tmp00_110_34;
	wire [WIDTH*2-1+0:0] tmp00_110_35;
	wire [WIDTH*2-1+0:0] tmp00_110_36;
	wire [WIDTH*2-1+0:0] tmp00_110_37;
	wire [WIDTH*2-1+0:0] tmp00_110_38;
	wire [WIDTH*2-1+0:0] tmp00_110_39;
	wire [WIDTH*2-1+0:0] tmp00_110_40;
	wire [WIDTH*2-1+0:0] tmp00_110_41;
	wire [WIDTH*2-1+0:0] tmp00_110_42;
	wire [WIDTH*2-1+0:0] tmp00_110_43;
	wire [WIDTH*2-1+0:0] tmp00_110_44;
	wire [WIDTH*2-1+0:0] tmp00_110_45;
	wire [WIDTH*2-1+0:0] tmp00_110_46;
	wire [WIDTH*2-1+0:0] tmp00_110_47;
	wire [WIDTH*2-1+0:0] tmp00_110_48;
	wire [WIDTH*2-1+0:0] tmp00_110_49;
	wire [WIDTH*2-1+0:0] tmp00_110_50;
	wire [WIDTH*2-1+0:0] tmp00_110_51;
	wire [WIDTH*2-1+0:0] tmp00_110_52;
	wire [WIDTH*2-1+0:0] tmp00_110_53;
	wire [WIDTH*2-1+0:0] tmp00_110_54;
	wire [WIDTH*2-1+0:0] tmp00_110_55;
	wire [WIDTH*2-1+0:0] tmp00_110_56;
	wire [WIDTH*2-1+0:0] tmp00_110_57;
	wire [WIDTH*2-1+0:0] tmp00_110_58;
	wire [WIDTH*2-1+0:0] tmp00_110_59;
	wire [WIDTH*2-1+0:0] tmp00_110_60;
	wire [WIDTH*2-1+0:0] tmp00_110_61;
	wire [WIDTH*2-1+0:0] tmp00_110_62;
	wire [WIDTH*2-1+0:0] tmp00_110_63;
	wire [WIDTH*2-1+0:0] tmp00_110_64;
	wire [WIDTH*2-1+0:0] tmp00_110_65;
	wire [WIDTH*2-1+0:0] tmp00_110_66;
	wire [WIDTH*2-1+0:0] tmp00_110_67;
	wire [WIDTH*2-1+0:0] tmp00_110_68;
	wire [WIDTH*2-1+0:0] tmp00_110_69;
	wire [WIDTH*2-1+0:0] tmp00_110_70;
	wire [WIDTH*2-1+0:0] tmp00_110_71;
	wire [WIDTH*2-1+0:0] tmp00_110_72;
	wire [WIDTH*2-1+0:0] tmp00_110_73;
	wire [WIDTH*2-1+0:0] tmp00_110_74;
	wire [WIDTH*2-1+0:0] tmp00_110_75;
	wire [WIDTH*2-1+0:0] tmp00_110_76;
	wire [WIDTH*2-1+0:0] tmp00_110_77;
	wire [WIDTH*2-1+0:0] tmp00_110_78;
	wire [WIDTH*2-1+0:0] tmp00_110_79;
	wire [WIDTH*2-1+0:0] tmp00_110_80;
	wire [WIDTH*2-1+0:0] tmp00_110_81;
	wire [WIDTH*2-1+0:0] tmp00_110_82;
	wire [WIDTH*2-1+0:0] tmp00_110_83;
	wire [WIDTH*2-1+0:0] tmp00_111_0;
	wire [WIDTH*2-1+0:0] tmp00_111_1;
	wire [WIDTH*2-1+0:0] tmp00_111_2;
	wire [WIDTH*2-1+0:0] tmp00_111_3;
	wire [WIDTH*2-1+0:0] tmp00_111_4;
	wire [WIDTH*2-1+0:0] tmp00_111_5;
	wire [WIDTH*2-1+0:0] tmp00_111_6;
	wire [WIDTH*2-1+0:0] tmp00_111_7;
	wire [WIDTH*2-1+0:0] tmp00_111_8;
	wire [WIDTH*2-1+0:0] tmp00_111_9;
	wire [WIDTH*2-1+0:0] tmp00_111_10;
	wire [WIDTH*2-1+0:0] tmp00_111_11;
	wire [WIDTH*2-1+0:0] tmp00_111_12;
	wire [WIDTH*2-1+0:0] tmp00_111_13;
	wire [WIDTH*2-1+0:0] tmp00_111_14;
	wire [WIDTH*2-1+0:0] tmp00_111_15;
	wire [WIDTH*2-1+0:0] tmp00_111_16;
	wire [WIDTH*2-1+0:0] tmp00_111_17;
	wire [WIDTH*2-1+0:0] tmp00_111_18;
	wire [WIDTH*2-1+0:0] tmp00_111_19;
	wire [WIDTH*2-1+0:0] tmp00_111_20;
	wire [WIDTH*2-1+0:0] tmp00_111_21;
	wire [WIDTH*2-1+0:0] tmp00_111_22;
	wire [WIDTH*2-1+0:0] tmp00_111_23;
	wire [WIDTH*2-1+0:0] tmp00_111_24;
	wire [WIDTH*2-1+0:0] tmp00_111_25;
	wire [WIDTH*2-1+0:0] tmp00_111_26;
	wire [WIDTH*2-1+0:0] tmp00_111_27;
	wire [WIDTH*2-1+0:0] tmp00_111_28;
	wire [WIDTH*2-1+0:0] tmp00_111_29;
	wire [WIDTH*2-1+0:0] tmp00_111_30;
	wire [WIDTH*2-1+0:0] tmp00_111_31;
	wire [WIDTH*2-1+0:0] tmp00_111_32;
	wire [WIDTH*2-1+0:0] tmp00_111_33;
	wire [WIDTH*2-1+0:0] tmp00_111_34;
	wire [WIDTH*2-1+0:0] tmp00_111_35;
	wire [WIDTH*2-1+0:0] tmp00_111_36;
	wire [WIDTH*2-1+0:0] tmp00_111_37;
	wire [WIDTH*2-1+0:0] tmp00_111_38;
	wire [WIDTH*2-1+0:0] tmp00_111_39;
	wire [WIDTH*2-1+0:0] tmp00_111_40;
	wire [WIDTH*2-1+0:0] tmp00_111_41;
	wire [WIDTH*2-1+0:0] tmp00_111_42;
	wire [WIDTH*2-1+0:0] tmp00_111_43;
	wire [WIDTH*2-1+0:0] tmp00_111_44;
	wire [WIDTH*2-1+0:0] tmp00_111_45;
	wire [WIDTH*2-1+0:0] tmp00_111_46;
	wire [WIDTH*2-1+0:0] tmp00_111_47;
	wire [WIDTH*2-1+0:0] tmp00_111_48;
	wire [WIDTH*2-1+0:0] tmp00_111_49;
	wire [WIDTH*2-1+0:0] tmp00_111_50;
	wire [WIDTH*2-1+0:0] tmp00_111_51;
	wire [WIDTH*2-1+0:0] tmp00_111_52;
	wire [WIDTH*2-1+0:0] tmp00_111_53;
	wire [WIDTH*2-1+0:0] tmp00_111_54;
	wire [WIDTH*2-1+0:0] tmp00_111_55;
	wire [WIDTH*2-1+0:0] tmp00_111_56;
	wire [WIDTH*2-1+0:0] tmp00_111_57;
	wire [WIDTH*2-1+0:0] tmp00_111_58;
	wire [WIDTH*2-1+0:0] tmp00_111_59;
	wire [WIDTH*2-1+0:0] tmp00_111_60;
	wire [WIDTH*2-1+0:0] tmp00_111_61;
	wire [WIDTH*2-1+0:0] tmp00_111_62;
	wire [WIDTH*2-1+0:0] tmp00_111_63;
	wire [WIDTH*2-1+0:0] tmp00_111_64;
	wire [WIDTH*2-1+0:0] tmp00_111_65;
	wire [WIDTH*2-1+0:0] tmp00_111_66;
	wire [WIDTH*2-1+0:0] tmp00_111_67;
	wire [WIDTH*2-1+0:0] tmp00_111_68;
	wire [WIDTH*2-1+0:0] tmp00_111_69;
	wire [WIDTH*2-1+0:0] tmp00_111_70;
	wire [WIDTH*2-1+0:0] tmp00_111_71;
	wire [WIDTH*2-1+0:0] tmp00_111_72;
	wire [WIDTH*2-1+0:0] tmp00_111_73;
	wire [WIDTH*2-1+0:0] tmp00_111_74;
	wire [WIDTH*2-1+0:0] tmp00_111_75;
	wire [WIDTH*2-1+0:0] tmp00_111_76;
	wire [WIDTH*2-1+0:0] tmp00_111_77;
	wire [WIDTH*2-1+0:0] tmp00_111_78;
	wire [WIDTH*2-1+0:0] tmp00_111_79;
	wire [WIDTH*2-1+0:0] tmp00_111_80;
	wire [WIDTH*2-1+0:0] tmp00_111_81;
	wire [WIDTH*2-1+0:0] tmp00_111_82;
	wire [WIDTH*2-1+0:0] tmp00_111_83;
	wire [WIDTH*2-1+0:0] tmp00_112_0;
	wire [WIDTH*2-1+0:0] tmp00_112_1;
	wire [WIDTH*2-1+0:0] tmp00_112_2;
	wire [WIDTH*2-1+0:0] tmp00_112_3;
	wire [WIDTH*2-1+0:0] tmp00_112_4;
	wire [WIDTH*2-1+0:0] tmp00_112_5;
	wire [WIDTH*2-1+0:0] tmp00_112_6;
	wire [WIDTH*2-1+0:0] tmp00_112_7;
	wire [WIDTH*2-1+0:0] tmp00_112_8;
	wire [WIDTH*2-1+0:0] tmp00_112_9;
	wire [WIDTH*2-1+0:0] tmp00_112_10;
	wire [WIDTH*2-1+0:0] tmp00_112_11;
	wire [WIDTH*2-1+0:0] tmp00_112_12;
	wire [WIDTH*2-1+0:0] tmp00_112_13;
	wire [WIDTH*2-1+0:0] tmp00_112_14;
	wire [WIDTH*2-1+0:0] tmp00_112_15;
	wire [WIDTH*2-1+0:0] tmp00_112_16;
	wire [WIDTH*2-1+0:0] tmp00_112_17;
	wire [WIDTH*2-1+0:0] tmp00_112_18;
	wire [WIDTH*2-1+0:0] tmp00_112_19;
	wire [WIDTH*2-1+0:0] tmp00_112_20;
	wire [WIDTH*2-1+0:0] tmp00_112_21;
	wire [WIDTH*2-1+0:0] tmp00_112_22;
	wire [WIDTH*2-1+0:0] tmp00_112_23;
	wire [WIDTH*2-1+0:0] tmp00_112_24;
	wire [WIDTH*2-1+0:0] tmp00_112_25;
	wire [WIDTH*2-1+0:0] tmp00_112_26;
	wire [WIDTH*2-1+0:0] tmp00_112_27;
	wire [WIDTH*2-1+0:0] tmp00_112_28;
	wire [WIDTH*2-1+0:0] tmp00_112_29;
	wire [WIDTH*2-1+0:0] tmp00_112_30;
	wire [WIDTH*2-1+0:0] tmp00_112_31;
	wire [WIDTH*2-1+0:0] tmp00_112_32;
	wire [WIDTH*2-1+0:0] tmp00_112_33;
	wire [WIDTH*2-1+0:0] tmp00_112_34;
	wire [WIDTH*2-1+0:0] tmp00_112_35;
	wire [WIDTH*2-1+0:0] tmp00_112_36;
	wire [WIDTH*2-1+0:0] tmp00_112_37;
	wire [WIDTH*2-1+0:0] tmp00_112_38;
	wire [WIDTH*2-1+0:0] tmp00_112_39;
	wire [WIDTH*2-1+0:0] tmp00_112_40;
	wire [WIDTH*2-1+0:0] tmp00_112_41;
	wire [WIDTH*2-1+0:0] tmp00_112_42;
	wire [WIDTH*2-1+0:0] tmp00_112_43;
	wire [WIDTH*2-1+0:0] tmp00_112_44;
	wire [WIDTH*2-1+0:0] tmp00_112_45;
	wire [WIDTH*2-1+0:0] tmp00_112_46;
	wire [WIDTH*2-1+0:0] tmp00_112_47;
	wire [WIDTH*2-1+0:0] tmp00_112_48;
	wire [WIDTH*2-1+0:0] tmp00_112_49;
	wire [WIDTH*2-1+0:0] tmp00_112_50;
	wire [WIDTH*2-1+0:0] tmp00_112_51;
	wire [WIDTH*2-1+0:0] tmp00_112_52;
	wire [WIDTH*2-1+0:0] tmp00_112_53;
	wire [WIDTH*2-1+0:0] tmp00_112_54;
	wire [WIDTH*2-1+0:0] tmp00_112_55;
	wire [WIDTH*2-1+0:0] tmp00_112_56;
	wire [WIDTH*2-1+0:0] tmp00_112_57;
	wire [WIDTH*2-1+0:0] tmp00_112_58;
	wire [WIDTH*2-1+0:0] tmp00_112_59;
	wire [WIDTH*2-1+0:0] tmp00_112_60;
	wire [WIDTH*2-1+0:0] tmp00_112_61;
	wire [WIDTH*2-1+0:0] tmp00_112_62;
	wire [WIDTH*2-1+0:0] tmp00_112_63;
	wire [WIDTH*2-1+0:0] tmp00_112_64;
	wire [WIDTH*2-1+0:0] tmp00_112_65;
	wire [WIDTH*2-1+0:0] tmp00_112_66;
	wire [WIDTH*2-1+0:0] tmp00_112_67;
	wire [WIDTH*2-1+0:0] tmp00_112_68;
	wire [WIDTH*2-1+0:0] tmp00_112_69;
	wire [WIDTH*2-1+0:0] tmp00_112_70;
	wire [WIDTH*2-1+0:0] tmp00_112_71;
	wire [WIDTH*2-1+0:0] tmp00_112_72;
	wire [WIDTH*2-1+0:0] tmp00_112_73;
	wire [WIDTH*2-1+0:0] tmp00_112_74;
	wire [WIDTH*2-1+0:0] tmp00_112_75;
	wire [WIDTH*2-1+0:0] tmp00_112_76;
	wire [WIDTH*2-1+0:0] tmp00_112_77;
	wire [WIDTH*2-1+0:0] tmp00_112_78;
	wire [WIDTH*2-1+0:0] tmp00_112_79;
	wire [WIDTH*2-1+0:0] tmp00_112_80;
	wire [WIDTH*2-1+0:0] tmp00_112_81;
	wire [WIDTH*2-1+0:0] tmp00_112_82;
	wire [WIDTH*2-1+0:0] tmp00_112_83;
	wire [WIDTH*2-1+0:0] tmp00_113_0;
	wire [WIDTH*2-1+0:0] tmp00_113_1;
	wire [WIDTH*2-1+0:0] tmp00_113_2;
	wire [WIDTH*2-1+0:0] tmp00_113_3;
	wire [WIDTH*2-1+0:0] tmp00_113_4;
	wire [WIDTH*2-1+0:0] tmp00_113_5;
	wire [WIDTH*2-1+0:0] tmp00_113_6;
	wire [WIDTH*2-1+0:0] tmp00_113_7;
	wire [WIDTH*2-1+0:0] tmp00_113_8;
	wire [WIDTH*2-1+0:0] tmp00_113_9;
	wire [WIDTH*2-1+0:0] tmp00_113_10;
	wire [WIDTH*2-1+0:0] tmp00_113_11;
	wire [WIDTH*2-1+0:0] tmp00_113_12;
	wire [WIDTH*2-1+0:0] tmp00_113_13;
	wire [WIDTH*2-1+0:0] tmp00_113_14;
	wire [WIDTH*2-1+0:0] tmp00_113_15;
	wire [WIDTH*2-1+0:0] tmp00_113_16;
	wire [WIDTH*2-1+0:0] tmp00_113_17;
	wire [WIDTH*2-1+0:0] tmp00_113_18;
	wire [WIDTH*2-1+0:0] tmp00_113_19;
	wire [WIDTH*2-1+0:0] tmp00_113_20;
	wire [WIDTH*2-1+0:0] tmp00_113_21;
	wire [WIDTH*2-1+0:0] tmp00_113_22;
	wire [WIDTH*2-1+0:0] tmp00_113_23;
	wire [WIDTH*2-1+0:0] tmp00_113_24;
	wire [WIDTH*2-1+0:0] tmp00_113_25;
	wire [WIDTH*2-1+0:0] tmp00_113_26;
	wire [WIDTH*2-1+0:0] tmp00_113_27;
	wire [WIDTH*2-1+0:0] tmp00_113_28;
	wire [WIDTH*2-1+0:0] tmp00_113_29;
	wire [WIDTH*2-1+0:0] tmp00_113_30;
	wire [WIDTH*2-1+0:0] tmp00_113_31;
	wire [WIDTH*2-1+0:0] tmp00_113_32;
	wire [WIDTH*2-1+0:0] tmp00_113_33;
	wire [WIDTH*2-1+0:0] tmp00_113_34;
	wire [WIDTH*2-1+0:0] tmp00_113_35;
	wire [WIDTH*2-1+0:0] tmp00_113_36;
	wire [WIDTH*2-1+0:0] tmp00_113_37;
	wire [WIDTH*2-1+0:0] tmp00_113_38;
	wire [WIDTH*2-1+0:0] tmp00_113_39;
	wire [WIDTH*2-1+0:0] tmp00_113_40;
	wire [WIDTH*2-1+0:0] tmp00_113_41;
	wire [WIDTH*2-1+0:0] tmp00_113_42;
	wire [WIDTH*2-1+0:0] tmp00_113_43;
	wire [WIDTH*2-1+0:0] tmp00_113_44;
	wire [WIDTH*2-1+0:0] tmp00_113_45;
	wire [WIDTH*2-1+0:0] tmp00_113_46;
	wire [WIDTH*2-1+0:0] tmp00_113_47;
	wire [WIDTH*2-1+0:0] tmp00_113_48;
	wire [WIDTH*2-1+0:0] tmp00_113_49;
	wire [WIDTH*2-1+0:0] tmp00_113_50;
	wire [WIDTH*2-1+0:0] tmp00_113_51;
	wire [WIDTH*2-1+0:0] tmp00_113_52;
	wire [WIDTH*2-1+0:0] tmp00_113_53;
	wire [WIDTH*2-1+0:0] tmp00_113_54;
	wire [WIDTH*2-1+0:0] tmp00_113_55;
	wire [WIDTH*2-1+0:0] tmp00_113_56;
	wire [WIDTH*2-1+0:0] tmp00_113_57;
	wire [WIDTH*2-1+0:0] tmp00_113_58;
	wire [WIDTH*2-1+0:0] tmp00_113_59;
	wire [WIDTH*2-1+0:0] tmp00_113_60;
	wire [WIDTH*2-1+0:0] tmp00_113_61;
	wire [WIDTH*2-1+0:0] tmp00_113_62;
	wire [WIDTH*2-1+0:0] tmp00_113_63;
	wire [WIDTH*2-1+0:0] tmp00_113_64;
	wire [WIDTH*2-1+0:0] tmp00_113_65;
	wire [WIDTH*2-1+0:0] tmp00_113_66;
	wire [WIDTH*2-1+0:0] tmp00_113_67;
	wire [WIDTH*2-1+0:0] tmp00_113_68;
	wire [WIDTH*2-1+0:0] tmp00_113_69;
	wire [WIDTH*2-1+0:0] tmp00_113_70;
	wire [WIDTH*2-1+0:0] tmp00_113_71;
	wire [WIDTH*2-1+0:0] tmp00_113_72;
	wire [WIDTH*2-1+0:0] tmp00_113_73;
	wire [WIDTH*2-1+0:0] tmp00_113_74;
	wire [WIDTH*2-1+0:0] tmp00_113_75;
	wire [WIDTH*2-1+0:0] tmp00_113_76;
	wire [WIDTH*2-1+0:0] tmp00_113_77;
	wire [WIDTH*2-1+0:0] tmp00_113_78;
	wire [WIDTH*2-1+0:0] tmp00_113_79;
	wire [WIDTH*2-1+0:0] tmp00_113_80;
	wire [WIDTH*2-1+0:0] tmp00_113_81;
	wire [WIDTH*2-1+0:0] tmp00_113_82;
	wire [WIDTH*2-1+0:0] tmp00_113_83;
	wire [WIDTH*2-1+0:0] tmp00_114_0;
	wire [WIDTH*2-1+0:0] tmp00_114_1;
	wire [WIDTH*2-1+0:0] tmp00_114_2;
	wire [WIDTH*2-1+0:0] tmp00_114_3;
	wire [WIDTH*2-1+0:0] tmp00_114_4;
	wire [WIDTH*2-1+0:0] tmp00_114_5;
	wire [WIDTH*2-1+0:0] tmp00_114_6;
	wire [WIDTH*2-1+0:0] tmp00_114_7;
	wire [WIDTH*2-1+0:0] tmp00_114_8;
	wire [WIDTH*2-1+0:0] tmp00_114_9;
	wire [WIDTH*2-1+0:0] tmp00_114_10;
	wire [WIDTH*2-1+0:0] tmp00_114_11;
	wire [WIDTH*2-1+0:0] tmp00_114_12;
	wire [WIDTH*2-1+0:0] tmp00_114_13;
	wire [WIDTH*2-1+0:0] tmp00_114_14;
	wire [WIDTH*2-1+0:0] tmp00_114_15;
	wire [WIDTH*2-1+0:0] tmp00_114_16;
	wire [WIDTH*2-1+0:0] tmp00_114_17;
	wire [WIDTH*2-1+0:0] tmp00_114_18;
	wire [WIDTH*2-1+0:0] tmp00_114_19;
	wire [WIDTH*2-1+0:0] tmp00_114_20;
	wire [WIDTH*2-1+0:0] tmp00_114_21;
	wire [WIDTH*2-1+0:0] tmp00_114_22;
	wire [WIDTH*2-1+0:0] tmp00_114_23;
	wire [WIDTH*2-1+0:0] tmp00_114_24;
	wire [WIDTH*2-1+0:0] tmp00_114_25;
	wire [WIDTH*2-1+0:0] tmp00_114_26;
	wire [WIDTH*2-1+0:0] tmp00_114_27;
	wire [WIDTH*2-1+0:0] tmp00_114_28;
	wire [WIDTH*2-1+0:0] tmp00_114_29;
	wire [WIDTH*2-1+0:0] tmp00_114_30;
	wire [WIDTH*2-1+0:0] tmp00_114_31;
	wire [WIDTH*2-1+0:0] tmp00_114_32;
	wire [WIDTH*2-1+0:0] tmp00_114_33;
	wire [WIDTH*2-1+0:0] tmp00_114_34;
	wire [WIDTH*2-1+0:0] tmp00_114_35;
	wire [WIDTH*2-1+0:0] tmp00_114_36;
	wire [WIDTH*2-1+0:0] tmp00_114_37;
	wire [WIDTH*2-1+0:0] tmp00_114_38;
	wire [WIDTH*2-1+0:0] tmp00_114_39;
	wire [WIDTH*2-1+0:0] tmp00_114_40;
	wire [WIDTH*2-1+0:0] tmp00_114_41;
	wire [WIDTH*2-1+0:0] tmp00_114_42;
	wire [WIDTH*2-1+0:0] tmp00_114_43;
	wire [WIDTH*2-1+0:0] tmp00_114_44;
	wire [WIDTH*2-1+0:0] tmp00_114_45;
	wire [WIDTH*2-1+0:0] tmp00_114_46;
	wire [WIDTH*2-1+0:0] tmp00_114_47;
	wire [WIDTH*2-1+0:0] tmp00_114_48;
	wire [WIDTH*2-1+0:0] tmp00_114_49;
	wire [WIDTH*2-1+0:0] tmp00_114_50;
	wire [WIDTH*2-1+0:0] tmp00_114_51;
	wire [WIDTH*2-1+0:0] tmp00_114_52;
	wire [WIDTH*2-1+0:0] tmp00_114_53;
	wire [WIDTH*2-1+0:0] tmp00_114_54;
	wire [WIDTH*2-1+0:0] tmp00_114_55;
	wire [WIDTH*2-1+0:0] tmp00_114_56;
	wire [WIDTH*2-1+0:0] tmp00_114_57;
	wire [WIDTH*2-1+0:0] tmp00_114_58;
	wire [WIDTH*2-1+0:0] tmp00_114_59;
	wire [WIDTH*2-1+0:0] tmp00_114_60;
	wire [WIDTH*2-1+0:0] tmp00_114_61;
	wire [WIDTH*2-1+0:0] tmp00_114_62;
	wire [WIDTH*2-1+0:0] tmp00_114_63;
	wire [WIDTH*2-1+0:0] tmp00_114_64;
	wire [WIDTH*2-1+0:0] tmp00_114_65;
	wire [WIDTH*2-1+0:0] tmp00_114_66;
	wire [WIDTH*2-1+0:0] tmp00_114_67;
	wire [WIDTH*2-1+0:0] tmp00_114_68;
	wire [WIDTH*2-1+0:0] tmp00_114_69;
	wire [WIDTH*2-1+0:0] tmp00_114_70;
	wire [WIDTH*2-1+0:0] tmp00_114_71;
	wire [WIDTH*2-1+0:0] tmp00_114_72;
	wire [WIDTH*2-1+0:0] tmp00_114_73;
	wire [WIDTH*2-1+0:0] tmp00_114_74;
	wire [WIDTH*2-1+0:0] tmp00_114_75;
	wire [WIDTH*2-1+0:0] tmp00_114_76;
	wire [WIDTH*2-1+0:0] tmp00_114_77;
	wire [WIDTH*2-1+0:0] tmp00_114_78;
	wire [WIDTH*2-1+0:0] tmp00_114_79;
	wire [WIDTH*2-1+0:0] tmp00_114_80;
	wire [WIDTH*2-1+0:0] tmp00_114_81;
	wire [WIDTH*2-1+0:0] tmp00_114_82;
	wire [WIDTH*2-1+0:0] tmp00_114_83;
	wire [WIDTH*2-1+0:0] tmp00_115_0;
	wire [WIDTH*2-1+0:0] tmp00_115_1;
	wire [WIDTH*2-1+0:0] tmp00_115_2;
	wire [WIDTH*2-1+0:0] tmp00_115_3;
	wire [WIDTH*2-1+0:0] tmp00_115_4;
	wire [WIDTH*2-1+0:0] tmp00_115_5;
	wire [WIDTH*2-1+0:0] tmp00_115_6;
	wire [WIDTH*2-1+0:0] tmp00_115_7;
	wire [WIDTH*2-1+0:0] tmp00_115_8;
	wire [WIDTH*2-1+0:0] tmp00_115_9;
	wire [WIDTH*2-1+0:0] tmp00_115_10;
	wire [WIDTH*2-1+0:0] tmp00_115_11;
	wire [WIDTH*2-1+0:0] tmp00_115_12;
	wire [WIDTH*2-1+0:0] tmp00_115_13;
	wire [WIDTH*2-1+0:0] tmp00_115_14;
	wire [WIDTH*2-1+0:0] tmp00_115_15;
	wire [WIDTH*2-1+0:0] tmp00_115_16;
	wire [WIDTH*2-1+0:0] tmp00_115_17;
	wire [WIDTH*2-1+0:0] tmp00_115_18;
	wire [WIDTH*2-1+0:0] tmp00_115_19;
	wire [WIDTH*2-1+0:0] tmp00_115_20;
	wire [WIDTH*2-1+0:0] tmp00_115_21;
	wire [WIDTH*2-1+0:0] tmp00_115_22;
	wire [WIDTH*2-1+0:0] tmp00_115_23;
	wire [WIDTH*2-1+0:0] tmp00_115_24;
	wire [WIDTH*2-1+0:0] tmp00_115_25;
	wire [WIDTH*2-1+0:0] tmp00_115_26;
	wire [WIDTH*2-1+0:0] tmp00_115_27;
	wire [WIDTH*2-1+0:0] tmp00_115_28;
	wire [WIDTH*2-1+0:0] tmp00_115_29;
	wire [WIDTH*2-1+0:0] tmp00_115_30;
	wire [WIDTH*2-1+0:0] tmp00_115_31;
	wire [WIDTH*2-1+0:0] tmp00_115_32;
	wire [WIDTH*2-1+0:0] tmp00_115_33;
	wire [WIDTH*2-1+0:0] tmp00_115_34;
	wire [WIDTH*2-1+0:0] tmp00_115_35;
	wire [WIDTH*2-1+0:0] tmp00_115_36;
	wire [WIDTH*2-1+0:0] tmp00_115_37;
	wire [WIDTH*2-1+0:0] tmp00_115_38;
	wire [WIDTH*2-1+0:0] tmp00_115_39;
	wire [WIDTH*2-1+0:0] tmp00_115_40;
	wire [WIDTH*2-1+0:0] tmp00_115_41;
	wire [WIDTH*2-1+0:0] tmp00_115_42;
	wire [WIDTH*2-1+0:0] tmp00_115_43;
	wire [WIDTH*2-1+0:0] tmp00_115_44;
	wire [WIDTH*2-1+0:0] tmp00_115_45;
	wire [WIDTH*2-1+0:0] tmp00_115_46;
	wire [WIDTH*2-1+0:0] tmp00_115_47;
	wire [WIDTH*2-1+0:0] tmp00_115_48;
	wire [WIDTH*2-1+0:0] tmp00_115_49;
	wire [WIDTH*2-1+0:0] tmp00_115_50;
	wire [WIDTH*2-1+0:0] tmp00_115_51;
	wire [WIDTH*2-1+0:0] tmp00_115_52;
	wire [WIDTH*2-1+0:0] tmp00_115_53;
	wire [WIDTH*2-1+0:0] tmp00_115_54;
	wire [WIDTH*2-1+0:0] tmp00_115_55;
	wire [WIDTH*2-1+0:0] tmp00_115_56;
	wire [WIDTH*2-1+0:0] tmp00_115_57;
	wire [WIDTH*2-1+0:0] tmp00_115_58;
	wire [WIDTH*2-1+0:0] tmp00_115_59;
	wire [WIDTH*2-1+0:0] tmp00_115_60;
	wire [WIDTH*2-1+0:0] tmp00_115_61;
	wire [WIDTH*2-1+0:0] tmp00_115_62;
	wire [WIDTH*2-1+0:0] tmp00_115_63;
	wire [WIDTH*2-1+0:0] tmp00_115_64;
	wire [WIDTH*2-1+0:0] tmp00_115_65;
	wire [WIDTH*2-1+0:0] tmp00_115_66;
	wire [WIDTH*2-1+0:0] tmp00_115_67;
	wire [WIDTH*2-1+0:0] tmp00_115_68;
	wire [WIDTH*2-1+0:0] tmp00_115_69;
	wire [WIDTH*2-1+0:0] tmp00_115_70;
	wire [WIDTH*2-1+0:0] tmp00_115_71;
	wire [WIDTH*2-1+0:0] tmp00_115_72;
	wire [WIDTH*2-1+0:0] tmp00_115_73;
	wire [WIDTH*2-1+0:0] tmp00_115_74;
	wire [WIDTH*2-1+0:0] tmp00_115_75;
	wire [WIDTH*2-1+0:0] tmp00_115_76;
	wire [WIDTH*2-1+0:0] tmp00_115_77;
	wire [WIDTH*2-1+0:0] tmp00_115_78;
	wire [WIDTH*2-1+0:0] tmp00_115_79;
	wire [WIDTH*2-1+0:0] tmp00_115_80;
	wire [WIDTH*2-1+0:0] tmp00_115_81;
	wire [WIDTH*2-1+0:0] tmp00_115_82;
	wire [WIDTH*2-1+0:0] tmp00_115_83;
	wire [WIDTH*2-1+0:0] tmp00_116_0;
	wire [WIDTH*2-1+0:0] tmp00_116_1;
	wire [WIDTH*2-1+0:0] tmp00_116_2;
	wire [WIDTH*2-1+0:0] tmp00_116_3;
	wire [WIDTH*2-1+0:0] tmp00_116_4;
	wire [WIDTH*2-1+0:0] tmp00_116_5;
	wire [WIDTH*2-1+0:0] tmp00_116_6;
	wire [WIDTH*2-1+0:0] tmp00_116_7;
	wire [WIDTH*2-1+0:0] tmp00_116_8;
	wire [WIDTH*2-1+0:0] tmp00_116_9;
	wire [WIDTH*2-1+0:0] tmp00_116_10;
	wire [WIDTH*2-1+0:0] tmp00_116_11;
	wire [WIDTH*2-1+0:0] tmp00_116_12;
	wire [WIDTH*2-1+0:0] tmp00_116_13;
	wire [WIDTH*2-1+0:0] tmp00_116_14;
	wire [WIDTH*2-1+0:0] tmp00_116_15;
	wire [WIDTH*2-1+0:0] tmp00_116_16;
	wire [WIDTH*2-1+0:0] tmp00_116_17;
	wire [WIDTH*2-1+0:0] tmp00_116_18;
	wire [WIDTH*2-1+0:0] tmp00_116_19;
	wire [WIDTH*2-1+0:0] tmp00_116_20;
	wire [WIDTH*2-1+0:0] tmp00_116_21;
	wire [WIDTH*2-1+0:0] tmp00_116_22;
	wire [WIDTH*2-1+0:0] tmp00_116_23;
	wire [WIDTH*2-1+0:0] tmp00_116_24;
	wire [WIDTH*2-1+0:0] tmp00_116_25;
	wire [WIDTH*2-1+0:0] tmp00_116_26;
	wire [WIDTH*2-1+0:0] tmp00_116_27;
	wire [WIDTH*2-1+0:0] tmp00_116_28;
	wire [WIDTH*2-1+0:0] tmp00_116_29;
	wire [WIDTH*2-1+0:0] tmp00_116_30;
	wire [WIDTH*2-1+0:0] tmp00_116_31;
	wire [WIDTH*2-1+0:0] tmp00_116_32;
	wire [WIDTH*2-1+0:0] tmp00_116_33;
	wire [WIDTH*2-1+0:0] tmp00_116_34;
	wire [WIDTH*2-1+0:0] tmp00_116_35;
	wire [WIDTH*2-1+0:0] tmp00_116_36;
	wire [WIDTH*2-1+0:0] tmp00_116_37;
	wire [WIDTH*2-1+0:0] tmp00_116_38;
	wire [WIDTH*2-1+0:0] tmp00_116_39;
	wire [WIDTH*2-1+0:0] tmp00_116_40;
	wire [WIDTH*2-1+0:0] tmp00_116_41;
	wire [WIDTH*2-1+0:0] tmp00_116_42;
	wire [WIDTH*2-1+0:0] tmp00_116_43;
	wire [WIDTH*2-1+0:0] tmp00_116_44;
	wire [WIDTH*2-1+0:0] tmp00_116_45;
	wire [WIDTH*2-1+0:0] tmp00_116_46;
	wire [WIDTH*2-1+0:0] tmp00_116_47;
	wire [WIDTH*2-1+0:0] tmp00_116_48;
	wire [WIDTH*2-1+0:0] tmp00_116_49;
	wire [WIDTH*2-1+0:0] tmp00_116_50;
	wire [WIDTH*2-1+0:0] tmp00_116_51;
	wire [WIDTH*2-1+0:0] tmp00_116_52;
	wire [WIDTH*2-1+0:0] tmp00_116_53;
	wire [WIDTH*2-1+0:0] tmp00_116_54;
	wire [WIDTH*2-1+0:0] tmp00_116_55;
	wire [WIDTH*2-1+0:0] tmp00_116_56;
	wire [WIDTH*2-1+0:0] tmp00_116_57;
	wire [WIDTH*2-1+0:0] tmp00_116_58;
	wire [WIDTH*2-1+0:0] tmp00_116_59;
	wire [WIDTH*2-1+0:0] tmp00_116_60;
	wire [WIDTH*2-1+0:0] tmp00_116_61;
	wire [WIDTH*2-1+0:0] tmp00_116_62;
	wire [WIDTH*2-1+0:0] tmp00_116_63;
	wire [WIDTH*2-1+0:0] tmp00_116_64;
	wire [WIDTH*2-1+0:0] tmp00_116_65;
	wire [WIDTH*2-1+0:0] tmp00_116_66;
	wire [WIDTH*2-1+0:0] tmp00_116_67;
	wire [WIDTH*2-1+0:0] tmp00_116_68;
	wire [WIDTH*2-1+0:0] tmp00_116_69;
	wire [WIDTH*2-1+0:0] tmp00_116_70;
	wire [WIDTH*2-1+0:0] tmp00_116_71;
	wire [WIDTH*2-1+0:0] tmp00_116_72;
	wire [WIDTH*2-1+0:0] tmp00_116_73;
	wire [WIDTH*2-1+0:0] tmp00_116_74;
	wire [WIDTH*2-1+0:0] tmp00_116_75;
	wire [WIDTH*2-1+0:0] tmp00_116_76;
	wire [WIDTH*2-1+0:0] tmp00_116_77;
	wire [WIDTH*2-1+0:0] tmp00_116_78;
	wire [WIDTH*2-1+0:0] tmp00_116_79;
	wire [WIDTH*2-1+0:0] tmp00_116_80;
	wire [WIDTH*2-1+0:0] tmp00_116_81;
	wire [WIDTH*2-1+0:0] tmp00_116_82;
	wire [WIDTH*2-1+0:0] tmp00_116_83;
	wire [WIDTH*2-1+0:0] tmp00_117_0;
	wire [WIDTH*2-1+0:0] tmp00_117_1;
	wire [WIDTH*2-1+0:0] tmp00_117_2;
	wire [WIDTH*2-1+0:0] tmp00_117_3;
	wire [WIDTH*2-1+0:0] tmp00_117_4;
	wire [WIDTH*2-1+0:0] tmp00_117_5;
	wire [WIDTH*2-1+0:0] tmp00_117_6;
	wire [WIDTH*2-1+0:0] tmp00_117_7;
	wire [WIDTH*2-1+0:0] tmp00_117_8;
	wire [WIDTH*2-1+0:0] tmp00_117_9;
	wire [WIDTH*2-1+0:0] tmp00_117_10;
	wire [WIDTH*2-1+0:0] tmp00_117_11;
	wire [WIDTH*2-1+0:0] tmp00_117_12;
	wire [WIDTH*2-1+0:0] tmp00_117_13;
	wire [WIDTH*2-1+0:0] tmp00_117_14;
	wire [WIDTH*2-1+0:0] tmp00_117_15;
	wire [WIDTH*2-1+0:0] tmp00_117_16;
	wire [WIDTH*2-1+0:0] tmp00_117_17;
	wire [WIDTH*2-1+0:0] tmp00_117_18;
	wire [WIDTH*2-1+0:0] tmp00_117_19;
	wire [WIDTH*2-1+0:0] tmp00_117_20;
	wire [WIDTH*2-1+0:0] tmp00_117_21;
	wire [WIDTH*2-1+0:0] tmp00_117_22;
	wire [WIDTH*2-1+0:0] tmp00_117_23;
	wire [WIDTH*2-1+0:0] tmp00_117_24;
	wire [WIDTH*2-1+0:0] tmp00_117_25;
	wire [WIDTH*2-1+0:0] tmp00_117_26;
	wire [WIDTH*2-1+0:0] tmp00_117_27;
	wire [WIDTH*2-1+0:0] tmp00_117_28;
	wire [WIDTH*2-1+0:0] tmp00_117_29;
	wire [WIDTH*2-1+0:0] tmp00_117_30;
	wire [WIDTH*2-1+0:0] tmp00_117_31;
	wire [WIDTH*2-1+0:0] tmp00_117_32;
	wire [WIDTH*2-1+0:0] tmp00_117_33;
	wire [WIDTH*2-1+0:0] tmp00_117_34;
	wire [WIDTH*2-1+0:0] tmp00_117_35;
	wire [WIDTH*2-1+0:0] tmp00_117_36;
	wire [WIDTH*2-1+0:0] tmp00_117_37;
	wire [WIDTH*2-1+0:0] tmp00_117_38;
	wire [WIDTH*2-1+0:0] tmp00_117_39;
	wire [WIDTH*2-1+0:0] tmp00_117_40;
	wire [WIDTH*2-1+0:0] tmp00_117_41;
	wire [WIDTH*2-1+0:0] tmp00_117_42;
	wire [WIDTH*2-1+0:0] tmp00_117_43;
	wire [WIDTH*2-1+0:0] tmp00_117_44;
	wire [WIDTH*2-1+0:0] tmp00_117_45;
	wire [WIDTH*2-1+0:0] tmp00_117_46;
	wire [WIDTH*2-1+0:0] tmp00_117_47;
	wire [WIDTH*2-1+0:0] tmp00_117_48;
	wire [WIDTH*2-1+0:0] tmp00_117_49;
	wire [WIDTH*2-1+0:0] tmp00_117_50;
	wire [WIDTH*2-1+0:0] tmp00_117_51;
	wire [WIDTH*2-1+0:0] tmp00_117_52;
	wire [WIDTH*2-1+0:0] tmp00_117_53;
	wire [WIDTH*2-1+0:0] tmp00_117_54;
	wire [WIDTH*2-1+0:0] tmp00_117_55;
	wire [WIDTH*2-1+0:0] tmp00_117_56;
	wire [WIDTH*2-1+0:0] tmp00_117_57;
	wire [WIDTH*2-1+0:0] tmp00_117_58;
	wire [WIDTH*2-1+0:0] tmp00_117_59;
	wire [WIDTH*2-1+0:0] tmp00_117_60;
	wire [WIDTH*2-1+0:0] tmp00_117_61;
	wire [WIDTH*2-1+0:0] tmp00_117_62;
	wire [WIDTH*2-1+0:0] tmp00_117_63;
	wire [WIDTH*2-1+0:0] tmp00_117_64;
	wire [WIDTH*2-1+0:0] tmp00_117_65;
	wire [WIDTH*2-1+0:0] tmp00_117_66;
	wire [WIDTH*2-1+0:0] tmp00_117_67;
	wire [WIDTH*2-1+0:0] tmp00_117_68;
	wire [WIDTH*2-1+0:0] tmp00_117_69;
	wire [WIDTH*2-1+0:0] tmp00_117_70;
	wire [WIDTH*2-1+0:0] tmp00_117_71;
	wire [WIDTH*2-1+0:0] tmp00_117_72;
	wire [WIDTH*2-1+0:0] tmp00_117_73;
	wire [WIDTH*2-1+0:0] tmp00_117_74;
	wire [WIDTH*2-1+0:0] tmp00_117_75;
	wire [WIDTH*2-1+0:0] tmp00_117_76;
	wire [WIDTH*2-1+0:0] tmp00_117_77;
	wire [WIDTH*2-1+0:0] tmp00_117_78;
	wire [WIDTH*2-1+0:0] tmp00_117_79;
	wire [WIDTH*2-1+0:0] tmp00_117_80;
	wire [WIDTH*2-1+0:0] tmp00_117_81;
	wire [WIDTH*2-1+0:0] tmp00_117_82;
	wire [WIDTH*2-1+0:0] tmp00_117_83;
	wire [WIDTH*2-1+0:0] tmp00_118_0;
	wire [WIDTH*2-1+0:0] tmp00_118_1;
	wire [WIDTH*2-1+0:0] tmp00_118_2;
	wire [WIDTH*2-1+0:0] tmp00_118_3;
	wire [WIDTH*2-1+0:0] tmp00_118_4;
	wire [WIDTH*2-1+0:0] tmp00_118_5;
	wire [WIDTH*2-1+0:0] tmp00_118_6;
	wire [WIDTH*2-1+0:0] tmp00_118_7;
	wire [WIDTH*2-1+0:0] tmp00_118_8;
	wire [WIDTH*2-1+0:0] tmp00_118_9;
	wire [WIDTH*2-1+0:0] tmp00_118_10;
	wire [WIDTH*2-1+0:0] tmp00_118_11;
	wire [WIDTH*2-1+0:0] tmp00_118_12;
	wire [WIDTH*2-1+0:0] tmp00_118_13;
	wire [WIDTH*2-1+0:0] tmp00_118_14;
	wire [WIDTH*2-1+0:0] tmp00_118_15;
	wire [WIDTH*2-1+0:0] tmp00_118_16;
	wire [WIDTH*2-1+0:0] tmp00_118_17;
	wire [WIDTH*2-1+0:0] tmp00_118_18;
	wire [WIDTH*2-1+0:0] tmp00_118_19;
	wire [WIDTH*2-1+0:0] tmp00_118_20;
	wire [WIDTH*2-1+0:0] tmp00_118_21;
	wire [WIDTH*2-1+0:0] tmp00_118_22;
	wire [WIDTH*2-1+0:0] tmp00_118_23;
	wire [WIDTH*2-1+0:0] tmp00_118_24;
	wire [WIDTH*2-1+0:0] tmp00_118_25;
	wire [WIDTH*2-1+0:0] tmp00_118_26;
	wire [WIDTH*2-1+0:0] tmp00_118_27;
	wire [WIDTH*2-1+0:0] tmp00_118_28;
	wire [WIDTH*2-1+0:0] tmp00_118_29;
	wire [WIDTH*2-1+0:0] tmp00_118_30;
	wire [WIDTH*2-1+0:0] tmp00_118_31;
	wire [WIDTH*2-1+0:0] tmp00_118_32;
	wire [WIDTH*2-1+0:0] tmp00_118_33;
	wire [WIDTH*2-1+0:0] tmp00_118_34;
	wire [WIDTH*2-1+0:0] tmp00_118_35;
	wire [WIDTH*2-1+0:0] tmp00_118_36;
	wire [WIDTH*2-1+0:0] tmp00_118_37;
	wire [WIDTH*2-1+0:0] tmp00_118_38;
	wire [WIDTH*2-1+0:0] tmp00_118_39;
	wire [WIDTH*2-1+0:0] tmp00_118_40;
	wire [WIDTH*2-1+0:0] tmp00_118_41;
	wire [WIDTH*2-1+0:0] tmp00_118_42;
	wire [WIDTH*2-1+0:0] tmp00_118_43;
	wire [WIDTH*2-1+0:0] tmp00_118_44;
	wire [WIDTH*2-1+0:0] tmp00_118_45;
	wire [WIDTH*2-1+0:0] tmp00_118_46;
	wire [WIDTH*2-1+0:0] tmp00_118_47;
	wire [WIDTH*2-1+0:0] tmp00_118_48;
	wire [WIDTH*2-1+0:0] tmp00_118_49;
	wire [WIDTH*2-1+0:0] tmp00_118_50;
	wire [WIDTH*2-1+0:0] tmp00_118_51;
	wire [WIDTH*2-1+0:0] tmp00_118_52;
	wire [WIDTH*2-1+0:0] tmp00_118_53;
	wire [WIDTH*2-1+0:0] tmp00_118_54;
	wire [WIDTH*2-1+0:0] tmp00_118_55;
	wire [WIDTH*2-1+0:0] tmp00_118_56;
	wire [WIDTH*2-1+0:0] tmp00_118_57;
	wire [WIDTH*2-1+0:0] tmp00_118_58;
	wire [WIDTH*2-1+0:0] tmp00_118_59;
	wire [WIDTH*2-1+0:0] tmp00_118_60;
	wire [WIDTH*2-1+0:0] tmp00_118_61;
	wire [WIDTH*2-1+0:0] tmp00_118_62;
	wire [WIDTH*2-1+0:0] tmp00_118_63;
	wire [WIDTH*2-1+0:0] tmp00_118_64;
	wire [WIDTH*2-1+0:0] tmp00_118_65;
	wire [WIDTH*2-1+0:0] tmp00_118_66;
	wire [WIDTH*2-1+0:0] tmp00_118_67;
	wire [WIDTH*2-1+0:0] tmp00_118_68;
	wire [WIDTH*2-1+0:0] tmp00_118_69;
	wire [WIDTH*2-1+0:0] tmp00_118_70;
	wire [WIDTH*2-1+0:0] tmp00_118_71;
	wire [WIDTH*2-1+0:0] tmp00_118_72;
	wire [WIDTH*2-1+0:0] tmp00_118_73;
	wire [WIDTH*2-1+0:0] tmp00_118_74;
	wire [WIDTH*2-1+0:0] tmp00_118_75;
	wire [WIDTH*2-1+0:0] tmp00_118_76;
	wire [WIDTH*2-1+0:0] tmp00_118_77;
	wire [WIDTH*2-1+0:0] tmp00_118_78;
	wire [WIDTH*2-1+0:0] tmp00_118_79;
	wire [WIDTH*2-1+0:0] tmp00_118_80;
	wire [WIDTH*2-1+0:0] tmp00_118_81;
	wire [WIDTH*2-1+0:0] tmp00_118_82;
	wire [WIDTH*2-1+0:0] tmp00_118_83;
	wire [WIDTH*2-1+0:0] tmp00_119_0;
	wire [WIDTH*2-1+0:0] tmp00_119_1;
	wire [WIDTH*2-1+0:0] tmp00_119_2;
	wire [WIDTH*2-1+0:0] tmp00_119_3;
	wire [WIDTH*2-1+0:0] tmp00_119_4;
	wire [WIDTH*2-1+0:0] tmp00_119_5;
	wire [WIDTH*2-1+0:0] tmp00_119_6;
	wire [WIDTH*2-1+0:0] tmp00_119_7;
	wire [WIDTH*2-1+0:0] tmp00_119_8;
	wire [WIDTH*2-1+0:0] tmp00_119_9;
	wire [WIDTH*2-1+0:0] tmp00_119_10;
	wire [WIDTH*2-1+0:0] tmp00_119_11;
	wire [WIDTH*2-1+0:0] tmp00_119_12;
	wire [WIDTH*2-1+0:0] tmp00_119_13;
	wire [WIDTH*2-1+0:0] tmp00_119_14;
	wire [WIDTH*2-1+0:0] tmp00_119_15;
	wire [WIDTH*2-1+0:0] tmp00_119_16;
	wire [WIDTH*2-1+0:0] tmp00_119_17;
	wire [WIDTH*2-1+0:0] tmp00_119_18;
	wire [WIDTH*2-1+0:0] tmp00_119_19;
	wire [WIDTH*2-1+0:0] tmp00_119_20;
	wire [WIDTH*2-1+0:0] tmp00_119_21;
	wire [WIDTH*2-1+0:0] tmp00_119_22;
	wire [WIDTH*2-1+0:0] tmp00_119_23;
	wire [WIDTH*2-1+0:0] tmp00_119_24;
	wire [WIDTH*2-1+0:0] tmp00_119_25;
	wire [WIDTH*2-1+0:0] tmp00_119_26;
	wire [WIDTH*2-1+0:0] tmp00_119_27;
	wire [WIDTH*2-1+0:0] tmp00_119_28;
	wire [WIDTH*2-1+0:0] tmp00_119_29;
	wire [WIDTH*2-1+0:0] tmp00_119_30;
	wire [WIDTH*2-1+0:0] tmp00_119_31;
	wire [WIDTH*2-1+0:0] tmp00_119_32;
	wire [WIDTH*2-1+0:0] tmp00_119_33;
	wire [WIDTH*2-1+0:0] tmp00_119_34;
	wire [WIDTH*2-1+0:0] tmp00_119_35;
	wire [WIDTH*2-1+0:0] tmp00_119_36;
	wire [WIDTH*2-1+0:0] tmp00_119_37;
	wire [WIDTH*2-1+0:0] tmp00_119_38;
	wire [WIDTH*2-1+0:0] tmp00_119_39;
	wire [WIDTH*2-1+0:0] tmp00_119_40;
	wire [WIDTH*2-1+0:0] tmp00_119_41;
	wire [WIDTH*2-1+0:0] tmp00_119_42;
	wire [WIDTH*2-1+0:0] tmp00_119_43;
	wire [WIDTH*2-1+0:0] tmp00_119_44;
	wire [WIDTH*2-1+0:0] tmp00_119_45;
	wire [WIDTH*2-1+0:0] tmp00_119_46;
	wire [WIDTH*2-1+0:0] tmp00_119_47;
	wire [WIDTH*2-1+0:0] tmp00_119_48;
	wire [WIDTH*2-1+0:0] tmp00_119_49;
	wire [WIDTH*2-1+0:0] tmp00_119_50;
	wire [WIDTH*2-1+0:0] tmp00_119_51;
	wire [WIDTH*2-1+0:0] tmp00_119_52;
	wire [WIDTH*2-1+0:0] tmp00_119_53;
	wire [WIDTH*2-1+0:0] tmp00_119_54;
	wire [WIDTH*2-1+0:0] tmp00_119_55;
	wire [WIDTH*2-1+0:0] tmp00_119_56;
	wire [WIDTH*2-1+0:0] tmp00_119_57;
	wire [WIDTH*2-1+0:0] tmp00_119_58;
	wire [WIDTH*2-1+0:0] tmp00_119_59;
	wire [WIDTH*2-1+0:0] tmp00_119_60;
	wire [WIDTH*2-1+0:0] tmp00_119_61;
	wire [WIDTH*2-1+0:0] tmp00_119_62;
	wire [WIDTH*2-1+0:0] tmp00_119_63;
	wire [WIDTH*2-1+0:0] tmp00_119_64;
	wire [WIDTH*2-1+0:0] tmp00_119_65;
	wire [WIDTH*2-1+0:0] tmp00_119_66;
	wire [WIDTH*2-1+0:0] tmp00_119_67;
	wire [WIDTH*2-1+0:0] tmp00_119_68;
	wire [WIDTH*2-1+0:0] tmp00_119_69;
	wire [WIDTH*2-1+0:0] tmp00_119_70;
	wire [WIDTH*2-1+0:0] tmp00_119_71;
	wire [WIDTH*2-1+0:0] tmp00_119_72;
	wire [WIDTH*2-1+0:0] tmp00_119_73;
	wire [WIDTH*2-1+0:0] tmp00_119_74;
	wire [WIDTH*2-1+0:0] tmp00_119_75;
	wire [WIDTH*2-1+0:0] tmp00_119_76;
	wire [WIDTH*2-1+0:0] tmp00_119_77;
	wire [WIDTH*2-1+0:0] tmp00_119_78;
	wire [WIDTH*2-1+0:0] tmp00_119_79;
	wire [WIDTH*2-1+0:0] tmp00_119_80;
	wire [WIDTH*2-1+0:0] tmp00_119_81;
	wire [WIDTH*2-1+0:0] tmp00_119_82;
	wire [WIDTH*2-1+0:0] tmp00_119_83;
	wire [WIDTH*2-1+0:0] tmp00_120_0;
	wire [WIDTH*2-1+0:0] tmp00_120_1;
	wire [WIDTH*2-1+0:0] tmp00_120_2;
	wire [WIDTH*2-1+0:0] tmp00_120_3;
	wire [WIDTH*2-1+0:0] tmp00_120_4;
	wire [WIDTH*2-1+0:0] tmp00_120_5;
	wire [WIDTH*2-1+0:0] tmp00_120_6;
	wire [WIDTH*2-1+0:0] tmp00_120_7;
	wire [WIDTH*2-1+0:0] tmp00_120_8;
	wire [WIDTH*2-1+0:0] tmp00_120_9;
	wire [WIDTH*2-1+0:0] tmp00_120_10;
	wire [WIDTH*2-1+0:0] tmp00_120_11;
	wire [WIDTH*2-1+0:0] tmp00_120_12;
	wire [WIDTH*2-1+0:0] tmp00_120_13;
	wire [WIDTH*2-1+0:0] tmp00_120_14;
	wire [WIDTH*2-1+0:0] tmp00_120_15;
	wire [WIDTH*2-1+0:0] tmp00_120_16;
	wire [WIDTH*2-1+0:0] tmp00_120_17;
	wire [WIDTH*2-1+0:0] tmp00_120_18;
	wire [WIDTH*2-1+0:0] tmp00_120_19;
	wire [WIDTH*2-1+0:0] tmp00_120_20;
	wire [WIDTH*2-1+0:0] tmp00_120_21;
	wire [WIDTH*2-1+0:0] tmp00_120_22;
	wire [WIDTH*2-1+0:0] tmp00_120_23;
	wire [WIDTH*2-1+0:0] tmp00_120_24;
	wire [WIDTH*2-1+0:0] tmp00_120_25;
	wire [WIDTH*2-1+0:0] tmp00_120_26;
	wire [WIDTH*2-1+0:0] tmp00_120_27;
	wire [WIDTH*2-1+0:0] tmp00_120_28;
	wire [WIDTH*2-1+0:0] tmp00_120_29;
	wire [WIDTH*2-1+0:0] tmp00_120_30;
	wire [WIDTH*2-1+0:0] tmp00_120_31;
	wire [WIDTH*2-1+0:0] tmp00_120_32;
	wire [WIDTH*2-1+0:0] tmp00_120_33;
	wire [WIDTH*2-1+0:0] tmp00_120_34;
	wire [WIDTH*2-1+0:0] tmp00_120_35;
	wire [WIDTH*2-1+0:0] tmp00_120_36;
	wire [WIDTH*2-1+0:0] tmp00_120_37;
	wire [WIDTH*2-1+0:0] tmp00_120_38;
	wire [WIDTH*2-1+0:0] tmp00_120_39;
	wire [WIDTH*2-1+0:0] tmp00_120_40;
	wire [WIDTH*2-1+0:0] tmp00_120_41;
	wire [WIDTH*2-1+0:0] tmp00_120_42;
	wire [WIDTH*2-1+0:0] tmp00_120_43;
	wire [WIDTH*2-1+0:0] tmp00_120_44;
	wire [WIDTH*2-1+0:0] tmp00_120_45;
	wire [WIDTH*2-1+0:0] tmp00_120_46;
	wire [WIDTH*2-1+0:0] tmp00_120_47;
	wire [WIDTH*2-1+0:0] tmp00_120_48;
	wire [WIDTH*2-1+0:0] tmp00_120_49;
	wire [WIDTH*2-1+0:0] tmp00_120_50;
	wire [WIDTH*2-1+0:0] tmp00_120_51;
	wire [WIDTH*2-1+0:0] tmp00_120_52;
	wire [WIDTH*2-1+0:0] tmp00_120_53;
	wire [WIDTH*2-1+0:0] tmp00_120_54;
	wire [WIDTH*2-1+0:0] tmp00_120_55;
	wire [WIDTH*2-1+0:0] tmp00_120_56;
	wire [WIDTH*2-1+0:0] tmp00_120_57;
	wire [WIDTH*2-1+0:0] tmp00_120_58;
	wire [WIDTH*2-1+0:0] tmp00_120_59;
	wire [WIDTH*2-1+0:0] tmp00_120_60;
	wire [WIDTH*2-1+0:0] tmp00_120_61;
	wire [WIDTH*2-1+0:0] tmp00_120_62;
	wire [WIDTH*2-1+0:0] tmp00_120_63;
	wire [WIDTH*2-1+0:0] tmp00_120_64;
	wire [WIDTH*2-1+0:0] tmp00_120_65;
	wire [WIDTH*2-1+0:0] tmp00_120_66;
	wire [WIDTH*2-1+0:0] tmp00_120_67;
	wire [WIDTH*2-1+0:0] tmp00_120_68;
	wire [WIDTH*2-1+0:0] tmp00_120_69;
	wire [WIDTH*2-1+0:0] tmp00_120_70;
	wire [WIDTH*2-1+0:0] tmp00_120_71;
	wire [WIDTH*2-1+0:0] tmp00_120_72;
	wire [WIDTH*2-1+0:0] tmp00_120_73;
	wire [WIDTH*2-1+0:0] tmp00_120_74;
	wire [WIDTH*2-1+0:0] tmp00_120_75;
	wire [WIDTH*2-1+0:0] tmp00_120_76;
	wire [WIDTH*2-1+0:0] tmp00_120_77;
	wire [WIDTH*2-1+0:0] tmp00_120_78;
	wire [WIDTH*2-1+0:0] tmp00_120_79;
	wire [WIDTH*2-1+0:0] tmp00_120_80;
	wire [WIDTH*2-1+0:0] tmp00_120_81;
	wire [WIDTH*2-1+0:0] tmp00_120_82;
	wire [WIDTH*2-1+0:0] tmp00_120_83;
	wire [WIDTH*2-1+0:0] tmp00_121_0;
	wire [WIDTH*2-1+0:0] tmp00_121_1;
	wire [WIDTH*2-1+0:0] tmp00_121_2;
	wire [WIDTH*2-1+0:0] tmp00_121_3;
	wire [WIDTH*2-1+0:0] tmp00_121_4;
	wire [WIDTH*2-1+0:0] tmp00_121_5;
	wire [WIDTH*2-1+0:0] tmp00_121_6;
	wire [WIDTH*2-1+0:0] tmp00_121_7;
	wire [WIDTH*2-1+0:0] tmp00_121_8;
	wire [WIDTH*2-1+0:0] tmp00_121_9;
	wire [WIDTH*2-1+0:0] tmp00_121_10;
	wire [WIDTH*2-1+0:0] tmp00_121_11;
	wire [WIDTH*2-1+0:0] tmp00_121_12;
	wire [WIDTH*2-1+0:0] tmp00_121_13;
	wire [WIDTH*2-1+0:0] tmp00_121_14;
	wire [WIDTH*2-1+0:0] tmp00_121_15;
	wire [WIDTH*2-1+0:0] tmp00_121_16;
	wire [WIDTH*2-1+0:0] tmp00_121_17;
	wire [WIDTH*2-1+0:0] tmp00_121_18;
	wire [WIDTH*2-1+0:0] tmp00_121_19;
	wire [WIDTH*2-1+0:0] tmp00_121_20;
	wire [WIDTH*2-1+0:0] tmp00_121_21;
	wire [WIDTH*2-1+0:0] tmp00_121_22;
	wire [WIDTH*2-1+0:0] tmp00_121_23;
	wire [WIDTH*2-1+0:0] tmp00_121_24;
	wire [WIDTH*2-1+0:0] tmp00_121_25;
	wire [WIDTH*2-1+0:0] tmp00_121_26;
	wire [WIDTH*2-1+0:0] tmp00_121_27;
	wire [WIDTH*2-1+0:0] tmp00_121_28;
	wire [WIDTH*2-1+0:0] tmp00_121_29;
	wire [WIDTH*2-1+0:0] tmp00_121_30;
	wire [WIDTH*2-1+0:0] tmp00_121_31;
	wire [WIDTH*2-1+0:0] tmp00_121_32;
	wire [WIDTH*2-1+0:0] tmp00_121_33;
	wire [WIDTH*2-1+0:0] tmp00_121_34;
	wire [WIDTH*2-1+0:0] tmp00_121_35;
	wire [WIDTH*2-1+0:0] tmp00_121_36;
	wire [WIDTH*2-1+0:0] tmp00_121_37;
	wire [WIDTH*2-1+0:0] tmp00_121_38;
	wire [WIDTH*2-1+0:0] tmp00_121_39;
	wire [WIDTH*2-1+0:0] tmp00_121_40;
	wire [WIDTH*2-1+0:0] tmp00_121_41;
	wire [WIDTH*2-1+0:0] tmp00_121_42;
	wire [WIDTH*2-1+0:0] tmp00_121_43;
	wire [WIDTH*2-1+0:0] tmp00_121_44;
	wire [WIDTH*2-1+0:0] tmp00_121_45;
	wire [WIDTH*2-1+0:0] tmp00_121_46;
	wire [WIDTH*2-1+0:0] tmp00_121_47;
	wire [WIDTH*2-1+0:0] tmp00_121_48;
	wire [WIDTH*2-1+0:0] tmp00_121_49;
	wire [WIDTH*2-1+0:0] tmp00_121_50;
	wire [WIDTH*2-1+0:0] tmp00_121_51;
	wire [WIDTH*2-1+0:0] tmp00_121_52;
	wire [WIDTH*2-1+0:0] tmp00_121_53;
	wire [WIDTH*2-1+0:0] tmp00_121_54;
	wire [WIDTH*2-1+0:0] tmp00_121_55;
	wire [WIDTH*2-1+0:0] tmp00_121_56;
	wire [WIDTH*2-1+0:0] tmp00_121_57;
	wire [WIDTH*2-1+0:0] tmp00_121_58;
	wire [WIDTH*2-1+0:0] tmp00_121_59;
	wire [WIDTH*2-1+0:0] tmp00_121_60;
	wire [WIDTH*2-1+0:0] tmp00_121_61;
	wire [WIDTH*2-1+0:0] tmp00_121_62;
	wire [WIDTH*2-1+0:0] tmp00_121_63;
	wire [WIDTH*2-1+0:0] tmp00_121_64;
	wire [WIDTH*2-1+0:0] tmp00_121_65;
	wire [WIDTH*2-1+0:0] tmp00_121_66;
	wire [WIDTH*2-1+0:0] tmp00_121_67;
	wire [WIDTH*2-1+0:0] tmp00_121_68;
	wire [WIDTH*2-1+0:0] tmp00_121_69;
	wire [WIDTH*2-1+0:0] tmp00_121_70;
	wire [WIDTH*2-1+0:0] tmp00_121_71;
	wire [WIDTH*2-1+0:0] tmp00_121_72;
	wire [WIDTH*2-1+0:0] tmp00_121_73;
	wire [WIDTH*2-1+0:0] tmp00_121_74;
	wire [WIDTH*2-1+0:0] tmp00_121_75;
	wire [WIDTH*2-1+0:0] tmp00_121_76;
	wire [WIDTH*2-1+0:0] tmp00_121_77;
	wire [WIDTH*2-1+0:0] tmp00_121_78;
	wire [WIDTH*2-1+0:0] tmp00_121_79;
	wire [WIDTH*2-1+0:0] tmp00_121_80;
	wire [WIDTH*2-1+0:0] tmp00_121_81;
	wire [WIDTH*2-1+0:0] tmp00_121_82;
	wire [WIDTH*2-1+0:0] tmp00_121_83;
	wire [WIDTH*2-1+0:0] tmp00_122_0;
	wire [WIDTH*2-1+0:0] tmp00_122_1;
	wire [WIDTH*2-1+0:0] tmp00_122_2;
	wire [WIDTH*2-1+0:0] tmp00_122_3;
	wire [WIDTH*2-1+0:0] tmp00_122_4;
	wire [WIDTH*2-1+0:0] tmp00_122_5;
	wire [WIDTH*2-1+0:0] tmp00_122_6;
	wire [WIDTH*2-1+0:0] tmp00_122_7;
	wire [WIDTH*2-1+0:0] tmp00_122_8;
	wire [WIDTH*2-1+0:0] tmp00_122_9;
	wire [WIDTH*2-1+0:0] tmp00_122_10;
	wire [WIDTH*2-1+0:0] tmp00_122_11;
	wire [WIDTH*2-1+0:0] tmp00_122_12;
	wire [WIDTH*2-1+0:0] tmp00_122_13;
	wire [WIDTH*2-1+0:0] tmp00_122_14;
	wire [WIDTH*2-1+0:0] tmp00_122_15;
	wire [WIDTH*2-1+0:0] tmp00_122_16;
	wire [WIDTH*2-1+0:0] tmp00_122_17;
	wire [WIDTH*2-1+0:0] tmp00_122_18;
	wire [WIDTH*2-1+0:0] tmp00_122_19;
	wire [WIDTH*2-1+0:0] tmp00_122_20;
	wire [WIDTH*2-1+0:0] tmp00_122_21;
	wire [WIDTH*2-1+0:0] tmp00_122_22;
	wire [WIDTH*2-1+0:0] tmp00_122_23;
	wire [WIDTH*2-1+0:0] tmp00_122_24;
	wire [WIDTH*2-1+0:0] tmp00_122_25;
	wire [WIDTH*2-1+0:0] tmp00_122_26;
	wire [WIDTH*2-1+0:0] tmp00_122_27;
	wire [WIDTH*2-1+0:0] tmp00_122_28;
	wire [WIDTH*2-1+0:0] tmp00_122_29;
	wire [WIDTH*2-1+0:0] tmp00_122_30;
	wire [WIDTH*2-1+0:0] tmp00_122_31;
	wire [WIDTH*2-1+0:0] tmp00_122_32;
	wire [WIDTH*2-1+0:0] tmp00_122_33;
	wire [WIDTH*2-1+0:0] tmp00_122_34;
	wire [WIDTH*2-1+0:0] tmp00_122_35;
	wire [WIDTH*2-1+0:0] tmp00_122_36;
	wire [WIDTH*2-1+0:0] tmp00_122_37;
	wire [WIDTH*2-1+0:0] tmp00_122_38;
	wire [WIDTH*2-1+0:0] tmp00_122_39;
	wire [WIDTH*2-1+0:0] tmp00_122_40;
	wire [WIDTH*2-1+0:0] tmp00_122_41;
	wire [WIDTH*2-1+0:0] tmp00_122_42;
	wire [WIDTH*2-1+0:0] tmp00_122_43;
	wire [WIDTH*2-1+0:0] tmp00_122_44;
	wire [WIDTH*2-1+0:0] tmp00_122_45;
	wire [WIDTH*2-1+0:0] tmp00_122_46;
	wire [WIDTH*2-1+0:0] tmp00_122_47;
	wire [WIDTH*2-1+0:0] tmp00_122_48;
	wire [WIDTH*2-1+0:0] tmp00_122_49;
	wire [WIDTH*2-1+0:0] tmp00_122_50;
	wire [WIDTH*2-1+0:0] tmp00_122_51;
	wire [WIDTH*2-1+0:0] tmp00_122_52;
	wire [WIDTH*2-1+0:0] tmp00_122_53;
	wire [WIDTH*2-1+0:0] tmp00_122_54;
	wire [WIDTH*2-1+0:0] tmp00_122_55;
	wire [WIDTH*2-1+0:0] tmp00_122_56;
	wire [WIDTH*2-1+0:0] tmp00_122_57;
	wire [WIDTH*2-1+0:0] tmp00_122_58;
	wire [WIDTH*2-1+0:0] tmp00_122_59;
	wire [WIDTH*2-1+0:0] tmp00_122_60;
	wire [WIDTH*2-1+0:0] tmp00_122_61;
	wire [WIDTH*2-1+0:0] tmp00_122_62;
	wire [WIDTH*2-1+0:0] tmp00_122_63;
	wire [WIDTH*2-1+0:0] tmp00_122_64;
	wire [WIDTH*2-1+0:0] tmp00_122_65;
	wire [WIDTH*2-1+0:0] tmp00_122_66;
	wire [WIDTH*2-1+0:0] tmp00_122_67;
	wire [WIDTH*2-1+0:0] tmp00_122_68;
	wire [WIDTH*2-1+0:0] tmp00_122_69;
	wire [WIDTH*2-1+0:0] tmp00_122_70;
	wire [WIDTH*2-1+0:0] tmp00_122_71;
	wire [WIDTH*2-1+0:0] tmp00_122_72;
	wire [WIDTH*2-1+0:0] tmp00_122_73;
	wire [WIDTH*2-1+0:0] tmp00_122_74;
	wire [WIDTH*2-1+0:0] tmp00_122_75;
	wire [WIDTH*2-1+0:0] tmp00_122_76;
	wire [WIDTH*2-1+0:0] tmp00_122_77;
	wire [WIDTH*2-1+0:0] tmp00_122_78;
	wire [WIDTH*2-1+0:0] tmp00_122_79;
	wire [WIDTH*2-1+0:0] tmp00_122_80;
	wire [WIDTH*2-1+0:0] tmp00_122_81;
	wire [WIDTH*2-1+0:0] tmp00_122_82;
	wire [WIDTH*2-1+0:0] tmp00_122_83;
	wire [WIDTH*2-1+0:0] tmp00_123_0;
	wire [WIDTH*2-1+0:0] tmp00_123_1;
	wire [WIDTH*2-1+0:0] tmp00_123_2;
	wire [WIDTH*2-1+0:0] tmp00_123_3;
	wire [WIDTH*2-1+0:0] tmp00_123_4;
	wire [WIDTH*2-1+0:0] tmp00_123_5;
	wire [WIDTH*2-1+0:0] tmp00_123_6;
	wire [WIDTH*2-1+0:0] tmp00_123_7;
	wire [WIDTH*2-1+0:0] tmp00_123_8;
	wire [WIDTH*2-1+0:0] tmp00_123_9;
	wire [WIDTH*2-1+0:0] tmp00_123_10;
	wire [WIDTH*2-1+0:0] tmp00_123_11;
	wire [WIDTH*2-1+0:0] tmp00_123_12;
	wire [WIDTH*2-1+0:0] tmp00_123_13;
	wire [WIDTH*2-1+0:0] tmp00_123_14;
	wire [WIDTH*2-1+0:0] tmp00_123_15;
	wire [WIDTH*2-1+0:0] tmp00_123_16;
	wire [WIDTH*2-1+0:0] tmp00_123_17;
	wire [WIDTH*2-1+0:0] tmp00_123_18;
	wire [WIDTH*2-1+0:0] tmp00_123_19;
	wire [WIDTH*2-1+0:0] tmp00_123_20;
	wire [WIDTH*2-1+0:0] tmp00_123_21;
	wire [WIDTH*2-1+0:0] tmp00_123_22;
	wire [WIDTH*2-1+0:0] tmp00_123_23;
	wire [WIDTH*2-1+0:0] tmp00_123_24;
	wire [WIDTH*2-1+0:0] tmp00_123_25;
	wire [WIDTH*2-1+0:0] tmp00_123_26;
	wire [WIDTH*2-1+0:0] tmp00_123_27;
	wire [WIDTH*2-1+0:0] tmp00_123_28;
	wire [WIDTH*2-1+0:0] tmp00_123_29;
	wire [WIDTH*2-1+0:0] tmp00_123_30;
	wire [WIDTH*2-1+0:0] tmp00_123_31;
	wire [WIDTH*2-1+0:0] tmp00_123_32;
	wire [WIDTH*2-1+0:0] tmp00_123_33;
	wire [WIDTH*2-1+0:0] tmp00_123_34;
	wire [WIDTH*2-1+0:0] tmp00_123_35;
	wire [WIDTH*2-1+0:0] tmp00_123_36;
	wire [WIDTH*2-1+0:0] tmp00_123_37;
	wire [WIDTH*2-1+0:0] tmp00_123_38;
	wire [WIDTH*2-1+0:0] tmp00_123_39;
	wire [WIDTH*2-1+0:0] tmp00_123_40;
	wire [WIDTH*2-1+0:0] tmp00_123_41;
	wire [WIDTH*2-1+0:0] tmp00_123_42;
	wire [WIDTH*2-1+0:0] tmp00_123_43;
	wire [WIDTH*2-1+0:0] tmp00_123_44;
	wire [WIDTH*2-1+0:0] tmp00_123_45;
	wire [WIDTH*2-1+0:0] tmp00_123_46;
	wire [WIDTH*2-1+0:0] tmp00_123_47;
	wire [WIDTH*2-1+0:0] tmp00_123_48;
	wire [WIDTH*2-1+0:0] tmp00_123_49;
	wire [WIDTH*2-1+0:0] tmp00_123_50;
	wire [WIDTH*2-1+0:0] tmp00_123_51;
	wire [WIDTH*2-1+0:0] tmp00_123_52;
	wire [WIDTH*2-1+0:0] tmp00_123_53;
	wire [WIDTH*2-1+0:0] tmp00_123_54;
	wire [WIDTH*2-1+0:0] tmp00_123_55;
	wire [WIDTH*2-1+0:0] tmp00_123_56;
	wire [WIDTH*2-1+0:0] tmp00_123_57;
	wire [WIDTH*2-1+0:0] tmp00_123_58;
	wire [WIDTH*2-1+0:0] tmp00_123_59;
	wire [WIDTH*2-1+0:0] tmp00_123_60;
	wire [WIDTH*2-1+0:0] tmp00_123_61;
	wire [WIDTH*2-1+0:0] tmp00_123_62;
	wire [WIDTH*2-1+0:0] tmp00_123_63;
	wire [WIDTH*2-1+0:0] tmp00_123_64;
	wire [WIDTH*2-1+0:0] tmp00_123_65;
	wire [WIDTH*2-1+0:0] tmp00_123_66;
	wire [WIDTH*2-1+0:0] tmp00_123_67;
	wire [WIDTH*2-1+0:0] tmp00_123_68;
	wire [WIDTH*2-1+0:0] tmp00_123_69;
	wire [WIDTH*2-1+0:0] tmp00_123_70;
	wire [WIDTH*2-1+0:0] tmp00_123_71;
	wire [WIDTH*2-1+0:0] tmp00_123_72;
	wire [WIDTH*2-1+0:0] tmp00_123_73;
	wire [WIDTH*2-1+0:0] tmp00_123_74;
	wire [WIDTH*2-1+0:0] tmp00_123_75;
	wire [WIDTH*2-1+0:0] tmp00_123_76;
	wire [WIDTH*2-1+0:0] tmp00_123_77;
	wire [WIDTH*2-1+0:0] tmp00_123_78;
	wire [WIDTH*2-1+0:0] tmp00_123_79;
	wire [WIDTH*2-1+0:0] tmp00_123_80;
	wire [WIDTH*2-1+0:0] tmp00_123_81;
	wire [WIDTH*2-1+0:0] tmp00_123_82;
	wire [WIDTH*2-1+0:0] tmp00_123_83;
	wire [WIDTH*2-1+0:0] tmp00_124_0;
	wire [WIDTH*2-1+0:0] tmp00_124_1;
	wire [WIDTH*2-1+0:0] tmp00_124_2;
	wire [WIDTH*2-1+0:0] tmp00_124_3;
	wire [WIDTH*2-1+0:0] tmp00_124_4;
	wire [WIDTH*2-1+0:0] tmp00_124_5;
	wire [WIDTH*2-1+0:0] tmp00_124_6;
	wire [WIDTH*2-1+0:0] tmp00_124_7;
	wire [WIDTH*2-1+0:0] tmp00_124_8;
	wire [WIDTH*2-1+0:0] tmp00_124_9;
	wire [WIDTH*2-1+0:0] tmp00_124_10;
	wire [WIDTH*2-1+0:0] tmp00_124_11;
	wire [WIDTH*2-1+0:0] tmp00_124_12;
	wire [WIDTH*2-1+0:0] tmp00_124_13;
	wire [WIDTH*2-1+0:0] tmp00_124_14;
	wire [WIDTH*2-1+0:0] tmp00_124_15;
	wire [WIDTH*2-1+0:0] tmp00_124_16;
	wire [WIDTH*2-1+0:0] tmp00_124_17;
	wire [WIDTH*2-1+0:0] tmp00_124_18;
	wire [WIDTH*2-1+0:0] tmp00_124_19;
	wire [WIDTH*2-1+0:0] tmp00_124_20;
	wire [WIDTH*2-1+0:0] tmp00_124_21;
	wire [WIDTH*2-1+0:0] tmp00_124_22;
	wire [WIDTH*2-1+0:0] tmp00_124_23;
	wire [WIDTH*2-1+0:0] tmp00_124_24;
	wire [WIDTH*2-1+0:0] tmp00_124_25;
	wire [WIDTH*2-1+0:0] tmp00_124_26;
	wire [WIDTH*2-1+0:0] tmp00_124_27;
	wire [WIDTH*2-1+0:0] tmp00_124_28;
	wire [WIDTH*2-1+0:0] tmp00_124_29;
	wire [WIDTH*2-1+0:0] tmp00_124_30;
	wire [WIDTH*2-1+0:0] tmp00_124_31;
	wire [WIDTH*2-1+0:0] tmp00_124_32;
	wire [WIDTH*2-1+0:0] tmp00_124_33;
	wire [WIDTH*2-1+0:0] tmp00_124_34;
	wire [WIDTH*2-1+0:0] tmp00_124_35;
	wire [WIDTH*2-1+0:0] tmp00_124_36;
	wire [WIDTH*2-1+0:0] tmp00_124_37;
	wire [WIDTH*2-1+0:0] tmp00_124_38;
	wire [WIDTH*2-1+0:0] tmp00_124_39;
	wire [WIDTH*2-1+0:0] tmp00_124_40;
	wire [WIDTH*2-1+0:0] tmp00_124_41;
	wire [WIDTH*2-1+0:0] tmp00_124_42;
	wire [WIDTH*2-1+0:0] tmp00_124_43;
	wire [WIDTH*2-1+0:0] tmp00_124_44;
	wire [WIDTH*2-1+0:0] tmp00_124_45;
	wire [WIDTH*2-1+0:0] tmp00_124_46;
	wire [WIDTH*2-1+0:0] tmp00_124_47;
	wire [WIDTH*2-1+0:0] tmp00_124_48;
	wire [WIDTH*2-1+0:0] tmp00_124_49;
	wire [WIDTH*2-1+0:0] tmp00_124_50;
	wire [WIDTH*2-1+0:0] tmp00_124_51;
	wire [WIDTH*2-1+0:0] tmp00_124_52;
	wire [WIDTH*2-1+0:0] tmp00_124_53;
	wire [WIDTH*2-1+0:0] tmp00_124_54;
	wire [WIDTH*2-1+0:0] tmp00_124_55;
	wire [WIDTH*2-1+0:0] tmp00_124_56;
	wire [WIDTH*2-1+0:0] tmp00_124_57;
	wire [WIDTH*2-1+0:0] tmp00_124_58;
	wire [WIDTH*2-1+0:0] tmp00_124_59;
	wire [WIDTH*2-1+0:0] tmp00_124_60;
	wire [WIDTH*2-1+0:0] tmp00_124_61;
	wire [WIDTH*2-1+0:0] tmp00_124_62;
	wire [WIDTH*2-1+0:0] tmp00_124_63;
	wire [WIDTH*2-1+0:0] tmp00_124_64;
	wire [WIDTH*2-1+0:0] tmp00_124_65;
	wire [WIDTH*2-1+0:0] tmp00_124_66;
	wire [WIDTH*2-1+0:0] tmp00_124_67;
	wire [WIDTH*2-1+0:0] tmp00_124_68;
	wire [WIDTH*2-1+0:0] tmp00_124_69;
	wire [WIDTH*2-1+0:0] tmp00_124_70;
	wire [WIDTH*2-1+0:0] tmp00_124_71;
	wire [WIDTH*2-1+0:0] tmp00_124_72;
	wire [WIDTH*2-1+0:0] tmp00_124_73;
	wire [WIDTH*2-1+0:0] tmp00_124_74;
	wire [WIDTH*2-1+0:0] tmp00_124_75;
	wire [WIDTH*2-1+0:0] tmp00_124_76;
	wire [WIDTH*2-1+0:0] tmp00_124_77;
	wire [WIDTH*2-1+0:0] tmp00_124_78;
	wire [WIDTH*2-1+0:0] tmp00_124_79;
	wire [WIDTH*2-1+0:0] tmp00_124_80;
	wire [WIDTH*2-1+0:0] tmp00_124_81;
	wire [WIDTH*2-1+0:0] tmp00_124_82;
	wire [WIDTH*2-1+0:0] tmp00_124_83;
	wire [WIDTH*2-1+0:0] tmp00_125_0;
	wire [WIDTH*2-1+0:0] tmp00_125_1;
	wire [WIDTH*2-1+0:0] tmp00_125_2;
	wire [WIDTH*2-1+0:0] tmp00_125_3;
	wire [WIDTH*2-1+0:0] tmp00_125_4;
	wire [WIDTH*2-1+0:0] tmp00_125_5;
	wire [WIDTH*2-1+0:0] tmp00_125_6;
	wire [WIDTH*2-1+0:0] tmp00_125_7;
	wire [WIDTH*2-1+0:0] tmp00_125_8;
	wire [WIDTH*2-1+0:0] tmp00_125_9;
	wire [WIDTH*2-1+0:0] tmp00_125_10;
	wire [WIDTH*2-1+0:0] tmp00_125_11;
	wire [WIDTH*2-1+0:0] tmp00_125_12;
	wire [WIDTH*2-1+0:0] tmp00_125_13;
	wire [WIDTH*2-1+0:0] tmp00_125_14;
	wire [WIDTH*2-1+0:0] tmp00_125_15;
	wire [WIDTH*2-1+0:0] tmp00_125_16;
	wire [WIDTH*2-1+0:0] tmp00_125_17;
	wire [WIDTH*2-1+0:0] tmp00_125_18;
	wire [WIDTH*2-1+0:0] tmp00_125_19;
	wire [WIDTH*2-1+0:0] tmp00_125_20;
	wire [WIDTH*2-1+0:0] tmp00_125_21;
	wire [WIDTH*2-1+0:0] tmp00_125_22;
	wire [WIDTH*2-1+0:0] tmp00_125_23;
	wire [WIDTH*2-1+0:0] tmp00_125_24;
	wire [WIDTH*2-1+0:0] tmp00_125_25;
	wire [WIDTH*2-1+0:0] tmp00_125_26;
	wire [WIDTH*2-1+0:0] tmp00_125_27;
	wire [WIDTH*2-1+0:0] tmp00_125_28;
	wire [WIDTH*2-1+0:0] tmp00_125_29;
	wire [WIDTH*2-1+0:0] tmp00_125_30;
	wire [WIDTH*2-1+0:0] tmp00_125_31;
	wire [WIDTH*2-1+0:0] tmp00_125_32;
	wire [WIDTH*2-1+0:0] tmp00_125_33;
	wire [WIDTH*2-1+0:0] tmp00_125_34;
	wire [WIDTH*2-1+0:0] tmp00_125_35;
	wire [WIDTH*2-1+0:0] tmp00_125_36;
	wire [WIDTH*2-1+0:0] tmp00_125_37;
	wire [WIDTH*2-1+0:0] tmp00_125_38;
	wire [WIDTH*2-1+0:0] tmp00_125_39;
	wire [WIDTH*2-1+0:0] tmp00_125_40;
	wire [WIDTH*2-1+0:0] tmp00_125_41;
	wire [WIDTH*2-1+0:0] tmp00_125_42;
	wire [WIDTH*2-1+0:0] tmp00_125_43;
	wire [WIDTH*2-1+0:0] tmp00_125_44;
	wire [WIDTH*2-1+0:0] tmp00_125_45;
	wire [WIDTH*2-1+0:0] tmp00_125_46;
	wire [WIDTH*2-1+0:0] tmp00_125_47;
	wire [WIDTH*2-1+0:0] tmp00_125_48;
	wire [WIDTH*2-1+0:0] tmp00_125_49;
	wire [WIDTH*2-1+0:0] tmp00_125_50;
	wire [WIDTH*2-1+0:0] tmp00_125_51;
	wire [WIDTH*2-1+0:0] tmp00_125_52;
	wire [WIDTH*2-1+0:0] tmp00_125_53;
	wire [WIDTH*2-1+0:0] tmp00_125_54;
	wire [WIDTH*2-1+0:0] tmp00_125_55;
	wire [WIDTH*2-1+0:0] tmp00_125_56;
	wire [WIDTH*2-1+0:0] tmp00_125_57;
	wire [WIDTH*2-1+0:0] tmp00_125_58;
	wire [WIDTH*2-1+0:0] tmp00_125_59;
	wire [WIDTH*2-1+0:0] tmp00_125_60;
	wire [WIDTH*2-1+0:0] tmp00_125_61;
	wire [WIDTH*2-1+0:0] tmp00_125_62;
	wire [WIDTH*2-1+0:0] tmp00_125_63;
	wire [WIDTH*2-1+0:0] tmp00_125_64;
	wire [WIDTH*2-1+0:0] tmp00_125_65;
	wire [WIDTH*2-1+0:0] tmp00_125_66;
	wire [WIDTH*2-1+0:0] tmp00_125_67;
	wire [WIDTH*2-1+0:0] tmp00_125_68;
	wire [WIDTH*2-1+0:0] tmp00_125_69;
	wire [WIDTH*2-1+0:0] tmp00_125_70;
	wire [WIDTH*2-1+0:0] tmp00_125_71;
	wire [WIDTH*2-1+0:0] tmp00_125_72;
	wire [WIDTH*2-1+0:0] tmp00_125_73;
	wire [WIDTH*2-1+0:0] tmp00_125_74;
	wire [WIDTH*2-1+0:0] tmp00_125_75;
	wire [WIDTH*2-1+0:0] tmp00_125_76;
	wire [WIDTH*2-1+0:0] tmp00_125_77;
	wire [WIDTH*2-1+0:0] tmp00_125_78;
	wire [WIDTH*2-1+0:0] tmp00_125_79;
	wire [WIDTH*2-1+0:0] tmp00_125_80;
	wire [WIDTH*2-1+0:0] tmp00_125_81;
	wire [WIDTH*2-1+0:0] tmp00_125_82;
	wire [WIDTH*2-1+0:0] tmp00_125_83;
	wire [WIDTH*2-1+0:0] tmp00_126_0;
	wire [WIDTH*2-1+0:0] tmp00_126_1;
	wire [WIDTH*2-1+0:0] tmp00_126_2;
	wire [WIDTH*2-1+0:0] tmp00_126_3;
	wire [WIDTH*2-1+0:0] tmp00_126_4;
	wire [WIDTH*2-1+0:0] tmp00_126_5;
	wire [WIDTH*2-1+0:0] tmp00_126_6;
	wire [WIDTH*2-1+0:0] tmp00_126_7;
	wire [WIDTH*2-1+0:0] tmp00_126_8;
	wire [WIDTH*2-1+0:0] tmp00_126_9;
	wire [WIDTH*2-1+0:0] tmp00_126_10;
	wire [WIDTH*2-1+0:0] tmp00_126_11;
	wire [WIDTH*2-1+0:0] tmp00_126_12;
	wire [WIDTH*2-1+0:0] tmp00_126_13;
	wire [WIDTH*2-1+0:0] tmp00_126_14;
	wire [WIDTH*2-1+0:0] tmp00_126_15;
	wire [WIDTH*2-1+0:0] tmp00_126_16;
	wire [WIDTH*2-1+0:0] tmp00_126_17;
	wire [WIDTH*2-1+0:0] tmp00_126_18;
	wire [WIDTH*2-1+0:0] tmp00_126_19;
	wire [WIDTH*2-1+0:0] tmp00_126_20;
	wire [WIDTH*2-1+0:0] tmp00_126_21;
	wire [WIDTH*2-1+0:0] tmp00_126_22;
	wire [WIDTH*2-1+0:0] tmp00_126_23;
	wire [WIDTH*2-1+0:0] tmp00_126_24;
	wire [WIDTH*2-1+0:0] tmp00_126_25;
	wire [WIDTH*2-1+0:0] tmp00_126_26;
	wire [WIDTH*2-1+0:0] tmp00_126_27;
	wire [WIDTH*2-1+0:0] tmp00_126_28;
	wire [WIDTH*2-1+0:0] tmp00_126_29;
	wire [WIDTH*2-1+0:0] tmp00_126_30;
	wire [WIDTH*2-1+0:0] tmp00_126_31;
	wire [WIDTH*2-1+0:0] tmp00_126_32;
	wire [WIDTH*2-1+0:0] tmp00_126_33;
	wire [WIDTH*2-1+0:0] tmp00_126_34;
	wire [WIDTH*2-1+0:0] tmp00_126_35;
	wire [WIDTH*2-1+0:0] tmp00_126_36;
	wire [WIDTH*2-1+0:0] tmp00_126_37;
	wire [WIDTH*2-1+0:0] tmp00_126_38;
	wire [WIDTH*2-1+0:0] tmp00_126_39;
	wire [WIDTH*2-1+0:0] tmp00_126_40;
	wire [WIDTH*2-1+0:0] tmp00_126_41;
	wire [WIDTH*2-1+0:0] tmp00_126_42;
	wire [WIDTH*2-1+0:0] tmp00_126_43;
	wire [WIDTH*2-1+0:0] tmp00_126_44;
	wire [WIDTH*2-1+0:0] tmp00_126_45;
	wire [WIDTH*2-1+0:0] tmp00_126_46;
	wire [WIDTH*2-1+0:0] tmp00_126_47;
	wire [WIDTH*2-1+0:0] tmp00_126_48;
	wire [WIDTH*2-1+0:0] tmp00_126_49;
	wire [WIDTH*2-1+0:0] tmp00_126_50;
	wire [WIDTH*2-1+0:0] tmp00_126_51;
	wire [WIDTH*2-1+0:0] tmp00_126_52;
	wire [WIDTH*2-1+0:0] tmp00_126_53;
	wire [WIDTH*2-1+0:0] tmp00_126_54;
	wire [WIDTH*2-1+0:0] tmp00_126_55;
	wire [WIDTH*2-1+0:0] tmp00_126_56;
	wire [WIDTH*2-1+0:0] tmp00_126_57;
	wire [WIDTH*2-1+0:0] tmp00_126_58;
	wire [WIDTH*2-1+0:0] tmp00_126_59;
	wire [WIDTH*2-1+0:0] tmp00_126_60;
	wire [WIDTH*2-1+0:0] tmp00_126_61;
	wire [WIDTH*2-1+0:0] tmp00_126_62;
	wire [WIDTH*2-1+0:0] tmp00_126_63;
	wire [WIDTH*2-1+0:0] tmp00_126_64;
	wire [WIDTH*2-1+0:0] tmp00_126_65;
	wire [WIDTH*2-1+0:0] tmp00_126_66;
	wire [WIDTH*2-1+0:0] tmp00_126_67;
	wire [WIDTH*2-1+0:0] tmp00_126_68;
	wire [WIDTH*2-1+0:0] tmp00_126_69;
	wire [WIDTH*2-1+0:0] tmp00_126_70;
	wire [WIDTH*2-1+0:0] tmp00_126_71;
	wire [WIDTH*2-1+0:0] tmp00_126_72;
	wire [WIDTH*2-1+0:0] tmp00_126_73;
	wire [WIDTH*2-1+0:0] tmp00_126_74;
	wire [WIDTH*2-1+0:0] tmp00_126_75;
	wire [WIDTH*2-1+0:0] tmp00_126_76;
	wire [WIDTH*2-1+0:0] tmp00_126_77;
	wire [WIDTH*2-1+0:0] tmp00_126_78;
	wire [WIDTH*2-1+0:0] tmp00_126_79;
	wire [WIDTH*2-1+0:0] tmp00_126_80;
	wire [WIDTH*2-1+0:0] tmp00_126_81;
	wire [WIDTH*2-1+0:0] tmp00_126_82;
	wire [WIDTH*2-1+0:0] tmp00_126_83;
	wire [WIDTH*2-1+0:0] tmp00_127_0;
	wire [WIDTH*2-1+0:0] tmp00_127_1;
	wire [WIDTH*2-1+0:0] tmp00_127_2;
	wire [WIDTH*2-1+0:0] tmp00_127_3;
	wire [WIDTH*2-1+0:0] tmp00_127_4;
	wire [WIDTH*2-1+0:0] tmp00_127_5;
	wire [WIDTH*2-1+0:0] tmp00_127_6;
	wire [WIDTH*2-1+0:0] tmp00_127_7;
	wire [WIDTH*2-1+0:0] tmp00_127_8;
	wire [WIDTH*2-1+0:0] tmp00_127_9;
	wire [WIDTH*2-1+0:0] tmp00_127_10;
	wire [WIDTH*2-1+0:0] tmp00_127_11;
	wire [WIDTH*2-1+0:0] tmp00_127_12;
	wire [WIDTH*2-1+0:0] tmp00_127_13;
	wire [WIDTH*2-1+0:0] tmp00_127_14;
	wire [WIDTH*2-1+0:0] tmp00_127_15;
	wire [WIDTH*2-1+0:0] tmp00_127_16;
	wire [WIDTH*2-1+0:0] tmp00_127_17;
	wire [WIDTH*2-1+0:0] tmp00_127_18;
	wire [WIDTH*2-1+0:0] tmp00_127_19;
	wire [WIDTH*2-1+0:0] tmp00_127_20;
	wire [WIDTH*2-1+0:0] tmp00_127_21;
	wire [WIDTH*2-1+0:0] tmp00_127_22;
	wire [WIDTH*2-1+0:0] tmp00_127_23;
	wire [WIDTH*2-1+0:0] tmp00_127_24;
	wire [WIDTH*2-1+0:0] tmp00_127_25;
	wire [WIDTH*2-1+0:0] tmp00_127_26;
	wire [WIDTH*2-1+0:0] tmp00_127_27;
	wire [WIDTH*2-1+0:0] tmp00_127_28;
	wire [WIDTH*2-1+0:0] tmp00_127_29;
	wire [WIDTH*2-1+0:0] tmp00_127_30;
	wire [WIDTH*2-1+0:0] tmp00_127_31;
	wire [WIDTH*2-1+0:0] tmp00_127_32;
	wire [WIDTH*2-1+0:0] tmp00_127_33;
	wire [WIDTH*2-1+0:0] tmp00_127_34;
	wire [WIDTH*2-1+0:0] tmp00_127_35;
	wire [WIDTH*2-1+0:0] tmp00_127_36;
	wire [WIDTH*2-1+0:0] tmp00_127_37;
	wire [WIDTH*2-1+0:0] tmp00_127_38;
	wire [WIDTH*2-1+0:0] tmp00_127_39;
	wire [WIDTH*2-1+0:0] tmp00_127_40;
	wire [WIDTH*2-1+0:0] tmp00_127_41;
	wire [WIDTH*2-1+0:0] tmp00_127_42;
	wire [WIDTH*2-1+0:0] tmp00_127_43;
	wire [WIDTH*2-1+0:0] tmp00_127_44;
	wire [WIDTH*2-1+0:0] tmp00_127_45;
	wire [WIDTH*2-1+0:0] tmp00_127_46;
	wire [WIDTH*2-1+0:0] tmp00_127_47;
	wire [WIDTH*2-1+0:0] tmp00_127_48;
	wire [WIDTH*2-1+0:0] tmp00_127_49;
	wire [WIDTH*2-1+0:0] tmp00_127_50;
	wire [WIDTH*2-1+0:0] tmp00_127_51;
	wire [WIDTH*2-1+0:0] tmp00_127_52;
	wire [WIDTH*2-1+0:0] tmp00_127_53;
	wire [WIDTH*2-1+0:0] tmp00_127_54;
	wire [WIDTH*2-1+0:0] tmp00_127_55;
	wire [WIDTH*2-1+0:0] tmp00_127_56;
	wire [WIDTH*2-1+0:0] tmp00_127_57;
	wire [WIDTH*2-1+0:0] tmp00_127_58;
	wire [WIDTH*2-1+0:0] tmp00_127_59;
	wire [WIDTH*2-1+0:0] tmp00_127_60;
	wire [WIDTH*2-1+0:0] tmp00_127_61;
	wire [WIDTH*2-1+0:0] tmp00_127_62;
	wire [WIDTH*2-1+0:0] tmp00_127_63;
	wire [WIDTH*2-1+0:0] tmp00_127_64;
	wire [WIDTH*2-1+0:0] tmp00_127_65;
	wire [WIDTH*2-1+0:0] tmp00_127_66;
	wire [WIDTH*2-1+0:0] tmp00_127_67;
	wire [WIDTH*2-1+0:0] tmp00_127_68;
	wire [WIDTH*2-1+0:0] tmp00_127_69;
	wire [WIDTH*2-1+0:0] tmp00_127_70;
	wire [WIDTH*2-1+0:0] tmp00_127_71;
	wire [WIDTH*2-1+0:0] tmp00_127_72;
	wire [WIDTH*2-1+0:0] tmp00_127_73;
	wire [WIDTH*2-1+0:0] tmp00_127_74;
	wire [WIDTH*2-1+0:0] tmp00_127_75;
	wire [WIDTH*2-1+0:0] tmp00_127_76;
	wire [WIDTH*2-1+0:0] tmp00_127_77;
	wire [WIDTH*2-1+0:0] tmp00_127_78;
	wire [WIDTH*2-1+0:0] tmp00_127_79;
	wire [WIDTH*2-1+0:0] tmp00_127_80;
	wire [WIDTH*2-1+0:0] tmp00_127_81;
	wire [WIDTH*2-1+0:0] tmp00_127_82;
	wire [WIDTH*2-1+0:0] tmp00_127_83;
	wire [WIDTH*2-1+1:0] tmp01_0_0;
	wire [WIDTH*2-1+1:0] tmp01_0_1;
	wire [WIDTH*2-1+1:0] tmp01_0_2;
	wire [WIDTH*2-1+1:0] tmp01_0_3;
	wire [WIDTH*2-1+1:0] tmp01_0_4;
	wire [WIDTH*2-1+1:0] tmp01_0_5;
	wire [WIDTH*2-1+1:0] tmp01_0_6;
	wire [WIDTH*2-1+1:0] tmp01_0_7;
	wire [WIDTH*2-1+1:0] tmp01_0_8;
	wire [WIDTH*2-1+1:0] tmp01_0_9;
	wire [WIDTH*2-1+1:0] tmp01_0_10;
	wire [WIDTH*2-1+1:0] tmp01_0_11;
	wire [WIDTH*2-1+1:0] tmp01_0_12;
	wire [WIDTH*2-1+1:0] tmp01_0_13;
	wire [WIDTH*2-1+1:0] tmp01_0_14;
	wire [WIDTH*2-1+1:0] tmp01_0_15;
	wire [WIDTH*2-1+1:0] tmp01_0_16;
	wire [WIDTH*2-1+1:0] tmp01_0_17;
	wire [WIDTH*2-1+1:0] tmp01_0_18;
	wire [WIDTH*2-1+1:0] tmp01_0_19;
	wire [WIDTH*2-1+1:0] tmp01_0_20;
	wire [WIDTH*2-1+1:0] tmp01_0_21;
	wire [WIDTH*2-1+1:0] tmp01_0_22;
	wire [WIDTH*2-1+1:0] tmp01_0_23;
	wire [WIDTH*2-1+1:0] tmp01_0_24;
	wire [WIDTH*2-1+1:0] tmp01_0_25;
	wire [WIDTH*2-1+1:0] tmp01_0_26;
	wire [WIDTH*2-1+1:0] tmp01_0_27;
	wire [WIDTH*2-1+1:0] tmp01_0_28;
	wire [WIDTH*2-1+1:0] tmp01_0_29;
	wire [WIDTH*2-1+1:0] tmp01_0_30;
	wire [WIDTH*2-1+1:0] tmp01_0_31;
	wire [WIDTH*2-1+1:0] tmp01_0_32;
	wire [WIDTH*2-1+1:0] tmp01_0_33;
	wire [WIDTH*2-1+1:0] tmp01_0_34;
	wire [WIDTH*2-1+1:0] tmp01_0_35;
	wire [WIDTH*2-1+1:0] tmp01_0_36;
	wire [WIDTH*2-1+1:0] tmp01_0_37;
	wire [WIDTH*2-1+1:0] tmp01_0_38;
	wire [WIDTH*2-1+1:0] tmp01_0_39;
	wire [WIDTH*2-1+1:0] tmp01_0_40;
	wire [WIDTH*2-1+1:0] tmp01_0_41;
	wire [WIDTH*2-1+1:0] tmp01_0_42;
	wire [WIDTH*2-1+1:0] tmp01_0_43;
	wire [WIDTH*2-1+1:0] tmp01_0_44;
	wire [WIDTH*2-1+1:0] tmp01_0_45;
	wire [WIDTH*2-1+1:0] tmp01_0_46;
	wire [WIDTH*2-1+1:0] tmp01_0_47;
	wire [WIDTH*2-1+1:0] tmp01_0_48;
	wire [WIDTH*2-1+1:0] tmp01_0_49;
	wire [WIDTH*2-1+1:0] tmp01_0_50;
	wire [WIDTH*2-1+1:0] tmp01_0_51;
	wire [WIDTH*2-1+1:0] tmp01_0_52;
	wire [WIDTH*2-1+1:0] tmp01_0_53;
	wire [WIDTH*2-1+1:0] tmp01_0_54;
	wire [WIDTH*2-1+1:0] tmp01_0_55;
	wire [WIDTH*2-1+1:0] tmp01_0_56;
	wire [WIDTH*2-1+1:0] tmp01_0_57;
	wire [WIDTH*2-1+1:0] tmp01_0_58;
	wire [WIDTH*2-1+1:0] tmp01_0_59;
	wire [WIDTH*2-1+1:0] tmp01_0_60;
	wire [WIDTH*2-1+1:0] tmp01_0_61;
	wire [WIDTH*2-1+1:0] tmp01_0_62;
	wire [WIDTH*2-1+1:0] tmp01_0_63;
	wire [WIDTH*2-1+1:0] tmp01_0_64;
	wire [WIDTH*2-1+1:0] tmp01_0_65;
	wire [WIDTH*2-1+1:0] tmp01_0_66;
	wire [WIDTH*2-1+1:0] tmp01_0_67;
	wire [WIDTH*2-1+1:0] tmp01_0_68;
	wire [WIDTH*2-1+1:0] tmp01_0_69;
	wire [WIDTH*2-1+1:0] tmp01_0_70;
	wire [WIDTH*2-1+1:0] tmp01_0_71;
	wire [WIDTH*2-1+1:0] tmp01_0_72;
	wire [WIDTH*2-1+1:0] tmp01_0_73;
	wire [WIDTH*2-1+1:0] tmp01_0_74;
	wire [WIDTH*2-1+1:0] tmp01_0_75;
	wire [WIDTH*2-1+1:0] tmp01_0_76;
	wire [WIDTH*2-1+1:0] tmp01_0_77;
	wire [WIDTH*2-1+1:0] tmp01_0_78;
	wire [WIDTH*2-1+1:0] tmp01_0_79;
	wire [WIDTH*2-1+1:0] tmp01_0_80;
	wire [WIDTH*2-1+1:0] tmp01_0_81;
	wire [WIDTH*2-1+1:0] tmp01_0_82;
	wire [WIDTH*2-1+1:0] tmp01_0_83;
	wire [WIDTH*2-1+1:0] tmp01_1_0;
	wire [WIDTH*2-1+1:0] tmp01_1_1;
	wire [WIDTH*2-1+1:0] tmp01_1_2;
	wire [WIDTH*2-1+1:0] tmp01_1_3;
	wire [WIDTH*2-1+1:0] tmp01_1_4;
	wire [WIDTH*2-1+1:0] tmp01_1_5;
	wire [WIDTH*2-1+1:0] tmp01_1_6;
	wire [WIDTH*2-1+1:0] tmp01_1_7;
	wire [WIDTH*2-1+1:0] tmp01_1_8;
	wire [WIDTH*2-1+1:0] tmp01_1_9;
	wire [WIDTH*2-1+1:0] tmp01_1_10;
	wire [WIDTH*2-1+1:0] tmp01_1_11;
	wire [WIDTH*2-1+1:0] tmp01_1_12;
	wire [WIDTH*2-1+1:0] tmp01_1_13;
	wire [WIDTH*2-1+1:0] tmp01_1_14;
	wire [WIDTH*2-1+1:0] tmp01_1_15;
	wire [WIDTH*2-1+1:0] tmp01_1_16;
	wire [WIDTH*2-1+1:0] tmp01_1_17;
	wire [WIDTH*2-1+1:0] tmp01_1_18;
	wire [WIDTH*2-1+1:0] tmp01_1_19;
	wire [WIDTH*2-1+1:0] tmp01_1_20;
	wire [WIDTH*2-1+1:0] tmp01_1_21;
	wire [WIDTH*2-1+1:0] tmp01_1_22;
	wire [WIDTH*2-1+1:0] tmp01_1_23;
	wire [WIDTH*2-1+1:0] tmp01_1_24;
	wire [WIDTH*2-1+1:0] tmp01_1_25;
	wire [WIDTH*2-1+1:0] tmp01_1_26;
	wire [WIDTH*2-1+1:0] tmp01_1_27;
	wire [WIDTH*2-1+1:0] tmp01_1_28;
	wire [WIDTH*2-1+1:0] tmp01_1_29;
	wire [WIDTH*2-1+1:0] tmp01_1_30;
	wire [WIDTH*2-1+1:0] tmp01_1_31;
	wire [WIDTH*2-1+1:0] tmp01_1_32;
	wire [WIDTH*2-1+1:0] tmp01_1_33;
	wire [WIDTH*2-1+1:0] tmp01_1_34;
	wire [WIDTH*2-1+1:0] tmp01_1_35;
	wire [WIDTH*2-1+1:0] tmp01_1_36;
	wire [WIDTH*2-1+1:0] tmp01_1_37;
	wire [WIDTH*2-1+1:0] tmp01_1_38;
	wire [WIDTH*2-1+1:0] tmp01_1_39;
	wire [WIDTH*2-1+1:0] tmp01_1_40;
	wire [WIDTH*2-1+1:0] tmp01_1_41;
	wire [WIDTH*2-1+1:0] tmp01_1_42;
	wire [WIDTH*2-1+1:0] tmp01_1_43;
	wire [WIDTH*2-1+1:0] tmp01_1_44;
	wire [WIDTH*2-1+1:0] tmp01_1_45;
	wire [WIDTH*2-1+1:0] tmp01_1_46;
	wire [WIDTH*2-1+1:0] tmp01_1_47;
	wire [WIDTH*2-1+1:0] tmp01_1_48;
	wire [WIDTH*2-1+1:0] tmp01_1_49;
	wire [WIDTH*2-1+1:0] tmp01_1_50;
	wire [WIDTH*2-1+1:0] tmp01_1_51;
	wire [WIDTH*2-1+1:0] tmp01_1_52;
	wire [WIDTH*2-1+1:0] tmp01_1_53;
	wire [WIDTH*2-1+1:0] tmp01_1_54;
	wire [WIDTH*2-1+1:0] tmp01_1_55;
	wire [WIDTH*2-1+1:0] tmp01_1_56;
	wire [WIDTH*2-1+1:0] tmp01_1_57;
	wire [WIDTH*2-1+1:0] tmp01_1_58;
	wire [WIDTH*2-1+1:0] tmp01_1_59;
	wire [WIDTH*2-1+1:0] tmp01_1_60;
	wire [WIDTH*2-1+1:0] tmp01_1_61;
	wire [WIDTH*2-1+1:0] tmp01_1_62;
	wire [WIDTH*2-1+1:0] tmp01_1_63;
	wire [WIDTH*2-1+1:0] tmp01_1_64;
	wire [WIDTH*2-1+1:0] tmp01_1_65;
	wire [WIDTH*2-1+1:0] tmp01_1_66;
	wire [WIDTH*2-1+1:0] tmp01_1_67;
	wire [WIDTH*2-1+1:0] tmp01_1_68;
	wire [WIDTH*2-1+1:0] tmp01_1_69;
	wire [WIDTH*2-1+1:0] tmp01_1_70;
	wire [WIDTH*2-1+1:0] tmp01_1_71;
	wire [WIDTH*2-1+1:0] tmp01_1_72;
	wire [WIDTH*2-1+1:0] tmp01_1_73;
	wire [WIDTH*2-1+1:0] tmp01_1_74;
	wire [WIDTH*2-1+1:0] tmp01_1_75;
	wire [WIDTH*2-1+1:0] tmp01_1_76;
	wire [WIDTH*2-1+1:0] tmp01_1_77;
	wire [WIDTH*2-1+1:0] tmp01_1_78;
	wire [WIDTH*2-1+1:0] tmp01_1_79;
	wire [WIDTH*2-1+1:0] tmp01_1_80;
	wire [WIDTH*2-1+1:0] tmp01_1_81;
	wire [WIDTH*2-1+1:0] tmp01_1_82;
	wire [WIDTH*2-1+1:0] tmp01_1_83;
	wire [WIDTH*2-1+1:0] tmp01_2_0;
	wire [WIDTH*2-1+1:0] tmp01_2_1;
	wire [WIDTH*2-1+1:0] tmp01_2_2;
	wire [WIDTH*2-1+1:0] tmp01_2_3;
	wire [WIDTH*2-1+1:0] tmp01_2_4;
	wire [WIDTH*2-1+1:0] tmp01_2_5;
	wire [WIDTH*2-1+1:0] tmp01_2_6;
	wire [WIDTH*2-1+1:0] tmp01_2_7;
	wire [WIDTH*2-1+1:0] tmp01_2_8;
	wire [WIDTH*2-1+1:0] tmp01_2_9;
	wire [WIDTH*2-1+1:0] tmp01_2_10;
	wire [WIDTH*2-1+1:0] tmp01_2_11;
	wire [WIDTH*2-1+1:0] tmp01_2_12;
	wire [WIDTH*2-1+1:0] tmp01_2_13;
	wire [WIDTH*2-1+1:0] tmp01_2_14;
	wire [WIDTH*2-1+1:0] tmp01_2_15;
	wire [WIDTH*2-1+1:0] tmp01_2_16;
	wire [WIDTH*2-1+1:0] tmp01_2_17;
	wire [WIDTH*2-1+1:0] tmp01_2_18;
	wire [WIDTH*2-1+1:0] tmp01_2_19;
	wire [WIDTH*2-1+1:0] tmp01_2_20;
	wire [WIDTH*2-1+1:0] tmp01_2_21;
	wire [WIDTH*2-1+1:0] tmp01_2_22;
	wire [WIDTH*2-1+1:0] tmp01_2_23;
	wire [WIDTH*2-1+1:0] tmp01_2_24;
	wire [WIDTH*2-1+1:0] tmp01_2_25;
	wire [WIDTH*2-1+1:0] tmp01_2_26;
	wire [WIDTH*2-1+1:0] tmp01_2_27;
	wire [WIDTH*2-1+1:0] tmp01_2_28;
	wire [WIDTH*2-1+1:0] tmp01_2_29;
	wire [WIDTH*2-1+1:0] tmp01_2_30;
	wire [WIDTH*2-1+1:0] tmp01_2_31;
	wire [WIDTH*2-1+1:0] tmp01_2_32;
	wire [WIDTH*2-1+1:0] tmp01_2_33;
	wire [WIDTH*2-1+1:0] tmp01_2_34;
	wire [WIDTH*2-1+1:0] tmp01_2_35;
	wire [WIDTH*2-1+1:0] tmp01_2_36;
	wire [WIDTH*2-1+1:0] tmp01_2_37;
	wire [WIDTH*2-1+1:0] tmp01_2_38;
	wire [WIDTH*2-1+1:0] tmp01_2_39;
	wire [WIDTH*2-1+1:0] tmp01_2_40;
	wire [WIDTH*2-1+1:0] tmp01_2_41;
	wire [WIDTH*2-1+1:0] tmp01_2_42;
	wire [WIDTH*2-1+1:0] tmp01_2_43;
	wire [WIDTH*2-1+1:0] tmp01_2_44;
	wire [WIDTH*2-1+1:0] tmp01_2_45;
	wire [WIDTH*2-1+1:0] tmp01_2_46;
	wire [WIDTH*2-1+1:0] tmp01_2_47;
	wire [WIDTH*2-1+1:0] tmp01_2_48;
	wire [WIDTH*2-1+1:0] tmp01_2_49;
	wire [WIDTH*2-1+1:0] tmp01_2_50;
	wire [WIDTH*2-1+1:0] tmp01_2_51;
	wire [WIDTH*2-1+1:0] tmp01_2_52;
	wire [WIDTH*2-1+1:0] tmp01_2_53;
	wire [WIDTH*2-1+1:0] tmp01_2_54;
	wire [WIDTH*2-1+1:0] tmp01_2_55;
	wire [WIDTH*2-1+1:0] tmp01_2_56;
	wire [WIDTH*2-1+1:0] tmp01_2_57;
	wire [WIDTH*2-1+1:0] tmp01_2_58;
	wire [WIDTH*2-1+1:0] tmp01_2_59;
	wire [WIDTH*2-1+1:0] tmp01_2_60;
	wire [WIDTH*2-1+1:0] tmp01_2_61;
	wire [WIDTH*2-1+1:0] tmp01_2_62;
	wire [WIDTH*2-1+1:0] tmp01_2_63;
	wire [WIDTH*2-1+1:0] tmp01_2_64;
	wire [WIDTH*2-1+1:0] tmp01_2_65;
	wire [WIDTH*2-1+1:0] tmp01_2_66;
	wire [WIDTH*2-1+1:0] tmp01_2_67;
	wire [WIDTH*2-1+1:0] tmp01_2_68;
	wire [WIDTH*2-1+1:0] tmp01_2_69;
	wire [WIDTH*2-1+1:0] tmp01_2_70;
	wire [WIDTH*2-1+1:0] tmp01_2_71;
	wire [WIDTH*2-1+1:0] tmp01_2_72;
	wire [WIDTH*2-1+1:0] tmp01_2_73;
	wire [WIDTH*2-1+1:0] tmp01_2_74;
	wire [WIDTH*2-1+1:0] tmp01_2_75;
	wire [WIDTH*2-1+1:0] tmp01_2_76;
	wire [WIDTH*2-1+1:0] tmp01_2_77;
	wire [WIDTH*2-1+1:0] tmp01_2_78;
	wire [WIDTH*2-1+1:0] tmp01_2_79;
	wire [WIDTH*2-1+1:0] tmp01_2_80;
	wire [WIDTH*2-1+1:0] tmp01_2_81;
	wire [WIDTH*2-1+1:0] tmp01_2_82;
	wire [WIDTH*2-1+1:0] tmp01_2_83;
	wire [WIDTH*2-1+1:0] tmp01_3_0;
	wire [WIDTH*2-1+1:0] tmp01_3_1;
	wire [WIDTH*2-1+1:0] tmp01_3_2;
	wire [WIDTH*2-1+1:0] tmp01_3_3;
	wire [WIDTH*2-1+1:0] tmp01_3_4;
	wire [WIDTH*2-1+1:0] tmp01_3_5;
	wire [WIDTH*2-1+1:0] tmp01_3_6;
	wire [WIDTH*2-1+1:0] tmp01_3_7;
	wire [WIDTH*2-1+1:0] tmp01_3_8;
	wire [WIDTH*2-1+1:0] tmp01_3_9;
	wire [WIDTH*2-1+1:0] tmp01_3_10;
	wire [WIDTH*2-1+1:0] tmp01_3_11;
	wire [WIDTH*2-1+1:0] tmp01_3_12;
	wire [WIDTH*2-1+1:0] tmp01_3_13;
	wire [WIDTH*2-1+1:0] tmp01_3_14;
	wire [WIDTH*2-1+1:0] tmp01_3_15;
	wire [WIDTH*2-1+1:0] tmp01_3_16;
	wire [WIDTH*2-1+1:0] tmp01_3_17;
	wire [WIDTH*2-1+1:0] tmp01_3_18;
	wire [WIDTH*2-1+1:0] tmp01_3_19;
	wire [WIDTH*2-1+1:0] tmp01_3_20;
	wire [WIDTH*2-1+1:0] tmp01_3_21;
	wire [WIDTH*2-1+1:0] tmp01_3_22;
	wire [WIDTH*2-1+1:0] tmp01_3_23;
	wire [WIDTH*2-1+1:0] tmp01_3_24;
	wire [WIDTH*2-1+1:0] tmp01_3_25;
	wire [WIDTH*2-1+1:0] tmp01_3_26;
	wire [WIDTH*2-1+1:0] tmp01_3_27;
	wire [WIDTH*2-1+1:0] tmp01_3_28;
	wire [WIDTH*2-1+1:0] tmp01_3_29;
	wire [WIDTH*2-1+1:0] tmp01_3_30;
	wire [WIDTH*2-1+1:0] tmp01_3_31;
	wire [WIDTH*2-1+1:0] tmp01_3_32;
	wire [WIDTH*2-1+1:0] tmp01_3_33;
	wire [WIDTH*2-1+1:0] tmp01_3_34;
	wire [WIDTH*2-1+1:0] tmp01_3_35;
	wire [WIDTH*2-1+1:0] tmp01_3_36;
	wire [WIDTH*2-1+1:0] tmp01_3_37;
	wire [WIDTH*2-1+1:0] tmp01_3_38;
	wire [WIDTH*2-1+1:0] tmp01_3_39;
	wire [WIDTH*2-1+1:0] tmp01_3_40;
	wire [WIDTH*2-1+1:0] tmp01_3_41;
	wire [WIDTH*2-1+1:0] tmp01_3_42;
	wire [WIDTH*2-1+1:0] tmp01_3_43;
	wire [WIDTH*2-1+1:0] tmp01_3_44;
	wire [WIDTH*2-1+1:0] tmp01_3_45;
	wire [WIDTH*2-1+1:0] tmp01_3_46;
	wire [WIDTH*2-1+1:0] tmp01_3_47;
	wire [WIDTH*2-1+1:0] tmp01_3_48;
	wire [WIDTH*2-1+1:0] tmp01_3_49;
	wire [WIDTH*2-1+1:0] tmp01_3_50;
	wire [WIDTH*2-1+1:0] tmp01_3_51;
	wire [WIDTH*2-1+1:0] tmp01_3_52;
	wire [WIDTH*2-1+1:0] tmp01_3_53;
	wire [WIDTH*2-1+1:0] tmp01_3_54;
	wire [WIDTH*2-1+1:0] tmp01_3_55;
	wire [WIDTH*2-1+1:0] tmp01_3_56;
	wire [WIDTH*2-1+1:0] tmp01_3_57;
	wire [WIDTH*2-1+1:0] tmp01_3_58;
	wire [WIDTH*2-1+1:0] tmp01_3_59;
	wire [WIDTH*2-1+1:0] tmp01_3_60;
	wire [WIDTH*2-1+1:0] tmp01_3_61;
	wire [WIDTH*2-1+1:0] tmp01_3_62;
	wire [WIDTH*2-1+1:0] tmp01_3_63;
	wire [WIDTH*2-1+1:0] tmp01_3_64;
	wire [WIDTH*2-1+1:0] tmp01_3_65;
	wire [WIDTH*2-1+1:0] tmp01_3_66;
	wire [WIDTH*2-1+1:0] tmp01_3_67;
	wire [WIDTH*2-1+1:0] tmp01_3_68;
	wire [WIDTH*2-1+1:0] tmp01_3_69;
	wire [WIDTH*2-1+1:0] tmp01_3_70;
	wire [WIDTH*2-1+1:0] tmp01_3_71;
	wire [WIDTH*2-1+1:0] tmp01_3_72;
	wire [WIDTH*2-1+1:0] tmp01_3_73;
	wire [WIDTH*2-1+1:0] tmp01_3_74;
	wire [WIDTH*2-1+1:0] tmp01_3_75;
	wire [WIDTH*2-1+1:0] tmp01_3_76;
	wire [WIDTH*2-1+1:0] tmp01_3_77;
	wire [WIDTH*2-1+1:0] tmp01_3_78;
	wire [WIDTH*2-1+1:0] tmp01_3_79;
	wire [WIDTH*2-1+1:0] tmp01_3_80;
	wire [WIDTH*2-1+1:0] tmp01_3_81;
	wire [WIDTH*2-1+1:0] tmp01_3_82;
	wire [WIDTH*2-1+1:0] tmp01_3_83;
	wire [WIDTH*2-1+1:0] tmp01_4_0;
	wire [WIDTH*2-1+1:0] tmp01_4_1;
	wire [WIDTH*2-1+1:0] tmp01_4_2;
	wire [WIDTH*2-1+1:0] tmp01_4_3;
	wire [WIDTH*2-1+1:0] tmp01_4_4;
	wire [WIDTH*2-1+1:0] tmp01_4_5;
	wire [WIDTH*2-1+1:0] tmp01_4_6;
	wire [WIDTH*2-1+1:0] tmp01_4_7;
	wire [WIDTH*2-1+1:0] tmp01_4_8;
	wire [WIDTH*2-1+1:0] tmp01_4_9;
	wire [WIDTH*2-1+1:0] tmp01_4_10;
	wire [WIDTH*2-1+1:0] tmp01_4_11;
	wire [WIDTH*2-1+1:0] tmp01_4_12;
	wire [WIDTH*2-1+1:0] tmp01_4_13;
	wire [WIDTH*2-1+1:0] tmp01_4_14;
	wire [WIDTH*2-1+1:0] tmp01_4_15;
	wire [WIDTH*2-1+1:0] tmp01_4_16;
	wire [WIDTH*2-1+1:0] tmp01_4_17;
	wire [WIDTH*2-1+1:0] tmp01_4_18;
	wire [WIDTH*2-1+1:0] tmp01_4_19;
	wire [WIDTH*2-1+1:0] tmp01_4_20;
	wire [WIDTH*2-1+1:0] tmp01_4_21;
	wire [WIDTH*2-1+1:0] tmp01_4_22;
	wire [WIDTH*2-1+1:0] tmp01_4_23;
	wire [WIDTH*2-1+1:0] tmp01_4_24;
	wire [WIDTH*2-1+1:0] tmp01_4_25;
	wire [WIDTH*2-1+1:0] tmp01_4_26;
	wire [WIDTH*2-1+1:0] tmp01_4_27;
	wire [WIDTH*2-1+1:0] tmp01_4_28;
	wire [WIDTH*2-1+1:0] tmp01_4_29;
	wire [WIDTH*2-1+1:0] tmp01_4_30;
	wire [WIDTH*2-1+1:0] tmp01_4_31;
	wire [WIDTH*2-1+1:0] tmp01_4_32;
	wire [WIDTH*2-1+1:0] tmp01_4_33;
	wire [WIDTH*2-1+1:0] tmp01_4_34;
	wire [WIDTH*2-1+1:0] tmp01_4_35;
	wire [WIDTH*2-1+1:0] tmp01_4_36;
	wire [WIDTH*2-1+1:0] tmp01_4_37;
	wire [WIDTH*2-1+1:0] tmp01_4_38;
	wire [WIDTH*2-1+1:0] tmp01_4_39;
	wire [WIDTH*2-1+1:0] tmp01_4_40;
	wire [WIDTH*2-1+1:0] tmp01_4_41;
	wire [WIDTH*2-1+1:0] tmp01_4_42;
	wire [WIDTH*2-1+1:0] tmp01_4_43;
	wire [WIDTH*2-1+1:0] tmp01_4_44;
	wire [WIDTH*2-1+1:0] tmp01_4_45;
	wire [WIDTH*2-1+1:0] tmp01_4_46;
	wire [WIDTH*2-1+1:0] tmp01_4_47;
	wire [WIDTH*2-1+1:0] tmp01_4_48;
	wire [WIDTH*2-1+1:0] tmp01_4_49;
	wire [WIDTH*2-1+1:0] tmp01_4_50;
	wire [WIDTH*2-1+1:0] tmp01_4_51;
	wire [WIDTH*2-1+1:0] tmp01_4_52;
	wire [WIDTH*2-1+1:0] tmp01_4_53;
	wire [WIDTH*2-1+1:0] tmp01_4_54;
	wire [WIDTH*2-1+1:0] tmp01_4_55;
	wire [WIDTH*2-1+1:0] tmp01_4_56;
	wire [WIDTH*2-1+1:0] tmp01_4_57;
	wire [WIDTH*2-1+1:0] tmp01_4_58;
	wire [WIDTH*2-1+1:0] tmp01_4_59;
	wire [WIDTH*2-1+1:0] tmp01_4_60;
	wire [WIDTH*2-1+1:0] tmp01_4_61;
	wire [WIDTH*2-1+1:0] tmp01_4_62;
	wire [WIDTH*2-1+1:0] tmp01_4_63;
	wire [WIDTH*2-1+1:0] tmp01_4_64;
	wire [WIDTH*2-1+1:0] tmp01_4_65;
	wire [WIDTH*2-1+1:0] tmp01_4_66;
	wire [WIDTH*2-1+1:0] tmp01_4_67;
	wire [WIDTH*2-1+1:0] tmp01_4_68;
	wire [WIDTH*2-1+1:0] tmp01_4_69;
	wire [WIDTH*2-1+1:0] tmp01_4_70;
	wire [WIDTH*2-1+1:0] tmp01_4_71;
	wire [WIDTH*2-1+1:0] tmp01_4_72;
	wire [WIDTH*2-1+1:0] tmp01_4_73;
	wire [WIDTH*2-1+1:0] tmp01_4_74;
	wire [WIDTH*2-1+1:0] tmp01_4_75;
	wire [WIDTH*2-1+1:0] tmp01_4_76;
	wire [WIDTH*2-1+1:0] tmp01_4_77;
	wire [WIDTH*2-1+1:0] tmp01_4_78;
	wire [WIDTH*2-1+1:0] tmp01_4_79;
	wire [WIDTH*2-1+1:0] tmp01_4_80;
	wire [WIDTH*2-1+1:0] tmp01_4_81;
	wire [WIDTH*2-1+1:0] tmp01_4_82;
	wire [WIDTH*2-1+1:0] tmp01_4_83;
	wire [WIDTH*2-1+1:0] tmp01_5_0;
	wire [WIDTH*2-1+1:0] tmp01_5_1;
	wire [WIDTH*2-1+1:0] tmp01_5_2;
	wire [WIDTH*2-1+1:0] tmp01_5_3;
	wire [WIDTH*2-1+1:0] tmp01_5_4;
	wire [WIDTH*2-1+1:0] tmp01_5_5;
	wire [WIDTH*2-1+1:0] tmp01_5_6;
	wire [WIDTH*2-1+1:0] tmp01_5_7;
	wire [WIDTH*2-1+1:0] tmp01_5_8;
	wire [WIDTH*2-1+1:0] tmp01_5_9;
	wire [WIDTH*2-1+1:0] tmp01_5_10;
	wire [WIDTH*2-1+1:0] tmp01_5_11;
	wire [WIDTH*2-1+1:0] tmp01_5_12;
	wire [WIDTH*2-1+1:0] tmp01_5_13;
	wire [WIDTH*2-1+1:0] tmp01_5_14;
	wire [WIDTH*2-1+1:0] tmp01_5_15;
	wire [WIDTH*2-1+1:0] tmp01_5_16;
	wire [WIDTH*2-1+1:0] tmp01_5_17;
	wire [WIDTH*2-1+1:0] tmp01_5_18;
	wire [WIDTH*2-1+1:0] tmp01_5_19;
	wire [WIDTH*2-1+1:0] tmp01_5_20;
	wire [WIDTH*2-1+1:0] tmp01_5_21;
	wire [WIDTH*2-1+1:0] tmp01_5_22;
	wire [WIDTH*2-1+1:0] tmp01_5_23;
	wire [WIDTH*2-1+1:0] tmp01_5_24;
	wire [WIDTH*2-1+1:0] tmp01_5_25;
	wire [WIDTH*2-1+1:0] tmp01_5_26;
	wire [WIDTH*2-1+1:0] tmp01_5_27;
	wire [WIDTH*2-1+1:0] tmp01_5_28;
	wire [WIDTH*2-1+1:0] tmp01_5_29;
	wire [WIDTH*2-1+1:0] tmp01_5_30;
	wire [WIDTH*2-1+1:0] tmp01_5_31;
	wire [WIDTH*2-1+1:0] tmp01_5_32;
	wire [WIDTH*2-1+1:0] tmp01_5_33;
	wire [WIDTH*2-1+1:0] tmp01_5_34;
	wire [WIDTH*2-1+1:0] tmp01_5_35;
	wire [WIDTH*2-1+1:0] tmp01_5_36;
	wire [WIDTH*2-1+1:0] tmp01_5_37;
	wire [WIDTH*2-1+1:0] tmp01_5_38;
	wire [WIDTH*2-1+1:0] tmp01_5_39;
	wire [WIDTH*2-1+1:0] tmp01_5_40;
	wire [WIDTH*2-1+1:0] tmp01_5_41;
	wire [WIDTH*2-1+1:0] tmp01_5_42;
	wire [WIDTH*2-1+1:0] tmp01_5_43;
	wire [WIDTH*2-1+1:0] tmp01_5_44;
	wire [WIDTH*2-1+1:0] tmp01_5_45;
	wire [WIDTH*2-1+1:0] tmp01_5_46;
	wire [WIDTH*2-1+1:0] tmp01_5_47;
	wire [WIDTH*2-1+1:0] tmp01_5_48;
	wire [WIDTH*2-1+1:0] tmp01_5_49;
	wire [WIDTH*2-1+1:0] tmp01_5_50;
	wire [WIDTH*2-1+1:0] tmp01_5_51;
	wire [WIDTH*2-1+1:0] tmp01_5_52;
	wire [WIDTH*2-1+1:0] tmp01_5_53;
	wire [WIDTH*2-1+1:0] tmp01_5_54;
	wire [WIDTH*2-1+1:0] tmp01_5_55;
	wire [WIDTH*2-1+1:0] tmp01_5_56;
	wire [WIDTH*2-1+1:0] tmp01_5_57;
	wire [WIDTH*2-1+1:0] tmp01_5_58;
	wire [WIDTH*2-1+1:0] tmp01_5_59;
	wire [WIDTH*2-1+1:0] tmp01_5_60;
	wire [WIDTH*2-1+1:0] tmp01_5_61;
	wire [WIDTH*2-1+1:0] tmp01_5_62;
	wire [WIDTH*2-1+1:0] tmp01_5_63;
	wire [WIDTH*2-1+1:0] tmp01_5_64;
	wire [WIDTH*2-1+1:0] tmp01_5_65;
	wire [WIDTH*2-1+1:0] tmp01_5_66;
	wire [WIDTH*2-1+1:0] tmp01_5_67;
	wire [WIDTH*2-1+1:0] tmp01_5_68;
	wire [WIDTH*2-1+1:0] tmp01_5_69;
	wire [WIDTH*2-1+1:0] tmp01_5_70;
	wire [WIDTH*2-1+1:0] tmp01_5_71;
	wire [WIDTH*2-1+1:0] tmp01_5_72;
	wire [WIDTH*2-1+1:0] tmp01_5_73;
	wire [WIDTH*2-1+1:0] tmp01_5_74;
	wire [WIDTH*2-1+1:0] tmp01_5_75;
	wire [WIDTH*2-1+1:0] tmp01_5_76;
	wire [WIDTH*2-1+1:0] tmp01_5_77;
	wire [WIDTH*2-1+1:0] tmp01_5_78;
	wire [WIDTH*2-1+1:0] tmp01_5_79;
	wire [WIDTH*2-1+1:0] tmp01_5_80;
	wire [WIDTH*2-1+1:0] tmp01_5_81;
	wire [WIDTH*2-1+1:0] tmp01_5_82;
	wire [WIDTH*2-1+1:0] tmp01_5_83;
	wire [WIDTH*2-1+1:0] tmp01_6_0;
	wire [WIDTH*2-1+1:0] tmp01_6_1;
	wire [WIDTH*2-1+1:0] tmp01_6_2;
	wire [WIDTH*2-1+1:0] tmp01_6_3;
	wire [WIDTH*2-1+1:0] tmp01_6_4;
	wire [WIDTH*2-1+1:0] tmp01_6_5;
	wire [WIDTH*2-1+1:0] tmp01_6_6;
	wire [WIDTH*2-1+1:0] tmp01_6_7;
	wire [WIDTH*2-1+1:0] tmp01_6_8;
	wire [WIDTH*2-1+1:0] tmp01_6_9;
	wire [WIDTH*2-1+1:0] tmp01_6_10;
	wire [WIDTH*2-1+1:0] tmp01_6_11;
	wire [WIDTH*2-1+1:0] tmp01_6_12;
	wire [WIDTH*2-1+1:0] tmp01_6_13;
	wire [WIDTH*2-1+1:0] tmp01_6_14;
	wire [WIDTH*2-1+1:0] tmp01_6_15;
	wire [WIDTH*2-1+1:0] tmp01_6_16;
	wire [WIDTH*2-1+1:0] tmp01_6_17;
	wire [WIDTH*2-1+1:0] tmp01_6_18;
	wire [WIDTH*2-1+1:0] tmp01_6_19;
	wire [WIDTH*2-1+1:0] tmp01_6_20;
	wire [WIDTH*2-1+1:0] tmp01_6_21;
	wire [WIDTH*2-1+1:0] tmp01_6_22;
	wire [WIDTH*2-1+1:0] tmp01_6_23;
	wire [WIDTH*2-1+1:0] tmp01_6_24;
	wire [WIDTH*2-1+1:0] tmp01_6_25;
	wire [WIDTH*2-1+1:0] tmp01_6_26;
	wire [WIDTH*2-1+1:0] tmp01_6_27;
	wire [WIDTH*2-1+1:0] tmp01_6_28;
	wire [WIDTH*2-1+1:0] tmp01_6_29;
	wire [WIDTH*2-1+1:0] tmp01_6_30;
	wire [WIDTH*2-1+1:0] tmp01_6_31;
	wire [WIDTH*2-1+1:0] tmp01_6_32;
	wire [WIDTH*2-1+1:0] tmp01_6_33;
	wire [WIDTH*2-1+1:0] tmp01_6_34;
	wire [WIDTH*2-1+1:0] tmp01_6_35;
	wire [WIDTH*2-1+1:0] tmp01_6_36;
	wire [WIDTH*2-1+1:0] tmp01_6_37;
	wire [WIDTH*2-1+1:0] tmp01_6_38;
	wire [WIDTH*2-1+1:0] tmp01_6_39;
	wire [WIDTH*2-1+1:0] tmp01_6_40;
	wire [WIDTH*2-1+1:0] tmp01_6_41;
	wire [WIDTH*2-1+1:0] tmp01_6_42;
	wire [WIDTH*2-1+1:0] tmp01_6_43;
	wire [WIDTH*2-1+1:0] tmp01_6_44;
	wire [WIDTH*2-1+1:0] tmp01_6_45;
	wire [WIDTH*2-1+1:0] tmp01_6_46;
	wire [WIDTH*2-1+1:0] tmp01_6_47;
	wire [WIDTH*2-1+1:0] tmp01_6_48;
	wire [WIDTH*2-1+1:0] tmp01_6_49;
	wire [WIDTH*2-1+1:0] tmp01_6_50;
	wire [WIDTH*2-1+1:0] tmp01_6_51;
	wire [WIDTH*2-1+1:0] tmp01_6_52;
	wire [WIDTH*2-1+1:0] tmp01_6_53;
	wire [WIDTH*2-1+1:0] tmp01_6_54;
	wire [WIDTH*2-1+1:0] tmp01_6_55;
	wire [WIDTH*2-1+1:0] tmp01_6_56;
	wire [WIDTH*2-1+1:0] tmp01_6_57;
	wire [WIDTH*2-1+1:0] tmp01_6_58;
	wire [WIDTH*2-1+1:0] tmp01_6_59;
	wire [WIDTH*2-1+1:0] tmp01_6_60;
	wire [WIDTH*2-1+1:0] tmp01_6_61;
	wire [WIDTH*2-1+1:0] tmp01_6_62;
	wire [WIDTH*2-1+1:0] tmp01_6_63;
	wire [WIDTH*2-1+1:0] tmp01_6_64;
	wire [WIDTH*2-1+1:0] tmp01_6_65;
	wire [WIDTH*2-1+1:0] tmp01_6_66;
	wire [WIDTH*2-1+1:0] tmp01_6_67;
	wire [WIDTH*2-1+1:0] tmp01_6_68;
	wire [WIDTH*2-1+1:0] tmp01_6_69;
	wire [WIDTH*2-1+1:0] tmp01_6_70;
	wire [WIDTH*2-1+1:0] tmp01_6_71;
	wire [WIDTH*2-1+1:0] tmp01_6_72;
	wire [WIDTH*2-1+1:0] tmp01_6_73;
	wire [WIDTH*2-1+1:0] tmp01_6_74;
	wire [WIDTH*2-1+1:0] tmp01_6_75;
	wire [WIDTH*2-1+1:0] tmp01_6_76;
	wire [WIDTH*2-1+1:0] tmp01_6_77;
	wire [WIDTH*2-1+1:0] tmp01_6_78;
	wire [WIDTH*2-1+1:0] tmp01_6_79;
	wire [WIDTH*2-1+1:0] tmp01_6_80;
	wire [WIDTH*2-1+1:0] tmp01_6_81;
	wire [WIDTH*2-1+1:0] tmp01_6_82;
	wire [WIDTH*2-1+1:0] tmp01_6_83;
	wire [WIDTH*2-1+1:0] tmp01_7_0;
	wire [WIDTH*2-1+1:0] tmp01_7_1;
	wire [WIDTH*2-1+1:0] tmp01_7_2;
	wire [WIDTH*2-1+1:0] tmp01_7_3;
	wire [WIDTH*2-1+1:0] tmp01_7_4;
	wire [WIDTH*2-1+1:0] tmp01_7_5;
	wire [WIDTH*2-1+1:0] tmp01_7_6;
	wire [WIDTH*2-1+1:0] tmp01_7_7;
	wire [WIDTH*2-1+1:0] tmp01_7_8;
	wire [WIDTH*2-1+1:0] tmp01_7_9;
	wire [WIDTH*2-1+1:0] tmp01_7_10;
	wire [WIDTH*2-1+1:0] tmp01_7_11;
	wire [WIDTH*2-1+1:0] tmp01_7_12;
	wire [WIDTH*2-1+1:0] tmp01_7_13;
	wire [WIDTH*2-1+1:0] tmp01_7_14;
	wire [WIDTH*2-1+1:0] tmp01_7_15;
	wire [WIDTH*2-1+1:0] tmp01_7_16;
	wire [WIDTH*2-1+1:0] tmp01_7_17;
	wire [WIDTH*2-1+1:0] tmp01_7_18;
	wire [WIDTH*2-1+1:0] tmp01_7_19;
	wire [WIDTH*2-1+1:0] tmp01_7_20;
	wire [WIDTH*2-1+1:0] tmp01_7_21;
	wire [WIDTH*2-1+1:0] tmp01_7_22;
	wire [WIDTH*2-1+1:0] tmp01_7_23;
	wire [WIDTH*2-1+1:0] tmp01_7_24;
	wire [WIDTH*2-1+1:0] tmp01_7_25;
	wire [WIDTH*2-1+1:0] tmp01_7_26;
	wire [WIDTH*2-1+1:0] tmp01_7_27;
	wire [WIDTH*2-1+1:0] tmp01_7_28;
	wire [WIDTH*2-1+1:0] tmp01_7_29;
	wire [WIDTH*2-1+1:0] tmp01_7_30;
	wire [WIDTH*2-1+1:0] tmp01_7_31;
	wire [WIDTH*2-1+1:0] tmp01_7_32;
	wire [WIDTH*2-1+1:0] tmp01_7_33;
	wire [WIDTH*2-1+1:0] tmp01_7_34;
	wire [WIDTH*2-1+1:0] tmp01_7_35;
	wire [WIDTH*2-1+1:0] tmp01_7_36;
	wire [WIDTH*2-1+1:0] tmp01_7_37;
	wire [WIDTH*2-1+1:0] tmp01_7_38;
	wire [WIDTH*2-1+1:0] tmp01_7_39;
	wire [WIDTH*2-1+1:0] tmp01_7_40;
	wire [WIDTH*2-1+1:0] tmp01_7_41;
	wire [WIDTH*2-1+1:0] tmp01_7_42;
	wire [WIDTH*2-1+1:0] tmp01_7_43;
	wire [WIDTH*2-1+1:0] tmp01_7_44;
	wire [WIDTH*2-1+1:0] tmp01_7_45;
	wire [WIDTH*2-1+1:0] tmp01_7_46;
	wire [WIDTH*2-1+1:0] tmp01_7_47;
	wire [WIDTH*2-1+1:0] tmp01_7_48;
	wire [WIDTH*2-1+1:0] tmp01_7_49;
	wire [WIDTH*2-1+1:0] tmp01_7_50;
	wire [WIDTH*2-1+1:0] tmp01_7_51;
	wire [WIDTH*2-1+1:0] tmp01_7_52;
	wire [WIDTH*2-1+1:0] tmp01_7_53;
	wire [WIDTH*2-1+1:0] tmp01_7_54;
	wire [WIDTH*2-1+1:0] tmp01_7_55;
	wire [WIDTH*2-1+1:0] tmp01_7_56;
	wire [WIDTH*2-1+1:0] tmp01_7_57;
	wire [WIDTH*2-1+1:0] tmp01_7_58;
	wire [WIDTH*2-1+1:0] tmp01_7_59;
	wire [WIDTH*2-1+1:0] tmp01_7_60;
	wire [WIDTH*2-1+1:0] tmp01_7_61;
	wire [WIDTH*2-1+1:0] tmp01_7_62;
	wire [WIDTH*2-1+1:0] tmp01_7_63;
	wire [WIDTH*2-1+1:0] tmp01_7_64;
	wire [WIDTH*2-1+1:0] tmp01_7_65;
	wire [WIDTH*2-1+1:0] tmp01_7_66;
	wire [WIDTH*2-1+1:0] tmp01_7_67;
	wire [WIDTH*2-1+1:0] tmp01_7_68;
	wire [WIDTH*2-1+1:0] tmp01_7_69;
	wire [WIDTH*2-1+1:0] tmp01_7_70;
	wire [WIDTH*2-1+1:0] tmp01_7_71;
	wire [WIDTH*2-1+1:0] tmp01_7_72;
	wire [WIDTH*2-1+1:0] tmp01_7_73;
	wire [WIDTH*2-1+1:0] tmp01_7_74;
	wire [WIDTH*2-1+1:0] tmp01_7_75;
	wire [WIDTH*2-1+1:0] tmp01_7_76;
	wire [WIDTH*2-1+1:0] tmp01_7_77;
	wire [WIDTH*2-1+1:0] tmp01_7_78;
	wire [WIDTH*2-1+1:0] tmp01_7_79;
	wire [WIDTH*2-1+1:0] tmp01_7_80;
	wire [WIDTH*2-1+1:0] tmp01_7_81;
	wire [WIDTH*2-1+1:0] tmp01_7_82;
	wire [WIDTH*2-1+1:0] tmp01_7_83;
	wire [WIDTH*2-1+1:0] tmp01_8_0;
	wire [WIDTH*2-1+1:0] tmp01_8_1;
	wire [WIDTH*2-1+1:0] tmp01_8_2;
	wire [WIDTH*2-1+1:0] tmp01_8_3;
	wire [WIDTH*2-1+1:0] tmp01_8_4;
	wire [WIDTH*2-1+1:0] tmp01_8_5;
	wire [WIDTH*2-1+1:0] tmp01_8_6;
	wire [WIDTH*2-1+1:0] tmp01_8_7;
	wire [WIDTH*2-1+1:0] tmp01_8_8;
	wire [WIDTH*2-1+1:0] tmp01_8_9;
	wire [WIDTH*2-1+1:0] tmp01_8_10;
	wire [WIDTH*2-1+1:0] tmp01_8_11;
	wire [WIDTH*2-1+1:0] tmp01_8_12;
	wire [WIDTH*2-1+1:0] tmp01_8_13;
	wire [WIDTH*2-1+1:0] tmp01_8_14;
	wire [WIDTH*2-1+1:0] tmp01_8_15;
	wire [WIDTH*2-1+1:0] tmp01_8_16;
	wire [WIDTH*2-1+1:0] tmp01_8_17;
	wire [WIDTH*2-1+1:0] tmp01_8_18;
	wire [WIDTH*2-1+1:0] tmp01_8_19;
	wire [WIDTH*2-1+1:0] tmp01_8_20;
	wire [WIDTH*2-1+1:0] tmp01_8_21;
	wire [WIDTH*2-1+1:0] tmp01_8_22;
	wire [WIDTH*2-1+1:0] tmp01_8_23;
	wire [WIDTH*2-1+1:0] tmp01_8_24;
	wire [WIDTH*2-1+1:0] tmp01_8_25;
	wire [WIDTH*2-1+1:0] tmp01_8_26;
	wire [WIDTH*2-1+1:0] tmp01_8_27;
	wire [WIDTH*2-1+1:0] tmp01_8_28;
	wire [WIDTH*2-1+1:0] tmp01_8_29;
	wire [WIDTH*2-1+1:0] tmp01_8_30;
	wire [WIDTH*2-1+1:0] tmp01_8_31;
	wire [WIDTH*2-1+1:0] tmp01_8_32;
	wire [WIDTH*2-1+1:0] tmp01_8_33;
	wire [WIDTH*2-1+1:0] tmp01_8_34;
	wire [WIDTH*2-1+1:0] tmp01_8_35;
	wire [WIDTH*2-1+1:0] tmp01_8_36;
	wire [WIDTH*2-1+1:0] tmp01_8_37;
	wire [WIDTH*2-1+1:0] tmp01_8_38;
	wire [WIDTH*2-1+1:0] tmp01_8_39;
	wire [WIDTH*2-1+1:0] tmp01_8_40;
	wire [WIDTH*2-1+1:0] tmp01_8_41;
	wire [WIDTH*2-1+1:0] tmp01_8_42;
	wire [WIDTH*2-1+1:0] tmp01_8_43;
	wire [WIDTH*2-1+1:0] tmp01_8_44;
	wire [WIDTH*2-1+1:0] tmp01_8_45;
	wire [WIDTH*2-1+1:0] tmp01_8_46;
	wire [WIDTH*2-1+1:0] tmp01_8_47;
	wire [WIDTH*2-1+1:0] tmp01_8_48;
	wire [WIDTH*2-1+1:0] tmp01_8_49;
	wire [WIDTH*2-1+1:0] tmp01_8_50;
	wire [WIDTH*2-1+1:0] tmp01_8_51;
	wire [WIDTH*2-1+1:0] tmp01_8_52;
	wire [WIDTH*2-1+1:0] tmp01_8_53;
	wire [WIDTH*2-1+1:0] tmp01_8_54;
	wire [WIDTH*2-1+1:0] tmp01_8_55;
	wire [WIDTH*2-1+1:0] tmp01_8_56;
	wire [WIDTH*2-1+1:0] tmp01_8_57;
	wire [WIDTH*2-1+1:0] tmp01_8_58;
	wire [WIDTH*2-1+1:0] tmp01_8_59;
	wire [WIDTH*2-1+1:0] tmp01_8_60;
	wire [WIDTH*2-1+1:0] tmp01_8_61;
	wire [WIDTH*2-1+1:0] tmp01_8_62;
	wire [WIDTH*2-1+1:0] tmp01_8_63;
	wire [WIDTH*2-1+1:0] tmp01_8_64;
	wire [WIDTH*2-1+1:0] tmp01_8_65;
	wire [WIDTH*2-1+1:0] tmp01_8_66;
	wire [WIDTH*2-1+1:0] tmp01_8_67;
	wire [WIDTH*2-1+1:0] tmp01_8_68;
	wire [WIDTH*2-1+1:0] tmp01_8_69;
	wire [WIDTH*2-1+1:0] tmp01_8_70;
	wire [WIDTH*2-1+1:0] tmp01_8_71;
	wire [WIDTH*2-1+1:0] tmp01_8_72;
	wire [WIDTH*2-1+1:0] tmp01_8_73;
	wire [WIDTH*2-1+1:0] tmp01_8_74;
	wire [WIDTH*2-1+1:0] tmp01_8_75;
	wire [WIDTH*2-1+1:0] tmp01_8_76;
	wire [WIDTH*2-1+1:0] tmp01_8_77;
	wire [WIDTH*2-1+1:0] tmp01_8_78;
	wire [WIDTH*2-1+1:0] tmp01_8_79;
	wire [WIDTH*2-1+1:0] tmp01_8_80;
	wire [WIDTH*2-1+1:0] tmp01_8_81;
	wire [WIDTH*2-1+1:0] tmp01_8_82;
	wire [WIDTH*2-1+1:0] tmp01_8_83;
	wire [WIDTH*2-1+1:0] tmp01_9_0;
	wire [WIDTH*2-1+1:0] tmp01_9_1;
	wire [WIDTH*2-1+1:0] tmp01_9_2;
	wire [WIDTH*2-1+1:0] tmp01_9_3;
	wire [WIDTH*2-1+1:0] tmp01_9_4;
	wire [WIDTH*2-1+1:0] tmp01_9_5;
	wire [WIDTH*2-1+1:0] tmp01_9_6;
	wire [WIDTH*2-1+1:0] tmp01_9_7;
	wire [WIDTH*2-1+1:0] tmp01_9_8;
	wire [WIDTH*2-1+1:0] tmp01_9_9;
	wire [WIDTH*2-1+1:0] tmp01_9_10;
	wire [WIDTH*2-1+1:0] tmp01_9_11;
	wire [WIDTH*2-1+1:0] tmp01_9_12;
	wire [WIDTH*2-1+1:0] tmp01_9_13;
	wire [WIDTH*2-1+1:0] tmp01_9_14;
	wire [WIDTH*2-1+1:0] tmp01_9_15;
	wire [WIDTH*2-1+1:0] tmp01_9_16;
	wire [WIDTH*2-1+1:0] tmp01_9_17;
	wire [WIDTH*2-1+1:0] tmp01_9_18;
	wire [WIDTH*2-1+1:0] tmp01_9_19;
	wire [WIDTH*2-1+1:0] tmp01_9_20;
	wire [WIDTH*2-1+1:0] tmp01_9_21;
	wire [WIDTH*2-1+1:0] tmp01_9_22;
	wire [WIDTH*2-1+1:0] tmp01_9_23;
	wire [WIDTH*2-1+1:0] tmp01_9_24;
	wire [WIDTH*2-1+1:0] tmp01_9_25;
	wire [WIDTH*2-1+1:0] tmp01_9_26;
	wire [WIDTH*2-1+1:0] tmp01_9_27;
	wire [WIDTH*2-1+1:0] tmp01_9_28;
	wire [WIDTH*2-1+1:0] tmp01_9_29;
	wire [WIDTH*2-1+1:0] tmp01_9_30;
	wire [WIDTH*2-1+1:0] tmp01_9_31;
	wire [WIDTH*2-1+1:0] tmp01_9_32;
	wire [WIDTH*2-1+1:0] tmp01_9_33;
	wire [WIDTH*2-1+1:0] tmp01_9_34;
	wire [WIDTH*2-1+1:0] tmp01_9_35;
	wire [WIDTH*2-1+1:0] tmp01_9_36;
	wire [WIDTH*2-1+1:0] tmp01_9_37;
	wire [WIDTH*2-1+1:0] tmp01_9_38;
	wire [WIDTH*2-1+1:0] tmp01_9_39;
	wire [WIDTH*2-1+1:0] tmp01_9_40;
	wire [WIDTH*2-1+1:0] tmp01_9_41;
	wire [WIDTH*2-1+1:0] tmp01_9_42;
	wire [WIDTH*2-1+1:0] tmp01_9_43;
	wire [WIDTH*2-1+1:0] tmp01_9_44;
	wire [WIDTH*2-1+1:0] tmp01_9_45;
	wire [WIDTH*2-1+1:0] tmp01_9_46;
	wire [WIDTH*2-1+1:0] tmp01_9_47;
	wire [WIDTH*2-1+1:0] tmp01_9_48;
	wire [WIDTH*2-1+1:0] tmp01_9_49;
	wire [WIDTH*2-1+1:0] tmp01_9_50;
	wire [WIDTH*2-1+1:0] tmp01_9_51;
	wire [WIDTH*2-1+1:0] tmp01_9_52;
	wire [WIDTH*2-1+1:0] tmp01_9_53;
	wire [WIDTH*2-1+1:0] tmp01_9_54;
	wire [WIDTH*2-1+1:0] tmp01_9_55;
	wire [WIDTH*2-1+1:0] tmp01_9_56;
	wire [WIDTH*2-1+1:0] tmp01_9_57;
	wire [WIDTH*2-1+1:0] tmp01_9_58;
	wire [WIDTH*2-1+1:0] tmp01_9_59;
	wire [WIDTH*2-1+1:0] tmp01_9_60;
	wire [WIDTH*2-1+1:0] tmp01_9_61;
	wire [WIDTH*2-1+1:0] tmp01_9_62;
	wire [WIDTH*2-1+1:0] tmp01_9_63;
	wire [WIDTH*2-1+1:0] tmp01_9_64;
	wire [WIDTH*2-1+1:0] tmp01_9_65;
	wire [WIDTH*2-1+1:0] tmp01_9_66;
	wire [WIDTH*2-1+1:0] tmp01_9_67;
	wire [WIDTH*2-1+1:0] tmp01_9_68;
	wire [WIDTH*2-1+1:0] tmp01_9_69;
	wire [WIDTH*2-1+1:0] tmp01_9_70;
	wire [WIDTH*2-1+1:0] tmp01_9_71;
	wire [WIDTH*2-1+1:0] tmp01_9_72;
	wire [WIDTH*2-1+1:0] tmp01_9_73;
	wire [WIDTH*2-1+1:0] tmp01_9_74;
	wire [WIDTH*2-1+1:0] tmp01_9_75;
	wire [WIDTH*2-1+1:0] tmp01_9_76;
	wire [WIDTH*2-1+1:0] tmp01_9_77;
	wire [WIDTH*2-1+1:0] tmp01_9_78;
	wire [WIDTH*2-1+1:0] tmp01_9_79;
	wire [WIDTH*2-1+1:0] tmp01_9_80;
	wire [WIDTH*2-1+1:0] tmp01_9_81;
	wire [WIDTH*2-1+1:0] tmp01_9_82;
	wire [WIDTH*2-1+1:0] tmp01_9_83;
	wire [WIDTH*2-1+1:0] tmp01_10_0;
	wire [WIDTH*2-1+1:0] tmp01_10_1;
	wire [WIDTH*2-1+1:0] tmp01_10_2;
	wire [WIDTH*2-1+1:0] tmp01_10_3;
	wire [WIDTH*2-1+1:0] tmp01_10_4;
	wire [WIDTH*2-1+1:0] tmp01_10_5;
	wire [WIDTH*2-1+1:0] tmp01_10_6;
	wire [WIDTH*2-1+1:0] tmp01_10_7;
	wire [WIDTH*2-1+1:0] tmp01_10_8;
	wire [WIDTH*2-1+1:0] tmp01_10_9;
	wire [WIDTH*2-1+1:0] tmp01_10_10;
	wire [WIDTH*2-1+1:0] tmp01_10_11;
	wire [WIDTH*2-1+1:0] tmp01_10_12;
	wire [WIDTH*2-1+1:0] tmp01_10_13;
	wire [WIDTH*2-1+1:0] tmp01_10_14;
	wire [WIDTH*2-1+1:0] tmp01_10_15;
	wire [WIDTH*2-1+1:0] tmp01_10_16;
	wire [WIDTH*2-1+1:0] tmp01_10_17;
	wire [WIDTH*2-1+1:0] tmp01_10_18;
	wire [WIDTH*2-1+1:0] tmp01_10_19;
	wire [WIDTH*2-1+1:0] tmp01_10_20;
	wire [WIDTH*2-1+1:0] tmp01_10_21;
	wire [WIDTH*2-1+1:0] tmp01_10_22;
	wire [WIDTH*2-1+1:0] tmp01_10_23;
	wire [WIDTH*2-1+1:0] tmp01_10_24;
	wire [WIDTH*2-1+1:0] tmp01_10_25;
	wire [WIDTH*2-1+1:0] tmp01_10_26;
	wire [WIDTH*2-1+1:0] tmp01_10_27;
	wire [WIDTH*2-1+1:0] tmp01_10_28;
	wire [WIDTH*2-1+1:0] tmp01_10_29;
	wire [WIDTH*2-1+1:0] tmp01_10_30;
	wire [WIDTH*2-1+1:0] tmp01_10_31;
	wire [WIDTH*2-1+1:0] tmp01_10_32;
	wire [WIDTH*2-1+1:0] tmp01_10_33;
	wire [WIDTH*2-1+1:0] tmp01_10_34;
	wire [WIDTH*2-1+1:0] tmp01_10_35;
	wire [WIDTH*2-1+1:0] tmp01_10_36;
	wire [WIDTH*2-1+1:0] tmp01_10_37;
	wire [WIDTH*2-1+1:0] tmp01_10_38;
	wire [WIDTH*2-1+1:0] tmp01_10_39;
	wire [WIDTH*2-1+1:0] tmp01_10_40;
	wire [WIDTH*2-1+1:0] tmp01_10_41;
	wire [WIDTH*2-1+1:0] tmp01_10_42;
	wire [WIDTH*2-1+1:0] tmp01_10_43;
	wire [WIDTH*2-1+1:0] tmp01_10_44;
	wire [WIDTH*2-1+1:0] tmp01_10_45;
	wire [WIDTH*2-1+1:0] tmp01_10_46;
	wire [WIDTH*2-1+1:0] tmp01_10_47;
	wire [WIDTH*2-1+1:0] tmp01_10_48;
	wire [WIDTH*2-1+1:0] tmp01_10_49;
	wire [WIDTH*2-1+1:0] tmp01_10_50;
	wire [WIDTH*2-1+1:0] tmp01_10_51;
	wire [WIDTH*2-1+1:0] tmp01_10_52;
	wire [WIDTH*2-1+1:0] tmp01_10_53;
	wire [WIDTH*2-1+1:0] tmp01_10_54;
	wire [WIDTH*2-1+1:0] tmp01_10_55;
	wire [WIDTH*2-1+1:0] tmp01_10_56;
	wire [WIDTH*2-1+1:0] tmp01_10_57;
	wire [WIDTH*2-1+1:0] tmp01_10_58;
	wire [WIDTH*2-1+1:0] tmp01_10_59;
	wire [WIDTH*2-1+1:0] tmp01_10_60;
	wire [WIDTH*2-1+1:0] tmp01_10_61;
	wire [WIDTH*2-1+1:0] tmp01_10_62;
	wire [WIDTH*2-1+1:0] tmp01_10_63;
	wire [WIDTH*2-1+1:0] tmp01_10_64;
	wire [WIDTH*2-1+1:0] tmp01_10_65;
	wire [WIDTH*2-1+1:0] tmp01_10_66;
	wire [WIDTH*2-1+1:0] tmp01_10_67;
	wire [WIDTH*2-1+1:0] tmp01_10_68;
	wire [WIDTH*2-1+1:0] tmp01_10_69;
	wire [WIDTH*2-1+1:0] tmp01_10_70;
	wire [WIDTH*2-1+1:0] tmp01_10_71;
	wire [WIDTH*2-1+1:0] tmp01_10_72;
	wire [WIDTH*2-1+1:0] tmp01_10_73;
	wire [WIDTH*2-1+1:0] tmp01_10_74;
	wire [WIDTH*2-1+1:0] tmp01_10_75;
	wire [WIDTH*2-1+1:0] tmp01_10_76;
	wire [WIDTH*2-1+1:0] tmp01_10_77;
	wire [WIDTH*2-1+1:0] tmp01_10_78;
	wire [WIDTH*2-1+1:0] tmp01_10_79;
	wire [WIDTH*2-1+1:0] tmp01_10_80;
	wire [WIDTH*2-1+1:0] tmp01_10_81;
	wire [WIDTH*2-1+1:0] tmp01_10_82;
	wire [WIDTH*2-1+1:0] tmp01_10_83;
	wire [WIDTH*2-1+1:0] tmp01_11_0;
	wire [WIDTH*2-1+1:0] tmp01_11_1;
	wire [WIDTH*2-1+1:0] tmp01_11_2;
	wire [WIDTH*2-1+1:0] tmp01_11_3;
	wire [WIDTH*2-1+1:0] tmp01_11_4;
	wire [WIDTH*2-1+1:0] tmp01_11_5;
	wire [WIDTH*2-1+1:0] tmp01_11_6;
	wire [WIDTH*2-1+1:0] tmp01_11_7;
	wire [WIDTH*2-1+1:0] tmp01_11_8;
	wire [WIDTH*2-1+1:0] tmp01_11_9;
	wire [WIDTH*2-1+1:0] tmp01_11_10;
	wire [WIDTH*2-1+1:0] tmp01_11_11;
	wire [WIDTH*2-1+1:0] tmp01_11_12;
	wire [WIDTH*2-1+1:0] tmp01_11_13;
	wire [WIDTH*2-1+1:0] tmp01_11_14;
	wire [WIDTH*2-1+1:0] tmp01_11_15;
	wire [WIDTH*2-1+1:0] tmp01_11_16;
	wire [WIDTH*2-1+1:0] tmp01_11_17;
	wire [WIDTH*2-1+1:0] tmp01_11_18;
	wire [WIDTH*2-1+1:0] tmp01_11_19;
	wire [WIDTH*2-1+1:0] tmp01_11_20;
	wire [WIDTH*2-1+1:0] tmp01_11_21;
	wire [WIDTH*2-1+1:0] tmp01_11_22;
	wire [WIDTH*2-1+1:0] tmp01_11_23;
	wire [WIDTH*2-1+1:0] tmp01_11_24;
	wire [WIDTH*2-1+1:0] tmp01_11_25;
	wire [WIDTH*2-1+1:0] tmp01_11_26;
	wire [WIDTH*2-1+1:0] tmp01_11_27;
	wire [WIDTH*2-1+1:0] tmp01_11_28;
	wire [WIDTH*2-1+1:0] tmp01_11_29;
	wire [WIDTH*2-1+1:0] tmp01_11_30;
	wire [WIDTH*2-1+1:0] tmp01_11_31;
	wire [WIDTH*2-1+1:0] tmp01_11_32;
	wire [WIDTH*2-1+1:0] tmp01_11_33;
	wire [WIDTH*2-1+1:0] tmp01_11_34;
	wire [WIDTH*2-1+1:0] tmp01_11_35;
	wire [WIDTH*2-1+1:0] tmp01_11_36;
	wire [WIDTH*2-1+1:0] tmp01_11_37;
	wire [WIDTH*2-1+1:0] tmp01_11_38;
	wire [WIDTH*2-1+1:0] tmp01_11_39;
	wire [WIDTH*2-1+1:0] tmp01_11_40;
	wire [WIDTH*2-1+1:0] tmp01_11_41;
	wire [WIDTH*2-1+1:0] tmp01_11_42;
	wire [WIDTH*2-1+1:0] tmp01_11_43;
	wire [WIDTH*2-1+1:0] tmp01_11_44;
	wire [WIDTH*2-1+1:0] tmp01_11_45;
	wire [WIDTH*2-1+1:0] tmp01_11_46;
	wire [WIDTH*2-1+1:0] tmp01_11_47;
	wire [WIDTH*2-1+1:0] tmp01_11_48;
	wire [WIDTH*2-1+1:0] tmp01_11_49;
	wire [WIDTH*2-1+1:0] tmp01_11_50;
	wire [WIDTH*2-1+1:0] tmp01_11_51;
	wire [WIDTH*2-1+1:0] tmp01_11_52;
	wire [WIDTH*2-1+1:0] tmp01_11_53;
	wire [WIDTH*2-1+1:0] tmp01_11_54;
	wire [WIDTH*2-1+1:0] tmp01_11_55;
	wire [WIDTH*2-1+1:0] tmp01_11_56;
	wire [WIDTH*2-1+1:0] tmp01_11_57;
	wire [WIDTH*2-1+1:0] tmp01_11_58;
	wire [WIDTH*2-1+1:0] tmp01_11_59;
	wire [WIDTH*2-1+1:0] tmp01_11_60;
	wire [WIDTH*2-1+1:0] tmp01_11_61;
	wire [WIDTH*2-1+1:0] tmp01_11_62;
	wire [WIDTH*2-1+1:0] tmp01_11_63;
	wire [WIDTH*2-1+1:0] tmp01_11_64;
	wire [WIDTH*2-1+1:0] tmp01_11_65;
	wire [WIDTH*2-1+1:0] tmp01_11_66;
	wire [WIDTH*2-1+1:0] tmp01_11_67;
	wire [WIDTH*2-1+1:0] tmp01_11_68;
	wire [WIDTH*2-1+1:0] tmp01_11_69;
	wire [WIDTH*2-1+1:0] tmp01_11_70;
	wire [WIDTH*2-1+1:0] tmp01_11_71;
	wire [WIDTH*2-1+1:0] tmp01_11_72;
	wire [WIDTH*2-1+1:0] tmp01_11_73;
	wire [WIDTH*2-1+1:0] tmp01_11_74;
	wire [WIDTH*2-1+1:0] tmp01_11_75;
	wire [WIDTH*2-1+1:0] tmp01_11_76;
	wire [WIDTH*2-1+1:0] tmp01_11_77;
	wire [WIDTH*2-1+1:0] tmp01_11_78;
	wire [WIDTH*2-1+1:0] tmp01_11_79;
	wire [WIDTH*2-1+1:0] tmp01_11_80;
	wire [WIDTH*2-1+1:0] tmp01_11_81;
	wire [WIDTH*2-1+1:0] tmp01_11_82;
	wire [WIDTH*2-1+1:0] tmp01_11_83;
	wire [WIDTH*2-1+1:0] tmp01_12_0;
	wire [WIDTH*2-1+1:0] tmp01_12_1;
	wire [WIDTH*2-1+1:0] tmp01_12_2;
	wire [WIDTH*2-1+1:0] tmp01_12_3;
	wire [WIDTH*2-1+1:0] tmp01_12_4;
	wire [WIDTH*2-1+1:0] tmp01_12_5;
	wire [WIDTH*2-1+1:0] tmp01_12_6;
	wire [WIDTH*2-1+1:0] tmp01_12_7;
	wire [WIDTH*2-1+1:0] tmp01_12_8;
	wire [WIDTH*2-1+1:0] tmp01_12_9;
	wire [WIDTH*2-1+1:0] tmp01_12_10;
	wire [WIDTH*2-1+1:0] tmp01_12_11;
	wire [WIDTH*2-1+1:0] tmp01_12_12;
	wire [WIDTH*2-1+1:0] tmp01_12_13;
	wire [WIDTH*2-1+1:0] tmp01_12_14;
	wire [WIDTH*2-1+1:0] tmp01_12_15;
	wire [WIDTH*2-1+1:0] tmp01_12_16;
	wire [WIDTH*2-1+1:0] tmp01_12_17;
	wire [WIDTH*2-1+1:0] tmp01_12_18;
	wire [WIDTH*2-1+1:0] tmp01_12_19;
	wire [WIDTH*2-1+1:0] tmp01_12_20;
	wire [WIDTH*2-1+1:0] tmp01_12_21;
	wire [WIDTH*2-1+1:0] tmp01_12_22;
	wire [WIDTH*2-1+1:0] tmp01_12_23;
	wire [WIDTH*2-1+1:0] tmp01_12_24;
	wire [WIDTH*2-1+1:0] tmp01_12_25;
	wire [WIDTH*2-1+1:0] tmp01_12_26;
	wire [WIDTH*2-1+1:0] tmp01_12_27;
	wire [WIDTH*2-1+1:0] tmp01_12_28;
	wire [WIDTH*2-1+1:0] tmp01_12_29;
	wire [WIDTH*2-1+1:0] tmp01_12_30;
	wire [WIDTH*2-1+1:0] tmp01_12_31;
	wire [WIDTH*2-1+1:0] tmp01_12_32;
	wire [WIDTH*2-1+1:0] tmp01_12_33;
	wire [WIDTH*2-1+1:0] tmp01_12_34;
	wire [WIDTH*2-1+1:0] tmp01_12_35;
	wire [WIDTH*2-1+1:0] tmp01_12_36;
	wire [WIDTH*2-1+1:0] tmp01_12_37;
	wire [WIDTH*2-1+1:0] tmp01_12_38;
	wire [WIDTH*2-1+1:0] tmp01_12_39;
	wire [WIDTH*2-1+1:0] tmp01_12_40;
	wire [WIDTH*2-1+1:0] tmp01_12_41;
	wire [WIDTH*2-1+1:0] tmp01_12_42;
	wire [WIDTH*2-1+1:0] tmp01_12_43;
	wire [WIDTH*2-1+1:0] tmp01_12_44;
	wire [WIDTH*2-1+1:0] tmp01_12_45;
	wire [WIDTH*2-1+1:0] tmp01_12_46;
	wire [WIDTH*2-1+1:0] tmp01_12_47;
	wire [WIDTH*2-1+1:0] tmp01_12_48;
	wire [WIDTH*2-1+1:0] tmp01_12_49;
	wire [WIDTH*2-1+1:0] tmp01_12_50;
	wire [WIDTH*2-1+1:0] tmp01_12_51;
	wire [WIDTH*2-1+1:0] tmp01_12_52;
	wire [WIDTH*2-1+1:0] tmp01_12_53;
	wire [WIDTH*2-1+1:0] tmp01_12_54;
	wire [WIDTH*2-1+1:0] tmp01_12_55;
	wire [WIDTH*2-1+1:0] tmp01_12_56;
	wire [WIDTH*2-1+1:0] tmp01_12_57;
	wire [WIDTH*2-1+1:0] tmp01_12_58;
	wire [WIDTH*2-1+1:0] tmp01_12_59;
	wire [WIDTH*2-1+1:0] tmp01_12_60;
	wire [WIDTH*2-1+1:0] tmp01_12_61;
	wire [WIDTH*2-1+1:0] tmp01_12_62;
	wire [WIDTH*2-1+1:0] tmp01_12_63;
	wire [WIDTH*2-1+1:0] tmp01_12_64;
	wire [WIDTH*2-1+1:0] tmp01_12_65;
	wire [WIDTH*2-1+1:0] tmp01_12_66;
	wire [WIDTH*2-1+1:0] tmp01_12_67;
	wire [WIDTH*2-1+1:0] tmp01_12_68;
	wire [WIDTH*2-1+1:0] tmp01_12_69;
	wire [WIDTH*2-1+1:0] tmp01_12_70;
	wire [WIDTH*2-1+1:0] tmp01_12_71;
	wire [WIDTH*2-1+1:0] tmp01_12_72;
	wire [WIDTH*2-1+1:0] tmp01_12_73;
	wire [WIDTH*2-1+1:0] tmp01_12_74;
	wire [WIDTH*2-1+1:0] tmp01_12_75;
	wire [WIDTH*2-1+1:0] tmp01_12_76;
	wire [WIDTH*2-1+1:0] tmp01_12_77;
	wire [WIDTH*2-1+1:0] tmp01_12_78;
	wire [WIDTH*2-1+1:0] tmp01_12_79;
	wire [WIDTH*2-1+1:0] tmp01_12_80;
	wire [WIDTH*2-1+1:0] tmp01_12_81;
	wire [WIDTH*2-1+1:0] tmp01_12_82;
	wire [WIDTH*2-1+1:0] tmp01_12_83;
	wire [WIDTH*2-1+1:0] tmp01_13_0;
	wire [WIDTH*2-1+1:0] tmp01_13_1;
	wire [WIDTH*2-1+1:0] tmp01_13_2;
	wire [WIDTH*2-1+1:0] tmp01_13_3;
	wire [WIDTH*2-1+1:0] tmp01_13_4;
	wire [WIDTH*2-1+1:0] tmp01_13_5;
	wire [WIDTH*2-1+1:0] tmp01_13_6;
	wire [WIDTH*2-1+1:0] tmp01_13_7;
	wire [WIDTH*2-1+1:0] tmp01_13_8;
	wire [WIDTH*2-1+1:0] tmp01_13_9;
	wire [WIDTH*2-1+1:0] tmp01_13_10;
	wire [WIDTH*2-1+1:0] tmp01_13_11;
	wire [WIDTH*2-1+1:0] tmp01_13_12;
	wire [WIDTH*2-1+1:0] tmp01_13_13;
	wire [WIDTH*2-1+1:0] tmp01_13_14;
	wire [WIDTH*2-1+1:0] tmp01_13_15;
	wire [WIDTH*2-1+1:0] tmp01_13_16;
	wire [WIDTH*2-1+1:0] tmp01_13_17;
	wire [WIDTH*2-1+1:0] tmp01_13_18;
	wire [WIDTH*2-1+1:0] tmp01_13_19;
	wire [WIDTH*2-1+1:0] tmp01_13_20;
	wire [WIDTH*2-1+1:0] tmp01_13_21;
	wire [WIDTH*2-1+1:0] tmp01_13_22;
	wire [WIDTH*2-1+1:0] tmp01_13_23;
	wire [WIDTH*2-1+1:0] tmp01_13_24;
	wire [WIDTH*2-1+1:0] tmp01_13_25;
	wire [WIDTH*2-1+1:0] tmp01_13_26;
	wire [WIDTH*2-1+1:0] tmp01_13_27;
	wire [WIDTH*2-1+1:0] tmp01_13_28;
	wire [WIDTH*2-1+1:0] tmp01_13_29;
	wire [WIDTH*2-1+1:0] tmp01_13_30;
	wire [WIDTH*2-1+1:0] tmp01_13_31;
	wire [WIDTH*2-1+1:0] tmp01_13_32;
	wire [WIDTH*2-1+1:0] tmp01_13_33;
	wire [WIDTH*2-1+1:0] tmp01_13_34;
	wire [WIDTH*2-1+1:0] tmp01_13_35;
	wire [WIDTH*2-1+1:0] tmp01_13_36;
	wire [WIDTH*2-1+1:0] tmp01_13_37;
	wire [WIDTH*2-1+1:0] tmp01_13_38;
	wire [WIDTH*2-1+1:0] tmp01_13_39;
	wire [WIDTH*2-1+1:0] tmp01_13_40;
	wire [WIDTH*2-1+1:0] tmp01_13_41;
	wire [WIDTH*2-1+1:0] tmp01_13_42;
	wire [WIDTH*2-1+1:0] tmp01_13_43;
	wire [WIDTH*2-1+1:0] tmp01_13_44;
	wire [WIDTH*2-1+1:0] tmp01_13_45;
	wire [WIDTH*2-1+1:0] tmp01_13_46;
	wire [WIDTH*2-1+1:0] tmp01_13_47;
	wire [WIDTH*2-1+1:0] tmp01_13_48;
	wire [WIDTH*2-1+1:0] tmp01_13_49;
	wire [WIDTH*2-1+1:0] tmp01_13_50;
	wire [WIDTH*2-1+1:0] tmp01_13_51;
	wire [WIDTH*2-1+1:0] tmp01_13_52;
	wire [WIDTH*2-1+1:0] tmp01_13_53;
	wire [WIDTH*2-1+1:0] tmp01_13_54;
	wire [WIDTH*2-1+1:0] tmp01_13_55;
	wire [WIDTH*2-1+1:0] tmp01_13_56;
	wire [WIDTH*2-1+1:0] tmp01_13_57;
	wire [WIDTH*2-1+1:0] tmp01_13_58;
	wire [WIDTH*2-1+1:0] tmp01_13_59;
	wire [WIDTH*2-1+1:0] tmp01_13_60;
	wire [WIDTH*2-1+1:0] tmp01_13_61;
	wire [WIDTH*2-1+1:0] tmp01_13_62;
	wire [WIDTH*2-1+1:0] tmp01_13_63;
	wire [WIDTH*2-1+1:0] tmp01_13_64;
	wire [WIDTH*2-1+1:0] tmp01_13_65;
	wire [WIDTH*2-1+1:0] tmp01_13_66;
	wire [WIDTH*2-1+1:0] tmp01_13_67;
	wire [WIDTH*2-1+1:0] tmp01_13_68;
	wire [WIDTH*2-1+1:0] tmp01_13_69;
	wire [WIDTH*2-1+1:0] tmp01_13_70;
	wire [WIDTH*2-1+1:0] tmp01_13_71;
	wire [WIDTH*2-1+1:0] tmp01_13_72;
	wire [WIDTH*2-1+1:0] tmp01_13_73;
	wire [WIDTH*2-1+1:0] tmp01_13_74;
	wire [WIDTH*2-1+1:0] tmp01_13_75;
	wire [WIDTH*2-1+1:0] tmp01_13_76;
	wire [WIDTH*2-1+1:0] tmp01_13_77;
	wire [WIDTH*2-1+1:0] tmp01_13_78;
	wire [WIDTH*2-1+1:0] tmp01_13_79;
	wire [WIDTH*2-1+1:0] tmp01_13_80;
	wire [WIDTH*2-1+1:0] tmp01_13_81;
	wire [WIDTH*2-1+1:0] tmp01_13_82;
	wire [WIDTH*2-1+1:0] tmp01_13_83;
	wire [WIDTH*2-1+1:0] tmp01_14_0;
	wire [WIDTH*2-1+1:0] tmp01_14_1;
	wire [WIDTH*2-1+1:0] tmp01_14_2;
	wire [WIDTH*2-1+1:0] tmp01_14_3;
	wire [WIDTH*2-1+1:0] tmp01_14_4;
	wire [WIDTH*2-1+1:0] tmp01_14_5;
	wire [WIDTH*2-1+1:0] tmp01_14_6;
	wire [WIDTH*2-1+1:0] tmp01_14_7;
	wire [WIDTH*2-1+1:0] tmp01_14_8;
	wire [WIDTH*2-1+1:0] tmp01_14_9;
	wire [WIDTH*2-1+1:0] tmp01_14_10;
	wire [WIDTH*2-1+1:0] tmp01_14_11;
	wire [WIDTH*2-1+1:0] tmp01_14_12;
	wire [WIDTH*2-1+1:0] tmp01_14_13;
	wire [WIDTH*2-1+1:0] tmp01_14_14;
	wire [WIDTH*2-1+1:0] tmp01_14_15;
	wire [WIDTH*2-1+1:0] tmp01_14_16;
	wire [WIDTH*2-1+1:0] tmp01_14_17;
	wire [WIDTH*2-1+1:0] tmp01_14_18;
	wire [WIDTH*2-1+1:0] tmp01_14_19;
	wire [WIDTH*2-1+1:0] tmp01_14_20;
	wire [WIDTH*2-1+1:0] tmp01_14_21;
	wire [WIDTH*2-1+1:0] tmp01_14_22;
	wire [WIDTH*2-1+1:0] tmp01_14_23;
	wire [WIDTH*2-1+1:0] tmp01_14_24;
	wire [WIDTH*2-1+1:0] tmp01_14_25;
	wire [WIDTH*2-1+1:0] tmp01_14_26;
	wire [WIDTH*2-1+1:0] tmp01_14_27;
	wire [WIDTH*2-1+1:0] tmp01_14_28;
	wire [WIDTH*2-1+1:0] tmp01_14_29;
	wire [WIDTH*2-1+1:0] tmp01_14_30;
	wire [WIDTH*2-1+1:0] tmp01_14_31;
	wire [WIDTH*2-1+1:0] tmp01_14_32;
	wire [WIDTH*2-1+1:0] tmp01_14_33;
	wire [WIDTH*2-1+1:0] tmp01_14_34;
	wire [WIDTH*2-1+1:0] tmp01_14_35;
	wire [WIDTH*2-1+1:0] tmp01_14_36;
	wire [WIDTH*2-1+1:0] tmp01_14_37;
	wire [WIDTH*2-1+1:0] tmp01_14_38;
	wire [WIDTH*2-1+1:0] tmp01_14_39;
	wire [WIDTH*2-1+1:0] tmp01_14_40;
	wire [WIDTH*2-1+1:0] tmp01_14_41;
	wire [WIDTH*2-1+1:0] tmp01_14_42;
	wire [WIDTH*2-1+1:0] tmp01_14_43;
	wire [WIDTH*2-1+1:0] tmp01_14_44;
	wire [WIDTH*2-1+1:0] tmp01_14_45;
	wire [WIDTH*2-1+1:0] tmp01_14_46;
	wire [WIDTH*2-1+1:0] tmp01_14_47;
	wire [WIDTH*2-1+1:0] tmp01_14_48;
	wire [WIDTH*2-1+1:0] tmp01_14_49;
	wire [WIDTH*2-1+1:0] tmp01_14_50;
	wire [WIDTH*2-1+1:0] tmp01_14_51;
	wire [WIDTH*2-1+1:0] tmp01_14_52;
	wire [WIDTH*2-1+1:0] tmp01_14_53;
	wire [WIDTH*2-1+1:0] tmp01_14_54;
	wire [WIDTH*2-1+1:0] tmp01_14_55;
	wire [WIDTH*2-1+1:0] tmp01_14_56;
	wire [WIDTH*2-1+1:0] tmp01_14_57;
	wire [WIDTH*2-1+1:0] tmp01_14_58;
	wire [WIDTH*2-1+1:0] tmp01_14_59;
	wire [WIDTH*2-1+1:0] tmp01_14_60;
	wire [WIDTH*2-1+1:0] tmp01_14_61;
	wire [WIDTH*2-1+1:0] tmp01_14_62;
	wire [WIDTH*2-1+1:0] tmp01_14_63;
	wire [WIDTH*2-1+1:0] tmp01_14_64;
	wire [WIDTH*2-1+1:0] tmp01_14_65;
	wire [WIDTH*2-1+1:0] tmp01_14_66;
	wire [WIDTH*2-1+1:0] tmp01_14_67;
	wire [WIDTH*2-1+1:0] tmp01_14_68;
	wire [WIDTH*2-1+1:0] tmp01_14_69;
	wire [WIDTH*2-1+1:0] tmp01_14_70;
	wire [WIDTH*2-1+1:0] tmp01_14_71;
	wire [WIDTH*2-1+1:0] tmp01_14_72;
	wire [WIDTH*2-1+1:0] tmp01_14_73;
	wire [WIDTH*2-1+1:0] tmp01_14_74;
	wire [WIDTH*2-1+1:0] tmp01_14_75;
	wire [WIDTH*2-1+1:0] tmp01_14_76;
	wire [WIDTH*2-1+1:0] tmp01_14_77;
	wire [WIDTH*2-1+1:0] tmp01_14_78;
	wire [WIDTH*2-1+1:0] tmp01_14_79;
	wire [WIDTH*2-1+1:0] tmp01_14_80;
	wire [WIDTH*2-1+1:0] tmp01_14_81;
	wire [WIDTH*2-1+1:0] tmp01_14_82;
	wire [WIDTH*2-1+1:0] tmp01_14_83;
	wire [WIDTH*2-1+1:0] tmp01_15_0;
	wire [WIDTH*2-1+1:0] tmp01_15_1;
	wire [WIDTH*2-1+1:0] tmp01_15_2;
	wire [WIDTH*2-1+1:0] tmp01_15_3;
	wire [WIDTH*2-1+1:0] tmp01_15_4;
	wire [WIDTH*2-1+1:0] tmp01_15_5;
	wire [WIDTH*2-1+1:0] tmp01_15_6;
	wire [WIDTH*2-1+1:0] tmp01_15_7;
	wire [WIDTH*2-1+1:0] tmp01_15_8;
	wire [WIDTH*2-1+1:0] tmp01_15_9;
	wire [WIDTH*2-1+1:0] tmp01_15_10;
	wire [WIDTH*2-1+1:0] tmp01_15_11;
	wire [WIDTH*2-1+1:0] tmp01_15_12;
	wire [WIDTH*2-1+1:0] tmp01_15_13;
	wire [WIDTH*2-1+1:0] tmp01_15_14;
	wire [WIDTH*2-1+1:0] tmp01_15_15;
	wire [WIDTH*2-1+1:0] tmp01_15_16;
	wire [WIDTH*2-1+1:0] tmp01_15_17;
	wire [WIDTH*2-1+1:0] tmp01_15_18;
	wire [WIDTH*2-1+1:0] tmp01_15_19;
	wire [WIDTH*2-1+1:0] tmp01_15_20;
	wire [WIDTH*2-1+1:0] tmp01_15_21;
	wire [WIDTH*2-1+1:0] tmp01_15_22;
	wire [WIDTH*2-1+1:0] tmp01_15_23;
	wire [WIDTH*2-1+1:0] tmp01_15_24;
	wire [WIDTH*2-1+1:0] tmp01_15_25;
	wire [WIDTH*2-1+1:0] tmp01_15_26;
	wire [WIDTH*2-1+1:0] tmp01_15_27;
	wire [WIDTH*2-1+1:0] tmp01_15_28;
	wire [WIDTH*2-1+1:0] tmp01_15_29;
	wire [WIDTH*2-1+1:0] tmp01_15_30;
	wire [WIDTH*2-1+1:0] tmp01_15_31;
	wire [WIDTH*2-1+1:0] tmp01_15_32;
	wire [WIDTH*2-1+1:0] tmp01_15_33;
	wire [WIDTH*2-1+1:0] tmp01_15_34;
	wire [WIDTH*2-1+1:0] tmp01_15_35;
	wire [WIDTH*2-1+1:0] tmp01_15_36;
	wire [WIDTH*2-1+1:0] tmp01_15_37;
	wire [WIDTH*2-1+1:0] tmp01_15_38;
	wire [WIDTH*2-1+1:0] tmp01_15_39;
	wire [WIDTH*2-1+1:0] tmp01_15_40;
	wire [WIDTH*2-1+1:0] tmp01_15_41;
	wire [WIDTH*2-1+1:0] tmp01_15_42;
	wire [WIDTH*2-1+1:0] tmp01_15_43;
	wire [WIDTH*2-1+1:0] tmp01_15_44;
	wire [WIDTH*2-1+1:0] tmp01_15_45;
	wire [WIDTH*2-1+1:0] tmp01_15_46;
	wire [WIDTH*2-1+1:0] tmp01_15_47;
	wire [WIDTH*2-1+1:0] tmp01_15_48;
	wire [WIDTH*2-1+1:0] tmp01_15_49;
	wire [WIDTH*2-1+1:0] tmp01_15_50;
	wire [WIDTH*2-1+1:0] tmp01_15_51;
	wire [WIDTH*2-1+1:0] tmp01_15_52;
	wire [WIDTH*2-1+1:0] tmp01_15_53;
	wire [WIDTH*2-1+1:0] tmp01_15_54;
	wire [WIDTH*2-1+1:0] tmp01_15_55;
	wire [WIDTH*2-1+1:0] tmp01_15_56;
	wire [WIDTH*2-1+1:0] tmp01_15_57;
	wire [WIDTH*2-1+1:0] tmp01_15_58;
	wire [WIDTH*2-1+1:0] tmp01_15_59;
	wire [WIDTH*2-1+1:0] tmp01_15_60;
	wire [WIDTH*2-1+1:0] tmp01_15_61;
	wire [WIDTH*2-1+1:0] tmp01_15_62;
	wire [WIDTH*2-1+1:0] tmp01_15_63;
	wire [WIDTH*2-1+1:0] tmp01_15_64;
	wire [WIDTH*2-1+1:0] tmp01_15_65;
	wire [WIDTH*2-1+1:0] tmp01_15_66;
	wire [WIDTH*2-1+1:0] tmp01_15_67;
	wire [WIDTH*2-1+1:0] tmp01_15_68;
	wire [WIDTH*2-1+1:0] tmp01_15_69;
	wire [WIDTH*2-1+1:0] tmp01_15_70;
	wire [WIDTH*2-1+1:0] tmp01_15_71;
	wire [WIDTH*2-1+1:0] tmp01_15_72;
	wire [WIDTH*2-1+1:0] tmp01_15_73;
	wire [WIDTH*2-1+1:0] tmp01_15_74;
	wire [WIDTH*2-1+1:0] tmp01_15_75;
	wire [WIDTH*2-1+1:0] tmp01_15_76;
	wire [WIDTH*2-1+1:0] tmp01_15_77;
	wire [WIDTH*2-1+1:0] tmp01_15_78;
	wire [WIDTH*2-1+1:0] tmp01_15_79;
	wire [WIDTH*2-1+1:0] tmp01_15_80;
	wire [WIDTH*2-1+1:0] tmp01_15_81;
	wire [WIDTH*2-1+1:0] tmp01_15_82;
	wire [WIDTH*2-1+1:0] tmp01_15_83;
	wire [WIDTH*2-1+1:0] tmp01_16_0;
	wire [WIDTH*2-1+1:0] tmp01_16_1;
	wire [WIDTH*2-1+1:0] tmp01_16_2;
	wire [WIDTH*2-1+1:0] tmp01_16_3;
	wire [WIDTH*2-1+1:0] tmp01_16_4;
	wire [WIDTH*2-1+1:0] tmp01_16_5;
	wire [WIDTH*2-1+1:0] tmp01_16_6;
	wire [WIDTH*2-1+1:0] tmp01_16_7;
	wire [WIDTH*2-1+1:0] tmp01_16_8;
	wire [WIDTH*2-1+1:0] tmp01_16_9;
	wire [WIDTH*2-1+1:0] tmp01_16_10;
	wire [WIDTH*2-1+1:0] tmp01_16_11;
	wire [WIDTH*2-1+1:0] tmp01_16_12;
	wire [WIDTH*2-1+1:0] tmp01_16_13;
	wire [WIDTH*2-1+1:0] tmp01_16_14;
	wire [WIDTH*2-1+1:0] tmp01_16_15;
	wire [WIDTH*2-1+1:0] tmp01_16_16;
	wire [WIDTH*2-1+1:0] tmp01_16_17;
	wire [WIDTH*2-1+1:0] tmp01_16_18;
	wire [WIDTH*2-1+1:0] tmp01_16_19;
	wire [WIDTH*2-1+1:0] tmp01_16_20;
	wire [WIDTH*2-1+1:0] tmp01_16_21;
	wire [WIDTH*2-1+1:0] tmp01_16_22;
	wire [WIDTH*2-1+1:0] tmp01_16_23;
	wire [WIDTH*2-1+1:0] tmp01_16_24;
	wire [WIDTH*2-1+1:0] tmp01_16_25;
	wire [WIDTH*2-1+1:0] tmp01_16_26;
	wire [WIDTH*2-1+1:0] tmp01_16_27;
	wire [WIDTH*2-1+1:0] tmp01_16_28;
	wire [WIDTH*2-1+1:0] tmp01_16_29;
	wire [WIDTH*2-1+1:0] tmp01_16_30;
	wire [WIDTH*2-1+1:0] tmp01_16_31;
	wire [WIDTH*2-1+1:0] tmp01_16_32;
	wire [WIDTH*2-1+1:0] tmp01_16_33;
	wire [WIDTH*2-1+1:0] tmp01_16_34;
	wire [WIDTH*2-1+1:0] tmp01_16_35;
	wire [WIDTH*2-1+1:0] tmp01_16_36;
	wire [WIDTH*2-1+1:0] tmp01_16_37;
	wire [WIDTH*2-1+1:0] tmp01_16_38;
	wire [WIDTH*2-1+1:0] tmp01_16_39;
	wire [WIDTH*2-1+1:0] tmp01_16_40;
	wire [WIDTH*2-1+1:0] tmp01_16_41;
	wire [WIDTH*2-1+1:0] tmp01_16_42;
	wire [WIDTH*2-1+1:0] tmp01_16_43;
	wire [WIDTH*2-1+1:0] tmp01_16_44;
	wire [WIDTH*2-1+1:0] tmp01_16_45;
	wire [WIDTH*2-1+1:0] tmp01_16_46;
	wire [WIDTH*2-1+1:0] tmp01_16_47;
	wire [WIDTH*2-1+1:0] tmp01_16_48;
	wire [WIDTH*2-1+1:0] tmp01_16_49;
	wire [WIDTH*2-1+1:0] tmp01_16_50;
	wire [WIDTH*2-1+1:0] tmp01_16_51;
	wire [WIDTH*2-1+1:0] tmp01_16_52;
	wire [WIDTH*2-1+1:0] tmp01_16_53;
	wire [WIDTH*2-1+1:0] tmp01_16_54;
	wire [WIDTH*2-1+1:0] tmp01_16_55;
	wire [WIDTH*2-1+1:0] tmp01_16_56;
	wire [WIDTH*2-1+1:0] tmp01_16_57;
	wire [WIDTH*2-1+1:0] tmp01_16_58;
	wire [WIDTH*2-1+1:0] tmp01_16_59;
	wire [WIDTH*2-1+1:0] tmp01_16_60;
	wire [WIDTH*2-1+1:0] tmp01_16_61;
	wire [WIDTH*2-1+1:0] tmp01_16_62;
	wire [WIDTH*2-1+1:0] tmp01_16_63;
	wire [WIDTH*2-1+1:0] tmp01_16_64;
	wire [WIDTH*2-1+1:0] tmp01_16_65;
	wire [WIDTH*2-1+1:0] tmp01_16_66;
	wire [WIDTH*2-1+1:0] tmp01_16_67;
	wire [WIDTH*2-1+1:0] tmp01_16_68;
	wire [WIDTH*2-1+1:0] tmp01_16_69;
	wire [WIDTH*2-1+1:0] tmp01_16_70;
	wire [WIDTH*2-1+1:0] tmp01_16_71;
	wire [WIDTH*2-1+1:0] tmp01_16_72;
	wire [WIDTH*2-1+1:0] tmp01_16_73;
	wire [WIDTH*2-1+1:0] tmp01_16_74;
	wire [WIDTH*2-1+1:0] tmp01_16_75;
	wire [WIDTH*2-1+1:0] tmp01_16_76;
	wire [WIDTH*2-1+1:0] tmp01_16_77;
	wire [WIDTH*2-1+1:0] tmp01_16_78;
	wire [WIDTH*2-1+1:0] tmp01_16_79;
	wire [WIDTH*2-1+1:0] tmp01_16_80;
	wire [WIDTH*2-1+1:0] tmp01_16_81;
	wire [WIDTH*2-1+1:0] tmp01_16_82;
	wire [WIDTH*2-1+1:0] tmp01_16_83;
	wire [WIDTH*2-1+1:0] tmp01_17_0;
	wire [WIDTH*2-1+1:0] tmp01_17_1;
	wire [WIDTH*2-1+1:0] tmp01_17_2;
	wire [WIDTH*2-1+1:0] tmp01_17_3;
	wire [WIDTH*2-1+1:0] tmp01_17_4;
	wire [WIDTH*2-1+1:0] tmp01_17_5;
	wire [WIDTH*2-1+1:0] tmp01_17_6;
	wire [WIDTH*2-1+1:0] tmp01_17_7;
	wire [WIDTH*2-1+1:0] tmp01_17_8;
	wire [WIDTH*2-1+1:0] tmp01_17_9;
	wire [WIDTH*2-1+1:0] tmp01_17_10;
	wire [WIDTH*2-1+1:0] tmp01_17_11;
	wire [WIDTH*2-1+1:0] tmp01_17_12;
	wire [WIDTH*2-1+1:0] tmp01_17_13;
	wire [WIDTH*2-1+1:0] tmp01_17_14;
	wire [WIDTH*2-1+1:0] tmp01_17_15;
	wire [WIDTH*2-1+1:0] tmp01_17_16;
	wire [WIDTH*2-1+1:0] tmp01_17_17;
	wire [WIDTH*2-1+1:0] tmp01_17_18;
	wire [WIDTH*2-1+1:0] tmp01_17_19;
	wire [WIDTH*2-1+1:0] tmp01_17_20;
	wire [WIDTH*2-1+1:0] tmp01_17_21;
	wire [WIDTH*2-1+1:0] tmp01_17_22;
	wire [WIDTH*2-1+1:0] tmp01_17_23;
	wire [WIDTH*2-1+1:0] tmp01_17_24;
	wire [WIDTH*2-1+1:0] tmp01_17_25;
	wire [WIDTH*2-1+1:0] tmp01_17_26;
	wire [WIDTH*2-1+1:0] tmp01_17_27;
	wire [WIDTH*2-1+1:0] tmp01_17_28;
	wire [WIDTH*2-1+1:0] tmp01_17_29;
	wire [WIDTH*2-1+1:0] tmp01_17_30;
	wire [WIDTH*2-1+1:0] tmp01_17_31;
	wire [WIDTH*2-1+1:0] tmp01_17_32;
	wire [WIDTH*2-1+1:0] tmp01_17_33;
	wire [WIDTH*2-1+1:0] tmp01_17_34;
	wire [WIDTH*2-1+1:0] tmp01_17_35;
	wire [WIDTH*2-1+1:0] tmp01_17_36;
	wire [WIDTH*2-1+1:0] tmp01_17_37;
	wire [WIDTH*2-1+1:0] tmp01_17_38;
	wire [WIDTH*2-1+1:0] tmp01_17_39;
	wire [WIDTH*2-1+1:0] tmp01_17_40;
	wire [WIDTH*2-1+1:0] tmp01_17_41;
	wire [WIDTH*2-1+1:0] tmp01_17_42;
	wire [WIDTH*2-1+1:0] tmp01_17_43;
	wire [WIDTH*2-1+1:0] tmp01_17_44;
	wire [WIDTH*2-1+1:0] tmp01_17_45;
	wire [WIDTH*2-1+1:0] tmp01_17_46;
	wire [WIDTH*2-1+1:0] tmp01_17_47;
	wire [WIDTH*2-1+1:0] tmp01_17_48;
	wire [WIDTH*2-1+1:0] tmp01_17_49;
	wire [WIDTH*2-1+1:0] tmp01_17_50;
	wire [WIDTH*2-1+1:0] tmp01_17_51;
	wire [WIDTH*2-1+1:0] tmp01_17_52;
	wire [WIDTH*2-1+1:0] tmp01_17_53;
	wire [WIDTH*2-1+1:0] tmp01_17_54;
	wire [WIDTH*2-1+1:0] tmp01_17_55;
	wire [WIDTH*2-1+1:0] tmp01_17_56;
	wire [WIDTH*2-1+1:0] tmp01_17_57;
	wire [WIDTH*2-1+1:0] tmp01_17_58;
	wire [WIDTH*2-1+1:0] tmp01_17_59;
	wire [WIDTH*2-1+1:0] tmp01_17_60;
	wire [WIDTH*2-1+1:0] tmp01_17_61;
	wire [WIDTH*2-1+1:0] tmp01_17_62;
	wire [WIDTH*2-1+1:0] tmp01_17_63;
	wire [WIDTH*2-1+1:0] tmp01_17_64;
	wire [WIDTH*2-1+1:0] tmp01_17_65;
	wire [WIDTH*2-1+1:0] tmp01_17_66;
	wire [WIDTH*2-1+1:0] tmp01_17_67;
	wire [WIDTH*2-1+1:0] tmp01_17_68;
	wire [WIDTH*2-1+1:0] tmp01_17_69;
	wire [WIDTH*2-1+1:0] tmp01_17_70;
	wire [WIDTH*2-1+1:0] tmp01_17_71;
	wire [WIDTH*2-1+1:0] tmp01_17_72;
	wire [WIDTH*2-1+1:0] tmp01_17_73;
	wire [WIDTH*2-1+1:0] tmp01_17_74;
	wire [WIDTH*2-1+1:0] tmp01_17_75;
	wire [WIDTH*2-1+1:0] tmp01_17_76;
	wire [WIDTH*2-1+1:0] tmp01_17_77;
	wire [WIDTH*2-1+1:0] tmp01_17_78;
	wire [WIDTH*2-1+1:0] tmp01_17_79;
	wire [WIDTH*2-1+1:0] tmp01_17_80;
	wire [WIDTH*2-1+1:0] tmp01_17_81;
	wire [WIDTH*2-1+1:0] tmp01_17_82;
	wire [WIDTH*2-1+1:0] tmp01_17_83;
	wire [WIDTH*2-1+1:0] tmp01_18_0;
	wire [WIDTH*2-1+1:0] tmp01_18_1;
	wire [WIDTH*2-1+1:0] tmp01_18_2;
	wire [WIDTH*2-1+1:0] tmp01_18_3;
	wire [WIDTH*2-1+1:0] tmp01_18_4;
	wire [WIDTH*2-1+1:0] tmp01_18_5;
	wire [WIDTH*2-1+1:0] tmp01_18_6;
	wire [WIDTH*2-1+1:0] tmp01_18_7;
	wire [WIDTH*2-1+1:0] tmp01_18_8;
	wire [WIDTH*2-1+1:0] tmp01_18_9;
	wire [WIDTH*2-1+1:0] tmp01_18_10;
	wire [WIDTH*2-1+1:0] tmp01_18_11;
	wire [WIDTH*2-1+1:0] tmp01_18_12;
	wire [WIDTH*2-1+1:0] tmp01_18_13;
	wire [WIDTH*2-1+1:0] tmp01_18_14;
	wire [WIDTH*2-1+1:0] tmp01_18_15;
	wire [WIDTH*2-1+1:0] tmp01_18_16;
	wire [WIDTH*2-1+1:0] tmp01_18_17;
	wire [WIDTH*2-1+1:0] tmp01_18_18;
	wire [WIDTH*2-1+1:0] tmp01_18_19;
	wire [WIDTH*2-1+1:0] tmp01_18_20;
	wire [WIDTH*2-1+1:0] tmp01_18_21;
	wire [WIDTH*2-1+1:0] tmp01_18_22;
	wire [WIDTH*2-1+1:0] tmp01_18_23;
	wire [WIDTH*2-1+1:0] tmp01_18_24;
	wire [WIDTH*2-1+1:0] tmp01_18_25;
	wire [WIDTH*2-1+1:0] tmp01_18_26;
	wire [WIDTH*2-1+1:0] tmp01_18_27;
	wire [WIDTH*2-1+1:0] tmp01_18_28;
	wire [WIDTH*2-1+1:0] tmp01_18_29;
	wire [WIDTH*2-1+1:0] tmp01_18_30;
	wire [WIDTH*2-1+1:0] tmp01_18_31;
	wire [WIDTH*2-1+1:0] tmp01_18_32;
	wire [WIDTH*2-1+1:0] tmp01_18_33;
	wire [WIDTH*2-1+1:0] tmp01_18_34;
	wire [WIDTH*2-1+1:0] tmp01_18_35;
	wire [WIDTH*2-1+1:0] tmp01_18_36;
	wire [WIDTH*2-1+1:0] tmp01_18_37;
	wire [WIDTH*2-1+1:0] tmp01_18_38;
	wire [WIDTH*2-1+1:0] tmp01_18_39;
	wire [WIDTH*2-1+1:0] tmp01_18_40;
	wire [WIDTH*2-1+1:0] tmp01_18_41;
	wire [WIDTH*2-1+1:0] tmp01_18_42;
	wire [WIDTH*2-1+1:0] tmp01_18_43;
	wire [WIDTH*2-1+1:0] tmp01_18_44;
	wire [WIDTH*2-1+1:0] tmp01_18_45;
	wire [WIDTH*2-1+1:0] tmp01_18_46;
	wire [WIDTH*2-1+1:0] tmp01_18_47;
	wire [WIDTH*2-1+1:0] tmp01_18_48;
	wire [WIDTH*2-1+1:0] tmp01_18_49;
	wire [WIDTH*2-1+1:0] tmp01_18_50;
	wire [WIDTH*2-1+1:0] tmp01_18_51;
	wire [WIDTH*2-1+1:0] tmp01_18_52;
	wire [WIDTH*2-1+1:0] tmp01_18_53;
	wire [WIDTH*2-1+1:0] tmp01_18_54;
	wire [WIDTH*2-1+1:0] tmp01_18_55;
	wire [WIDTH*2-1+1:0] tmp01_18_56;
	wire [WIDTH*2-1+1:0] tmp01_18_57;
	wire [WIDTH*2-1+1:0] tmp01_18_58;
	wire [WIDTH*2-1+1:0] tmp01_18_59;
	wire [WIDTH*2-1+1:0] tmp01_18_60;
	wire [WIDTH*2-1+1:0] tmp01_18_61;
	wire [WIDTH*2-1+1:0] tmp01_18_62;
	wire [WIDTH*2-1+1:0] tmp01_18_63;
	wire [WIDTH*2-1+1:0] tmp01_18_64;
	wire [WIDTH*2-1+1:0] tmp01_18_65;
	wire [WIDTH*2-1+1:0] tmp01_18_66;
	wire [WIDTH*2-1+1:0] tmp01_18_67;
	wire [WIDTH*2-1+1:0] tmp01_18_68;
	wire [WIDTH*2-1+1:0] tmp01_18_69;
	wire [WIDTH*2-1+1:0] tmp01_18_70;
	wire [WIDTH*2-1+1:0] tmp01_18_71;
	wire [WIDTH*2-1+1:0] tmp01_18_72;
	wire [WIDTH*2-1+1:0] tmp01_18_73;
	wire [WIDTH*2-1+1:0] tmp01_18_74;
	wire [WIDTH*2-1+1:0] tmp01_18_75;
	wire [WIDTH*2-1+1:0] tmp01_18_76;
	wire [WIDTH*2-1+1:0] tmp01_18_77;
	wire [WIDTH*2-1+1:0] tmp01_18_78;
	wire [WIDTH*2-1+1:0] tmp01_18_79;
	wire [WIDTH*2-1+1:0] tmp01_18_80;
	wire [WIDTH*2-1+1:0] tmp01_18_81;
	wire [WIDTH*2-1+1:0] tmp01_18_82;
	wire [WIDTH*2-1+1:0] tmp01_18_83;
	wire [WIDTH*2-1+1:0] tmp01_19_0;
	wire [WIDTH*2-1+1:0] tmp01_19_1;
	wire [WIDTH*2-1+1:0] tmp01_19_2;
	wire [WIDTH*2-1+1:0] tmp01_19_3;
	wire [WIDTH*2-1+1:0] tmp01_19_4;
	wire [WIDTH*2-1+1:0] tmp01_19_5;
	wire [WIDTH*2-1+1:0] tmp01_19_6;
	wire [WIDTH*2-1+1:0] tmp01_19_7;
	wire [WIDTH*2-1+1:0] tmp01_19_8;
	wire [WIDTH*2-1+1:0] tmp01_19_9;
	wire [WIDTH*2-1+1:0] tmp01_19_10;
	wire [WIDTH*2-1+1:0] tmp01_19_11;
	wire [WIDTH*2-1+1:0] tmp01_19_12;
	wire [WIDTH*2-1+1:0] tmp01_19_13;
	wire [WIDTH*2-1+1:0] tmp01_19_14;
	wire [WIDTH*2-1+1:0] tmp01_19_15;
	wire [WIDTH*2-1+1:0] tmp01_19_16;
	wire [WIDTH*2-1+1:0] tmp01_19_17;
	wire [WIDTH*2-1+1:0] tmp01_19_18;
	wire [WIDTH*2-1+1:0] tmp01_19_19;
	wire [WIDTH*2-1+1:0] tmp01_19_20;
	wire [WIDTH*2-1+1:0] tmp01_19_21;
	wire [WIDTH*2-1+1:0] tmp01_19_22;
	wire [WIDTH*2-1+1:0] tmp01_19_23;
	wire [WIDTH*2-1+1:0] tmp01_19_24;
	wire [WIDTH*2-1+1:0] tmp01_19_25;
	wire [WIDTH*2-1+1:0] tmp01_19_26;
	wire [WIDTH*2-1+1:0] tmp01_19_27;
	wire [WIDTH*2-1+1:0] tmp01_19_28;
	wire [WIDTH*2-1+1:0] tmp01_19_29;
	wire [WIDTH*2-1+1:0] tmp01_19_30;
	wire [WIDTH*2-1+1:0] tmp01_19_31;
	wire [WIDTH*2-1+1:0] tmp01_19_32;
	wire [WIDTH*2-1+1:0] tmp01_19_33;
	wire [WIDTH*2-1+1:0] tmp01_19_34;
	wire [WIDTH*2-1+1:0] tmp01_19_35;
	wire [WIDTH*2-1+1:0] tmp01_19_36;
	wire [WIDTH*2-1+1:0] tmp01_19_37;
	wire [WIDTH*2-1+1:0] tmp01_19_38;
	wire [WIDTH*2-1+1:0] tmp01_19_39;
	wire [WIDTH*2-1+1:0] tmp01_19_40;
	wire [WIDTH*2-1+1:0] tmp01_19_41;
	wire [WIDTH*2-1+1:0] tmp01_19_42;
	wire [WIDTH*2-1+1:0] tmp01_19_43;
	wire [WIDTH*2-1+1:0] tmp01_19_44;
	wire [WIDTH*2-1+1:0] tmp01_19_45;
	wire [WIDTH*2-1+1:0] tmp01_19_46;
	wire [WIDTH*2-1+1:0] tmp01_19_47;
	wire [WIDTH*2-1+1:0] tmp01_19_48;
	wire [WIDTH*2-1+1:0] tmp01_19_49;
	wire [WIDTH*2-1+1:0] tmp01_19_50;
	wire [WIDTH*2-1+1:0] tmp01_19_51;
	wire [WIDTH*2-1+1:0] tmp01_19_52;
	wire [WIDTH*2-1+1:0] tmp01_19_53;
	wire [WIDTH*2-1+1:0] tmp01_19_54;
	wire [WIDTH*2-1+1:0] tmp01_19_55;
	wire [WIDTH*2-1+1:0] tmp01_19_56;
	wire [WIDTH*2-1+1:0] tmp01_19_57;
	wire [WIDTH*2-1+1:0] tmp01_19_58;
	wire [WIDTH*2-1+1:0] tmp01_19_59;
	wire [WIDTH*2-1+1:0] tmp01_19_60;
	wire [WIDTH*2-1+1:0] tmp01_19_61;
	wire [WIDTH*2-1+1:0] tmp01_19_62;
	wire [WIDTH*2-1+1:0] tmp01_19_63;
	wire [WIDTH*2-1+1:0] tmp01_19_64;
	wire [WIDTH*2-1+1:0] tmp01_19_65;
	wire [WIDTH*2-1+1:0] tmp01_19_66;
	wire [WIDTH*2-1+1:0] tmp01_19_67;
	wire [WIDTH*2-1+1:0] tmp01_19_68;
	wire [WIDTH*2-1+1:0] tmp01_19_69;
	wire [WIDTH*2-1+1:0] tmp01_19_70;
	wire [WIDTH*2-1+1:0] tmp01_19_71;
	wire [WIDTH*2-1+1:0] tmp01_19_72;
	wire [WIDTH*2-1+1:0] tmp01_19_73;
	wire [WIDTH*2-1+1:0] tmp01_19_74;
	wire [WIDTH*2-1+1:0] tmp01_19_75;
	wire [WIDTH*2-1+1:0] tmp01_19_76;
	wire [WIDTH*2-1+1:0] tmp01_19_77;
	wire [WIDTH*2-1+1:0] tmp01_19_78;
	wire [WIDTH*2-1+1:0] tmp01_19_79;
	wire [WIDTH*2-1+1:0] tmp01_19_80;
	wire [WIDTH*2-1+1:0] tmp01_19_81;
	wire [WIDTH*2-1+1:0] tmp01_19_82;
	wire [WIDTH*2-1+1:0] tmp01_19_83;
	wire [WIDTH*2-1+1:0] tmp01_20_0;
	wire [WIDTH*2-1+1:0] tmp01_20_1;
	wire [WIDTH*2-1+1:0] tmp01_20_2;
	wire [WIDTH*2-1+1:0] tmp01_20_3;
	wire [WIDTH*2-1+1:0] tmp01_20_4;
	wire [WIDTH*2-1+1:0] tmp01_20_5;
	wire [WIDTH*2-1+1:0] tmp01_20_6;
	wire [WIDTH*2-1+1:0] tmp01_20_7;
	wire [WIDTH*2-1+1:0] tmp01_20_8;
	wire [WIDTH*2-1+1:0] tmp01_20_9;
	wire [WIDTH*2-1+1:0] tmp01_20_10;
	wire [WIDTH*2-1+1:0] tmp01_20_11;
	wire [WIDTH*2-1+1:0] tmp01_20_12;
	wire [WIDTH*2-1+1:0] tmp01_20_13;
	wire [WIDTH*2-1+1:0] tmp01_20_14;
	wire [WIDTH*2-1+1:0] tmp01_20_15;
	wire [WIDTH*2-1+1:0] tmp01_20_16;
	wire [WIDTH*2-1+1:0] tmp01_20_17;
	wire [WIDTH*2-1+1:0] tmp01_20_18;
	wire [WIDTH*2-1+1:0] tmp01_20_19;
	wire [WIDTH*2-1+1:0] tmp01_20_20;
	wire [WIDTH*2-1+1:0] tmp01_20_21;
	wire [WIDTH*2-1+1:0] tmp01_20_22;
	wire [WIDTH*2-1+1:0] tmp01_20_23;
	wire [WIDTH*2-1+1:0] tmp01_20_24;
	wire [WIDTH*2-1+1:0] tmp01_20_25;
	wire [WIDTH*2-1+1:0] tmp01_20_26;
	wire [WIDTH*2-1+1:0] tmp01_20_27;
	wire [WIDTH*2-1+1:0] tmp01_20_28;
	wire [WIDTH*2-1+1:0] tmp01_20_29;
	wire [WIDTH*2-1+1:0] tmp01_20_30;
	wire [WIDTH*2-1+1:0] tmp01_20_31;
	wire [WIDTH*2-1+1:0] tmp01_20_32;
	wire [WIDTH*2-1+1:0] tmp01_20_33;
	wire [WIDTH*2-1+1:0] tmp01_20_34;
	wire [WIDTH*2-1+1:0] tmp01_20_35;
	wire [WIDTH*2-1+1:0] tmp01_20_36;
	wire [WIDTH*2-1+1:0] tmp01_20_37;
	wire [WIDTH*2-1+1:0] tmp01_20_38;
	wire [WIDTH*2-1+1:0] tmp01_20_39;
	wire [WIDTH*2-1+1:0] tmp01_20_40;
	wire [WIDTH*2-1+1:0] tmp01_20_41;
	wire [WIDTH*2-1+1:0] tmp01_20_42;
	wire [WIDTH*2-1+1:0] tmp01_20_43;
	wire [WIDTH*2-1+1:0] tmp01_20_44;
	wire [WIDTH*2-1+1:0] tmp01_20_45;
	wire [WIDTH*2-1+1:0] tmp01_20_46;
	wire [WIDTH*2-1+1:0] tmp01_20_47;
	wire [WIDTH*2-1+1:0] tmp01_20_48;
	wire [WIDTH*2-1+1:0] tmp01_20_49;
	wire [WIDTH*2-1+1:0] tmp01_20_50;
	wire [WIDTH*2-1+1:0] tmp01_20_51;
	wire [WIDTH*2-1+1:0] tmp01_20_52;
	wire [WIDTH*2-1+1:0] tmp01_20_53;
	wire [WIDTH*2-1+1:0] tmp01_20_54;
	wire [WIDTH*2-1+1:0] tmp01_20_55;
	wire [WIDTH*2-1+1:0] tmp01_20_56;
	wire [WIDTH*2-1+1:0] tmp01_20_57;
	wire [WIDTH*2-1+1:0] tmp01_20_58;
	wire [WIDTH*2-1+1:0] tmp01_20_59;
	wire [WIDTH*2-1+1:0] tmp01_20_60;
	wire [WIDTH*2-1+1:0] tmp01_20_61;
	wire [WIDTH*2-1+1:0] tmp01_20_62;
	wire [WIDTH*2-1+1:0] tmp01_20_63;
	wire [WIDTH*2-1+1:0] tmp01_20_64;
	wire [WIDTH*2-1+1:0] tmp01_20_65;
	wire [WIDTH*2-1+1:0] tmp01_20_66;
	wire [WIDTH*2-1+1:0] tmp01_20_67;
	wire [WIDTH*2-1+1:0] tmp01_20_68;
	wire [WIDTH*2-1+1:0] tmp01_20_69;
	wire [WIDTH*2-1+1:0] tmp01_20_70;
	wire [WIDTH*2-1+1:0] tmp01_20_71;
	wire [WIDTH*2-1+1:0] tmp01_20_72;
	wire [WIDTH*2-1+1:0] tmp01_20_73;
	wire [WIDTH*2-1+1:0] tmp01_20_74;
	wire [WIDTH*2-1+1:0] tmp01_20_75;
	wire [WIDTH*2-1+1:0] tmp01_20_76;
	wire [WIDTH*2-1+1:0] tmp01_20_77;
	wire [WIDTH*2-1+1:0] tmp01_20_78;
	wire [WIDTH*2-1+1:0] tmp01_20_79;
	wire [WIDTH*2-1+1:0] tmp01_20_80;
	wire [WIDTH*2-1+1:0] tmp01_20_81;
	wire [WIDTH*2-1+1:0] tmp01_20_82;
	wire [WIDTH*2-1+1:0] tmp01_20_83;
	wire [WIDTH*2-1+1:0] tmp01_21_0;
	wire [WIDTH*2-1+1:0] tmp01_21_1;
	wire [WIDTH*2-1+1:0] tmp01_21_2;
	wire [WIDTH*2-1+1:0] tmp01_21_3;
	wire [WIDTH*2-1+1:0] tmp01_21_4;
	wire [WIDTH*2-1+1:0] tmp01_21_5;
	wire [WIDTH*2-1+1:0] tmp01_21_6;
	wire [WIDTH*2-1+1:0] tmp01_21_7;
	wire [WIDTH*2-1+1:0] tmp01_21_8;
	wire [WIDTH*2-1+1:0] tmp01_21_9;
	wire [WIDTH*2-1+1:0] tmp01_21_10;
	wire [WIDTH*2-1+1:0] tmp01_21_11;
	wire [WIDTH*2-1+1:0] tmp01_21_12;
	wire [WIDTH*2-1+1:0] tmp01_21_13;
	wire [WIDTH*2-1+1:0] tmp01_21_14;
	wire [WIDTH*2-1+1:0] tmp01_21_15;
	wire [WIDTH*2-1+1:0] tmp01_21_16;
	wire [WIDTH*2-1+1:0] tmp01_21_17;
	wire [WIDTH*2-1+1:0] tmp01_21_18;
	wire [WIDTH*2-1+1:0] tmp01_21_19;
	wire [WIDTH*2-1+1:0] tmp01_21_20;
	wire [WIDTH*2-1+1:0] tmp01_21_21;
	wire [WIDTH*2-1+1:0] tmp01_21_22;
	wire [WIDTH*2-1+1:0] tmp01_21_23;
	wire [WIDTH*2-1+1:0] tmp01_21_24;
	wire [WIDTH*2-1+1:0] tmp01_21_25;
	wire [WIDTH*2-1+1:0] tmp01_21_26;
	wire [WIDTH*2-1+1:0] tmp01_21_27;
	wire [WIDTH*2-1+1:0] tmp01_21_28;
	wire [WIDTH*2-1+1:0] tmp01_21_29;
	wire [WIDTH*2-1+1:0] tmp01_21_30;
	wire [WIDTH*2-1+1:0] tmp01_21_31;
	wire [WIDTH*2-1+1:0] tmp01_21_32;
	wire [WIDTH*2-1+1:0] tmp01_21_33;
	wire [WIDTH*2-1+1:0] tmp01_21_34;
	wire [WIDTH*2-1+1:0] tmp01_21_35;
	wire [WIDTH*2-1+1:0] tmp01_21_36;
	wire [WIDTH*2-1+1:0] tmp01_21_37;
	wire [WIDTH*2-1+1:0] tmp01_21_38;
	wire [WIDTH*2-1+1:0] tmp01_21_39;
	wire [WIDTH*2-1+1:0] tmp01_21_40;
	wire [WIDTH*2-1+1:0] tmp01_21_41;
	wire [WIDTH*2-1+1:0] tmp01_21_42;
	wire [WIDTH*2-1+1:0] tmp01_21_43;
	wire [WIDTH*2-1+1:0] tmp01_21_44;
	wire [WIDTH*2-1+1:0] tmp01_21_45;
	wire [WIDTH*2-1+1:0] tmp01_21_46;
	wire [WIDTH*2-1+1:0] tmp01_21_47;
	wire [WIDTH*2-1+1:0] tmp01_21_48;
	wire [WIDTH*2-1+1:0] tmp01_21_49;
	wire [WIDTH*2-1+1:0] tmp01_21_50;
	wire [WIDTH*2-1+1:0] tmp01_21_51;
	wire [WIDTH*2-1+1:0] tmp01_21_52;
	wire [WIDTH*2-1+1:0] tmp01_21_53;
	wire [WIDTH*2-1+1:0] tmp01_21_54;
	wire [WIDTH*2-1+1:0] tmp01_21_55;
	wire [WIDTH*2-1+1:0] tmp01_21_56;
	wire [WIDTH*2-1+1:0] tmp01_21_57;
	wire [WIDTH*2-1+1:0] tmp01_21_58;
	wire [WIDTH*2-1+1:0] tmp01_21_59;
	wire [WIDTH*2-1+1:0] tmp01_21_60;
	wire [WIDTH*2-1+1:0] tmp01_21_61;
	wire [WIDTH*2-1+1:0] tmp01_21_62;
	wire [WIDTH*2-1+1:0] tmp01_21_63;
	wire [WIDTH*2-1+1:0] tmp01_21_64;
	wire [WIDTH*2-1+1:0] tmp01_21_65;
	wire [WIDTH*2-1+1:0] tmp01_21_66;
	wire [WIDTH*2-1+1:0] tmp01_21_67;
	wire [WIDTH*2-1+1:0] tmp01_21_68;
	wire [WIDTH*2-1+1:0] tmp01_21_69;
	wire [WIDTH*2-1+1:0] tmp01_21_70;
	wire [WIDTH*2-1+1:0] tmp01_21_71;
	wire [WIDTH*2-1+1:0] tmp01_21_72;
	wire [WIDTH*2-1+1:0] tmp01_21_73;
	wire [WIDTH*2-1+1:0] tmp01_21_74;
	wire [WIDTH*2-1+1:0] tmp01_21_75;
	wire [WIDTH*2-1+1:0] tmp01_21_76;
	wire [WIDTH*2-1+1:0] tmp01_21_77;
	wire [WIDTH*2-1+1:0] tmp01_21_78;
	wire [WIDTH*2-1+1:0] tmp01_21_79;
	wire [WIDTH*2-1+1:0] tmp01_21_80;
	wire [WIDTH*2-1+1:0] tmp01_21_81;
	wire [WIDTH*2-1+1:0] tmp01_21_82;
	wire [WIDTH*2-1+1:0] tmp01_21_83;
	wire [WIDTH*2-1+1:0] tmp01_22_0;
	wire [WIDTH*2-1+1:0] tmp01_22_1;
	wire [WIDTH*2-1+1:0] tmp01_22_2;
	wire [WIDTH*2-1+1:0] tmp01_22_3;
	wire [WIDTH*2-1+1:0] tmp01_22_4;
	wire [WIDTH*2-1+1:0] tmp01_22_5;
	wire [WIDTH*2-1+1:0] tmp01_22_6;
	wire [WIDTH*2-1+1:0] tmp01_22_7;
	wire [WIDTH*2-1+1:0] tmp01_22_8;
	wire [WIDTH*2-1+1:0] tmp01_22_9;
	wire [WIDTH*2-1+1:0] tmp01_22_10;
	wire [WIDTH*2-1+1:0] tmp01_22_11;
	wire [WIDTH*2-1+1:0] tmp01_22_12;
	wire [WIDTH*2-1+1:0] tmp01_22_13;
	wire [WIDTH*2-1+1:0] tmp01_22_14;
	wire [WIDTH*2-1+1:0] tmp01_22_15;
	wire [WIDTH*2-1+1:0] tmp01_22_16;
	wire [WIDTH*2-1+1:0] tmp01_22_17;
	wire [WIDTH*2-1+1:0] tmp01_22_18;
	wire [WIDTH*2-1+1:0] tmp01_22_19;
	wire [WIDTH*2-1+1:0] tmp01_22_20;
	wire [WIDTH*2-1+1:0] tmp01_22_21;
	wire [WIDTH*2-1+1:0] tmp01_22_22;
	wire [WIDTH*2-1+1:0] tmp01_22_23;
	wire [WIDTH*2-1+1:0] tmp01_22_24;
	wire [WIDTH*2-1+1:0] tmp01_22_25;
	wire [WIDTH*2-1+1:0] tmp01_22_26;
	wire [WIDTH*2-1+1:0] tmp01_22_27;
	wire [WIDTH*2-1+1:0] tmp01_22_28;
	wire [WIDTH*2-1+1:0] tmp01_22_29;
	wire [WIDTH*2-1+1:0] tmp01_22_30;
	wire [WIDTH*2-1+1:0] tmp01_22_31;
	wire [WIDTH*2-1+1:0] tmp01_22_32;
	wire [WIDTH*2-1+1:0] tmp01_22_33;
	wire [WIDTH*2-1+1:0] tmp01_22_34;
	wire [WIDTH*2-1+1:0] tmp01_22_35;
	wire [WIDTH*2-1+1:0] tmp01_22_36;
	wire [WIDTH*2-1+1:0] tmp01_22_37;
	wire [WIDTH*2-1+1:0] tmp01_22_38;
	wire [WIDTH*2-1+1:0] tmp01_22_39;
	wire [WIDTH*2-1+1:0] tmp01_22_40;
	wire [WIDTH*2-1+1:0] tmp01_22_41;
	wire [WIDTH*2-1+1:0] tmp01_22_42;
	wire [WIDTH*2-1+1:0] tmp01_22_43;
	wire [WIDTH*2-1+1:0] tmp01_22_44;
	wire [WIDTH*2-1+1:0] tmp01_22_45;
	wire [WIDTH*2-1+1:0] tmp01_22_46;
	wire [WIDTH*2-1+1:0] tmp01_22_47;
	wire [WIDTH*2-1+1:0] tmp01_22_48;
	wire [WIDTH*2-1+1:0] tmp01_22_49;
	wire [WIDTH*2-1+1:0] tmp01_22_50;
	wire [WIDTH*2-1+1:0] tmp01_22_51;
	wire [WIDTH*2-1+1:0] tmp01_22_52;
	wire [WIDTH*2-1+1:0] tmp01_22_53;
	wire [WIDTH*2-1+1:0] tmp01_22_54;
	wire [WIDTH*2-1+1:0] tmp01_22_55;
	wire [WIDTH*2-1+1:0] tmp01_22_56;
	wire [WIDTH*2-1+1:0] tmp01_22_57;
	wire [WIDTH*2-1+1:0] tmp01_22_58;
	wire [WIDTH*2-1+1:0] tmp01_22_59;
	wire [WIDTH*2-1+1:0] tmp01_22_60;
	wire [WIDTH*2-1+1:0] tmp01_22_61;
	wire [WIDTH*2-1+1:0] tmp01_22_62;
	wire [WIDTH*2-1+1:0] tmp01_22_63;
	wire [WIDTH*2-1+1:0] tmp01_22_64;
	wire [WIDTH*2-1+1:0] tmp01_22_65;
	wire [WIDTH*2-1+1:0] tmp01_22_66;
	wire [WIDTH*2-1+1:0] tmp01_22_67;
	wire [WIDTH*2-1+1:0] tmp01_22_68;
	wire [WIDTH*2-1+1:0] tmp01_22_69;
	wire [WIDTH*2-1+1:0] tmp01_22_70;
	wire [WIDTH*2-1+1:0] tmp01_22_71;
	wire [WIDTH*2-1+1:0] tmp01_22_72;
	wire [WIDTH*2-1+1:0] tmp01_22_73;
	wire [WIDTH*2-1+1:0] tmp01_22_74;
	wire [WIDTH*2-1+1:0] tmp01_22_75;
	wire [WIDTH*2-1+1:0] tmp01_22_76;
	wire [WIDTH*2-1+1:0] tmp01_22_77;
	wire [WIDTH*2-1+1:0] tmp01_22_78;
	wire [WIDTH*2-1+1:0] tmp01_22_79;
	wire [WIDTH*2-1+1:0] tmp01_22_80;
	wire [WIDTH*2-1+1:0] tmp01_22_81;
	wire [WIDTH*2-1+1:0] tmp01_22_82;
	wire [WIDTH*2-1+1:0] tmp01_22_83;
	wire [WIDTH*2-1+1:0] tmp01_23_0;
	wire [WIDTH*2-1+1:0] tmp01_23_1;
	wire [WIDTH*2-1+1:0] tmp01_23_2;
	wire [WIDTH*2-1+1:0] tmp01_23_3;
	wire [WIDTH*2-1+1:0] tmp01_23_4;
	wire [WIDTH*2-1+1:0] tmp01_23_5;
	wire [WIDTH*2-1+1:0] tmp01_23_6;
	wire [WIDTH*2-1+1:0] tmp01_23_7;
	wire [WIDTH*2-1+1:0] tmp01_23_8;
	wire [WIDTH*2-1+1:0] tmp01_23_9;
	wire [WIDTH*2-1+1:0] tmp01_23_10;
	wire [WIDTH*2-1+1:0] tmp01_23_11;
	wire [WIDTH*2-1+1:0] tmp01_23_12;
	wire [WIDTH*2-1+1:0] tmp01_23_13;
	wire [WIDTH*2-1+1:0] tmp01_23_14;
	wire [WIDTH*2-1+1:0] tmp01_23_15;
	wire [WIDTH*2-1+1:0] tmp01_23_16;
	wire [WIDTH*2-1+1:0] tmp01_23_17;
	wire [WIDTH*2-1+1:0] tmp01_23_18;
	wire [WIDTH*2-1+1:0] tmp01_23_19;
	wire [WIDTH*2-1+1:0] tmp01_23_20;
	wire [WIDTH*2-1+1:0] tmp01_23_21;
	wire [WIDTH*2-1+1:0] tmp01_23_22;
	wire [WIDTH*2-1+1:0] tmp01_23_23;
	wire [WIDTH*2-1+1:0] tmp01_23_24;
	wire [WIDTH*2-1+1:0] tmp01_23_25;
	wire [WIDTH*2-1+1:0] tmp01_23_26;
	wire [WIDTH*2-1+1:0] tmp01_23_27;
	wire [WIDTH*2-1+1:0] tmp01_23_28;
	wire [WIDTH*2-1+1:0] tmp01_23_29;
	wire [WIDTH*2-1+1:0] tmp01_23_30;
	wire [WIDTH*2-1+1:0] tmp01_23_31;
	wire [WIDTH*2-1+1:0] tmp01_23_32;
	wire [WIDTH*2-1+1:0] tmp01_23_33;
	wire [WIDTH*2-1+1:0] tmp01_23_34;
	wire [WIDTH*2-1+1:0] tmp01_23_35;
	wire [WIDTH*2-1+1:0] tmp01_23_36;
	wire [WIDTH*2-1+1:0] tmp01_23_37;
	wire [WIDTH*2-1+1:0] tmp01_23_38;
	wire [WIDTH*2-1+1:0] tmp01_23_39;
	wire [WIDTH*2-1+1:0] tmp01_23_40;
	wire [WIDTH*2-1+1:0] tmp01_23_41;
	wire [WIDTH*2-1+1:0] tmp01_23_42;
	wire [WIDTH*2-1+1:0] tmp01_23_43;
	wire [WIDTH*2-1+1:0] tmp01_23_44;
	wire [WIDTH*2-1+1:0] tmp01_23_45;
	wire [WIDTH*2-1+1:0] tmp01_23_46;
	wire [WIDTH*2-1+1:0] tmp01_23_47;
	wire [WIDTH*2-1+1:0] tmp01_23_48;
	wire [WIDTH*2-1+1:0] tmp01_23_49;
	wire [WIDTH*2-1+1:0] tmp01_23_50;
	wire [WIDTH*2-1+1:0] tmp01_23_51;
	wire [WIDTH*2-1+1:0] tmp01_23_52;
	wire [WIDTH*2-1+1:0] tmp01_23_53;
	wire [WIDTH*2-1+1:0] tmp01_23_54;
	wire [WIDTH*2-1+1:0] tmp01_23_55;
	wire [WIDTH*2-1+1:0] tmp01_23_56;
	wire [WIDTH*2-1+1:0] tmp01_23_57;
	wire [WIDTH*2-1+1:0] tmp01_23_58;
	wire [WIDTH*2-1+1:0] tmp01_23_59;
	wire [WIDTH*2-1+1:0] tmp01_23_60;
	wire [WIDTH*2-1+1:0] tmp01_23_61;
	wire [WIDTH*2-1+1:0] tmp01_23_62;
	wire [WIDTH*2-1+1:0] tmp01_23_63;
	wire [WIDTH*2-1+1:0] tmp01_23_64;
	wire [WIDTH*2-1+1:0] tmp01_23_65;
	wire [WIDTH*2-1+1:0] tmp01_23_66;
	wire [WIDTH*2-1+1:0] tmp01_23_67;
	wire [WIDTH*2-1+1:0] tmp01_23_68;
	wire [WIDTH*2-1+1:0] tmp01_23_69;
	wire [WIDTH*2-1+1:0] tmp01_23_70;
	wire [WIDTH*2-1+1:0] tmp01_23_71;
	wire [WIDTH*2-1+1:0] tmp01_23_72;
	wire [WIDTH*2-1+1:0] tmp01_23_73;
	wire [WIDTH*2-1+1:0] tmp01_23_74;
	wire [WIDTH*2-1+1:0] tmp01_23_75;
	wire [WIDTH*2-1+1:0] tmp01_23_76;
	wire [WIDTH*2-1+1:0] tmp01_23_77;
	wire [WIDTH*2-1+1:0] tmp01_23_78;
	wire [WIDTH*2-1+1:0] tmp01_23_79;
	wire [WIDTH*2-1+1:0] tmp01_23_80;
	wire [WIDTH*2-1+1:0] tmp01_23_81;
	wire [WIDTH*2-1+1:0] tmp01_23_82;
	wire [WIDTH*2-1+1:0] tmp01_23_83;
	wire [WIDTH*2-1+1:0] tmp01_24_0;
	wire [WIDTH*2-1+1:0] tmp01_24_1;
	wire [WIDTH*2-1+1:0] tmp01_24_2;
	wire [WIDTH*2-1+1:0] tmp01_24_3;
	wire [WIDTH*2-1+1:0] tmp01_24_4;
	wire [WIDTH*2-1+1:0] tmp01_24_5;
	wire [WIDTH*2-1+1:0] tmp01_24_6;
	wire [WIDTH*2-1+1:0] tmp01_24_7;
	wire [WIDTH*2-1+1:0] tmp01_24_8;
	wire [WIDTH*2-1+1:0] tmp01_24_9;
	wire [WIDTH*2-1+1:0] tmp01_24_10;
	wire [WIDTH*2-1+1:0] tmp01_24_11;
	wire [WIDTH*2-1+1:0] tmp01_24_12;
	wire [WIDTH*2-1+1:0] tmp01_24_13;
	wire [WIDTH*2-1+1:0] tmp01_24_14;
	wire [WIDTH*2-1+1:0] tmp01_24_15;
	wire [WIDTH*2-1+1:0] tmp01_24_16;
	wire [WIDTH*2-1+1:0] tmp01_24_17;
	wire [WIDTH*2-1+1:0] tmp01_24_18;
	wire [WIDTH*2-1+1:0] tmp01_24_19;
	wire [WIDTH*2-1+1:0] tmp01_24_20;
	wire [WIDTH*2-1+1:0] tmp01_24_21;
	wire [WIDTH*2-1+1:0] tmp01_24_22;
	wire [WIDTH*2-1+1:0] tmp01_24_23;
	wire [WIDTH*2-1+1:0] tmp01_24_24;
	wire [WIDTH*2-1+1:0] tmp01_24_25;
	wire [WIDTH*2-1+1:0] tmp01_24_26;
	wire [WIDTH*2-1+1:0] tmp01_24_27;
	wire [WIDTH*2-1+1:0] tmp01_24_28;
	wire [WIDTH*2-1+1:0] tmp01_24_29;
	wire [WIDTH*2-1+1:0] tmp01_24_30;
	wire [WIDTH*2-1+1:0] tmp01_24_31;
	wire [WIDTH*2-1+1:0] tmp01_24_32;
	wire [WIDTH*2-1+1:0] tmp01_24_33;
	wire [WIDTH*2-1+1:0] tmp01_24_34;
	wire [WIDTH*2-1+1:0] tmp01_24_35;
	wire [WIDTH*2-1+1:0] tmp01_24_36;
	wire [WIDTH*2-1+1:0] tmp01_24_37;
	wire [WIDTH*2-1+1:0] tmp01_24_38;
	wire [WIDTH*2-1+1:0] tmp01_24_39;
	wire [WIDTH*2-1+1:0] tmp01_24_40;
	wire [WIDTH*2-1+1:0] tmp01_24_41;
	wire [WIDTH*2-1+1:0] tmp01_24_42;
	wire [WIDTH*2-1+1:0] tmp01_24_43;
	wire [WIDTH*2-1+1:0] tmp01_24_44;
	wire [WIDTH*2-1+1:0] tmp01_24_45;
	wire [WIDTH*2-1+1:0] tmp01_24_46;
	wire [WIDTH*2-1+1:0] tmp01_24_47;
	wire [WIDTH*2-1+1:0] tmp01_24_48;
	wire [WIDTH*2-1+1:0] tmp01_24_49;
	wire [WIDTH*2-1+1:0] tmp01_24_50;
	wire [WIDTH*2-1+1:0] tmp01_24_51;
	wire [WIDTH*2-1+1:0] tmp01_24_52;
	wire [WIDTH*2-1+1:0] tmp01_24_53;
	wire [WIDTH*2-1+1:0] tmp01_24_54;
	wire [WIDTH*2-1+1:0] tmp01_24_55;
	wire [WIDTH*2-1+1:0] tmp01_24_56;
	wire [WIDTH*2-1+1:0] tmp01_24_57;
	wire [WIDTH*2-1+1:0] tmp01_24_58;
	wire [WIDTH*2-1+1:0] tmp01_24_59;
	wire [WIDTH*2-1+1:0] tmp01_24_60;
	wire [WIDTH*2-1+1:0] tmp01_24_61;
	wire [WIDTH*2-1+1:0] tmp01_24_62;
	wire [WIDTH*2-1+1:0] tmp01_24_63;
	wire [WIDTH*2-1+1:0] tmp01_24_64;
	wire [WIDTH*2-1+1:0] tmp01_24_65;
	wire [WIDTH*2-1+1:0] tmp01_24_66;
	wire [WIDTH*2-1+1:0] tmp01_24_67;
	wire [WIDTH*2-1+1:0] tmp01_24_68;
	wire [WIDTH*2-1+1:0] tmp01_24_69;
	wire [WIDTH*2-1+1:0] tmp01_24_70;
	wire [WIDTH*2-1+1:0] tmp01_24_71;
	wire [WIDTH*2-1+1:0] tmp01_24_72;
	wire [WIDTH*2-1+1:0] tmp01_24_73;
	wire [WIDTH*2-1+1:0] tmp01_24_74;
	wire [WIDTH*2-1+1:0] tmp01_24_75;
	wire [WIDTH*2-1+1:0] tmp01_24_76;
	wire [WIDTH*2-1+1:0] tmp01_24_77;
	wire [WIDTH*2-1+1:0] tmp01_24_78;
	wire [WIDTH*2-1+1:0] tmp01_24_79;
	wire [WIDTH*2-1+1:0] tmp01_24_80;
	wire [WIDTH*2-1+1:0] tmp01_24_81;
	wire [WIDTH*2-1+1:0] tmp01_24_82;
	wire [WIDTH*2-1+1:0] tmp01_24_83;
	wire [WIDTH*2-1+1:0] tmp01_25_0;
	wire [WIDTH*2-1+1:0] tmp01_25_1;
	wire [WIDTH*2-1+1:0] tmp01_25_2;
	wire [WIDTH*2-1+1:0] tmp01_25_3;
	wire [WIDTH*2-1+1:0] tmp01_25_4;
	wire [WIDTH*2-1+1:0] tmp01_25_5;
	wire [WIDTH*2-1+1:0] tmp01_25_6;
	wire [WIDTH*2-1+1:0] tmp01_25_7;
	wire [WIDTH*2-1+1:0] tmp01_25_8;
	wire [WIDTH*2-1+1:0] tmp01_25_9;
	wire [WIDTH*2-1+1:0] tmp01_25_10;
	wire [WIDTH*2-1+1:0] tmp01_25_11;
	wire [WIDTH*2-1+1:0] tmp01_25_12;
	wire [WIDTH*2-1+1:0] tmp01_25_13;
	wire [WIDTH*2-1+1:0] tmp01_25_14;
	wire [WIDTH*2-1+1:0] tmp01_25_15;
	wire [WIDTH*2-1+1:0] tmp01_25_16;
	wire [WIDTH*2-1+1:0] tmp01_25_17;
	wire [WIDTH*2-1+1:0] tmp01_25_18;
	wire [WIDTH*2-1+1:0] tmp01_25_19;
	wire [WIDTH*2-1+1:0] tmp01_25_20;
	wire [WIDTH*2-1+1:0] tmp01_25_21;
	wire [WIDTH*2-1+1:0] tmp01_25_22;
	wire [WIDTH*2-1+1:0] tmp01_25_23;
	wire [WIDTH*2-1+1:0] tmp01_25_24;
	wire [WIDTH*2-1+1:0] tmp01_25_25;
	wire [WIDTH*2-1+1:0] tmp01_25_26;
	wire [WIDTH*2-1+1:0] tmp01_25_27;
	wire [WIDTH*2-1+1:0] tmp01_25_28;
	wire [WIDTH*2-1+1:0] tmp01_25_29;
	wire [WIDTH*2-1+1:0] tmp01_25_30;
	wire [WIDTH*2-1+1:0] tmp01_25_31;
	wire [WIDTH*2-1+1:0] tmp01_25_32;
	wire [WIDTH*2-1+1:0] tmp01_25_33;
	wire [WIDTH*2-1+1:0] tmp01_25_34;
	wire [WIDTH*2-1+1:0] tmp01_25_35;
	wire [WIDTH*2-1+1:0] tmp01_25_36;
	wire [WIDTH*2-1+1:0] tmp01_25_37;
	wire [WIDTH*2-1+1:0] tmp01_25_38;
	wire [WIDTH*2-1+1:0] tmp01_25_39;
	wire [WIDTH*2-1+1:0] tmp01_25_40;
	wire [WIDTH*2-1+1:0] tmp01_25_41;
	wire [WIDTH*2-1+1:0] tmp01_25_42;
	wire [WIDTH*2-1+1:0] tmp01_25_43;
	wire [WIDTH*2-1+1:0] tmp01_25_44;
	wire [WIDTH*2-1+1:0] tmp01_25_45;
	wire [WIDTH*2-1+1:0] tmp01_25_46;
	wire [WIDTH*2-1+1:0] tmp01_25_47;
	wire [WIDTH*2-1+1:0] tmp01_25_48;
	wire [WIDTH*2-1+1:0] tmp01_25_49;
	wire [WIDTH*2-1+1:0] tmp01_25_50;
	wire [WIDTH*2-1+1:0] tmp01_25_51;
	wire [WIDTH*2-1+1:0] tmp01_25_52;
	wire [WIDTH*2-1+1:0] tmp01_25_53;
	wire [WIDTH*2-1+1:0] tmp01_25_54;
	wire [WIDTH*2-1+1:0] tmp01_25_55;
	wire [WIDTH*2-1+1:0] tmp01_25_56;
	wire [WIDTH*2-1+1:0] tmp01_25_57;
	wire [WIDTH*2-1+1:0] tmp01_25_58;
	wire [WIDTH*2-1+1:0] tmp01_25_59;
	wire [WIDTH*2-1+1:0] tmp01_25_60;
	wire [WIDTH*2-1+1:0] tmp01_25_61;
	wire [WIDTH*2-1+1:0] tmp01_25_62;
	wire [WIDTH*2-1+1:0] tmp01_25_63;
	wire [WIDTH*2-1+1:0] tmp01_25_64;
	wire [WIDTH*2-1+1:0] tmp01_25_65;
	wire [WIDTH*2-1+1:0] tmp01_25_66;
	wire [WIDTH*2-1+1:0] tmp01_25_67;
	wire [WIDTH*2-1+1:0] tmp01_25_68;
	wire [WIDTH*2-1+1:0] tmp01_25_69;
	wire [WIDTH*2-1+1:0] tmp01_25_70;
	wire [WIDTH*2-1+1:0] tmp01_25_71;
	wire [WIDTH*2-1+1:0] tmp01_25_72;
	wire [WIDTH*2-1+1:0] tmp01_25_73;
	wire [WIDTH*2-1+1:0] tmp01_25_74;
	wire [WIDTH*2-1+1:0] tmp01_25_75;
	wire [WIDTH*2-1+1:0] tmp01_25_76;
	wire [WIDTH*2-1+1:0] tmp01_25_77;
	wire [WIDTH*2-1+1:0] tmp01_25_78;
	wire [WIDTH*2-1+1:0] tmp01_25_79;
	wire [WIDTH*2-1+1:0] tmp01_25_80;
	wire [WIDTH*2-1+1:0] tmp01_25_81;
	wire [WIDTH*2-1+1:0] tmp01_25_82;
	wire [WIDTH*2-1+1:0] tmp01_25_83;
	wire [WIDTH*2-1+1:0] tmp01_26_0;
	wire [WIDTH*2-1+1:0] tmp01_26_1;
	wire [WIDTH*2-1+1:0] tmp01_26_2;
	wire [WIDTH*2-1+1:0] tmp01_26_3;
	wire [WIDTH*2-1+1:0] tmp01_26_4;
	wire [WIDTH*2-1+1:0] tmp01_26_5;
	wire [WIDTH*2-1+1:0] tmp01_26_6;
	wire [WIDTH*2-1+1:0] tmp01_26_7;
	wire [WIDTH*2-1+1:0] tmp01_26_8;
	wire [WIDTH*2-1+1:0] tmp01_26_9;
	wire [WIDTH*2-1+1:0] tmp01_26_10;
	wire [WIDTH*2-1+1:0] tmp01_26_11;
	wire [WIDTH*2-1+1:0] tmp01_26_12;
	wire [WIDTH*2-1+1:0] tmp01_26_13;
	wire [WIDTH*2-1+1:0] tmp01_26_14;
	wire [WIDTH*2-1+1:0] tmp01_26_15;
	wire [WIDTH*2-1+1:0] tmp01_26_16;
	wire [WIDTH*2-1+1:0] tmp01_26_17;
	wire [WIDTH*2-1+1:0] tmp01_26_18;
	wire [WIDTH*2-1+1:0] tmp01_26_19;
	wire [WIDTH*2-1+1:0] tmp01_26_20;
	wire [WIDTH*2-1+1:0] tmp01_26_21;
	wire [WIDTH*2-1+1:0] tmp01_26_22;
	wire [WIDTH*2-1+1:0] tmp01_26_23;
	wire [WIDTH*2-1+1:0] tmp01_26_24;
	wire [WIDTH*2-1+1:0] tmp01_26_25;
	wire [WIDTH*2-1+1:0] tmp01_26_26;
	wire [WIDTH*2-1+1:0] tmp01_26_27;
	wire [WIDTH*2-1+1:0] tmp01_26_28;
	wire [WIDTH*2-1+1:0] tmp01_26_29;
	wire [WIDTH*2-1+1:0] tmp01_26_30;
	wire [WIDTH*2-1+1:0] tmp01_26_31;
	wire [WIDTH*2-1+1:0] tmp01_26_32;
	wire [WIDTH*2-1+1:0] tmp01_26_33;
	wire [WIDTH*2-1+1:0] tmp01_26_34;
	wire [WIDTH*2-1+1:0] tmp01_26_35;
	wire [WIDTH*2-1+1:0] tmp01_26_36;
	wire [WIDTH*2-1+1:0] tmp01_26_37;
	wire [WIDTH*2-1+1:0] tmp01_26_38;
	wire [WIDTH*2-1+1:0] tmp01_26_39;
	wire [WIDTH*2-1+1:0] tmp01_26_40;
	wire [WIDTH*2-1+1:0] tmp01_26_41;
	wire [WIDTH*2-1+1:0] tmp01_26_42;
	wire [WIDTH*2-1+1:0] tmp01_26_43;
	wire [WIDTH*2-1+1:0] tmp01_26_44;
	wire [WIDTH*2-1+1:0] tmp01_26_45;
	wire [WIDTH*2-1+1:0] tmp01_26_46;
	wire [WIDTH*2-1+1:0] tmp01_26_47;
	wire [WIDTH*2-1+1:0] tmp01_26_48;
	wire [WIDTH*2-1+1:0] tmp01_26_49;
	wire [WIDTH*2-1+1:0] tmp01_26_50;
	wire [WIDTH*2-1+1:0] tmp01_26_51;
	wire [WIDTH*2-1+1:0] tmp01_26_52;
	wire [WIDTH*2-1+1:0] tmp01_26_53;
	wire [WIDTH*2-1+1:0] tmp01_26_54;
	wire [WIDTH*2-1+1:0] tmp01_26_55;
	wire [WIDTH*2-1+1:0] tmp01_26_56;
	wire [WIDTH*2-1+1:0] tmp01_26_57;
	wire [WIDTH*2-1+1:0] tmp01_26_58;
	wire [WIDTH*2-1+1:0] tmp01_26_59;
	wire [WIDTH*2-1+1:0] tmp01_26_60;
	wire [WIDTH*2-1+1:0] tmp01_26_61;
	wire [WIDTH*2-1+1:0] tmp01_26_62;
	wire [WIDTH*2-1+1:0] tmp01_26_63;
	wire [WIDTH*2-1+1:0] tmp01_26_64;
	wire [WIDTH*2-1+1:0] tmp01_26_65;
	wire [WIDTH*2-1+1:0] tmp01_26_66;
	wire [WIDTH*2-1+1:0] tmp01_26_67;
	wire [WIDTH*2-1+1:0] tmp01_26_68;
	wire [WIDTH*2-1+1:0] tmp01_26_69;
	wire [WIDTH*2-1+1:0] tmp01_26_70;
	wire [WIDTH*2-1+1:0] tmp01_26_71;
	wire [WIDTH*2-1+1:0] tmp01_26_72;
	wire [WIDTH*2-1+1:0] tmp01_26_73;
	wire [WIDTH*2-1+1:0] tmp01_26_74;
	wire [WIDTH*2-1+1:0] tmp01_26_75;
	wire [WIDTH*2-1+1:0] tmp01_26_76;
	wire [WIDTH*2-1+1:0] tmp01_26_77;
	wire [WIDTH*2-1+1:0] tmp01_26_78;
	wire [WIDTH*2-1+1:0] tmp01_26_79;
	wire [WIDTH*2-1+1:0] tmp01_26_80;
	wire [WIDTH*2-1+1:0] tmp01_26_81;
	wire [WIDTH*2-1+1:0] tmp01_26_82;
	wire [WIDTH*2-1+1:0] tmp01_26_83;
	wire [WIDTH*2-1+1:0] tmp01_27_0;
	wire [WIDTH*2-1+1:0] tmp01_27_1;
	wire [WIDTH*2-1+1:0] tmp01_27_2;
	wire [WIDTH*2-1+1:0] tmp01_27_3;
	wire [WIDTH*2-1+1:0] tmp01_27_4;
	wire [WIDTH*2-1+1:0] tmp01_27_5;
	wire [WIDTH*2-1+1:0] tmp01_27_6;
	wire [WIDTH*2-1+1:0] tmp01_27_7;
	wire [WIDTH*2-1+1:0] tmp01_27_8;
	wire [WIDTH*2-1+1:0] tmp01_27_9;
	wire [WIDTH*2-1+1:0] tmp01_27_10;
	wire [WIDTH*2-1+1:0] tmp01_27_11;
	wire [WIDTH*2-1+1:0] tmp01_27_12;
	wire [WIDTH*2-1+1:0] tmp01_27_13;
	wire [WIDTH*2-1+1:0] tmp01_27_14;
	wire [WIDTH*2-1+1:0] tmp01_27_15;
	wire [WIDTH*2-1+1:0] tmp01_27_16;
	wire [WIDTH*2-1+1:0] tmp01_27_17;
	wire [WIDTH*2-1+1:0] tmp01_27_18;
	wire [WIDTH*2-1+1:0] tmp01_27_19;
	wire [WIDTH*2-1+1:0] tmp01_27_20;
	wire [WIDTH*2-1+1:0] tmp01_27_21;
	wire [WIDTH*2-1+1:0] tmp01_27_22;
	wire [WIDTH*2-1+1:0] tmp01_27_23;
	wire [WIDTH*2-1+1:0] tmp01_27_24;
	wire [WIDTH*2-1+1:0] tmp01_27_25;
	wire [WIDTH*2-1+1:0] tmp01_27_26;
	wire [WIDTH*2-1+1:0] tmp01_27_27;
	wire [WIDTH*2-1+1:0] tmp01_27_28;
	wire [WIDTH*2-1+1:0] tmp01_27_29;
	wire [WIDTH*2-1+1:0] tmp01_27_30;
	wire [WIDTH*2-1+1:0] tmp01_27_31;
	wire [WIDTH*2-1+1:0] tmp01_27_32;
	wire [WIDTH*2-1+1:0] tmp01_27_33;
	wire [WIDTH*2-1+1:0] tmp01_27_34;
	wire [WIDTH*2-1+1:0] tmp01_27_35;
	wire [WIDTH*2-1+1:0] tmp01_27_36;
	wire [WIDTH*2-1+1:0] tmp01_27_37;
	wire [WIDTH*2-1+1:0] tmp01_27_38;
	wire [WIDTH*2-1+1:0] tmp01_27_39;
	wire [WIDTH*2-1+1:0] tmp01_27_40;
	wire [WIDTH*2-1+1:0] tmp01_27_41;
	wire [WIDTH*2-1+1:0] tmp01_27_42;
	wire [WIDTH*2-1+1:0] tmp01_27_43;
	wire [WIDTH*2-1+1:0] tmp01_27_44;
	wire [WIDTH*2-1+1:0] tmp01_27_45;
	wire [WIDTH*2-1+1:0] tmp01_27_46;
	wire [WIDTH*2-1+1:0] tmp01_27_47;
	wire [WIDTH*2-1+1:0] tmp01_27_48;
	wire [WIDTH*2-1+1:0] tmp01_27_49;
	wire [WIDTH*2-1+1:0] tmp01_27_50;
	wire [WIDTH*2-1+1:0] tmp01_27_51;
	wire [WIDTH*2-1+1:0] tmp01_27_52;
	wire [WIDTH*2-1+1:0] tmp01_27_53;
	wire [WIDTH*2-1+1:0] tmp01_27_54;
	wire [WIDTH*2-1+1:0] tmp01_27_55;
	wire [WIDTH*2-1+1:0] tmp01_27_56;
	wire [WIDTH*2-1+1:0] tmp01_27_57;
	wire [WIDTH*2-1+1:0] tmp01_27_58;
	wire [WIDTH*2-1+1:0] tmp01_27_59;
	wire [WIDTH*2-1+1:0] tmp01_27_60;
	wire [WIDTH*2-1+1:0] tmp01_27_61;
	wire [WIDTH*2-1+1:0] tmp01_27_62;
	wire [WIDTH*2-1+1:0] tmp01_27_63;
	wire [WIDTH*2-1+1:0] tmp01_27_64;
	wire [WIDTH*2-1+1:0] tmp01_27_65;
	wire [WIDTH*2-1+1:0] tmp01_27_66;
	wire [WIDTH*2-1+1:0] tmp01_27_67;
	wire [WIDTH*2-1+1:0] tmp01_27_68;
	wire [WIDTH*2-1+1:0] tmp01_27_69;
	wire [WIDTH*2-1+1:0] tmp01_27_70;
	wire [WIDTH*2-1+1:0] tmp01_27_71;
	wire [WIDTH*2-1+1:0] tmp01_27_72;
	wire [WIDTH*2-1+1:0] tmp01_27_73;
	wire [WIDTH*2-1+1:0] tmp01_27_74;
	wire [WIDTH*2-1+1:0] tmp01_27_75;
	wire [WIDTH*2-1+1:0] tmp01_27_76;
	wire [WIDTH*2-1+1:0] tmp01_27_77;
	wire [WIDTH*2-1+1:0] tmp01_27_78;
	wire [WIDTH*2-1+1:0] tmp01_27_79;
	wire [WIDTH*2-1+1:0] tmp01_27_80;
	wire [WIDTH*2-1+1:0] tmp01_27_81;
	wire [WIDTH*2-1+1:0] tmp01_27_82;
	wire [WIDTH*2-1+1:0] tmp01_27_83;
	wire [WIDTH*2-1+1:0] tmp01_28_0;
	wire [WIDTH*2-1+1:0] tmp01_28_1;
	wire [WIDTH*2-1+1:0] tmp01_28_2;
	wire [WIDTH*2-1+1:0] tmp01_28_3;
	wire [WIDTH*2-1+1:0] tmp01_28_4;
	wire [WIDTH*2-1+1:0] tmp01_28_5;
	wire [WIDTH*2-1+1:0] tmp01_28_6;
	wire [WIDTH*2-1+1:0] tmp01_28_7;
	wire [WIDTH*2-1+1:0] tmp01_28_8;
	wire [WIDTH*2-1+1:0] tmp01_28_9;
	wire [WIDTH*2-1+1:0] tmp01_28_10;
	wire [WIDTH*2-1+1:0] tmp01_28_11;
	wire [WIDTH*2-1+1:0] tmp01_28_12;
	wire [WIDTH*2-1+1:0] tmp01_28_13;
	wire [WIDTH*2-1+1:0] tmp01_28_14;
	wire [WIDTH*2-1+1:0] tmp01_28_15;
	wire [WIDTH*2-1+1:0] tmp01_28_16;
	wire [WIDTH*2-1+1:0] tmp01_28_17;
	wire [WIDTH*2-1+1:0] tmp01_28_18;
	wire [WIDTH*2-1+1:0] tmp01_28_19;
	wire [WIDTH*2-1+1:0] tmp01_28_20;
	wire [WIDTH*2-1+1:0] tmp01_28_21;
	wire [WIDTH*2-1+1:0] tmp01_28_22;
	wire [WIDTH*2-1+1:0] tmp01_28_23;
	wire [WIDTH*2-1+1:0] tmp01_28_24;
	wire [WIDTH*2-1+1:0] tmp01_28_25;
	wire [WIDTH*2-1+1:0] tmp01_28_26;
	wire [WIDTH*2-1+1:0] tmp01_28_27;
	wire [WIDTH*2-1+1:0] tmp01_28_28;
	wire [WIDTH*2-1+1:0] tmp01_28_29;
	wire [WIDTH*2-1+1:0] tmp01_28_30;
	wire [WIDTH*2-1+1:0] tmp01_28_31;
	wire [WIDTH*2-1+1:0] tmp01_28_32;
	wire [WIDTH*2-1+1:0] tmp01_28_33;
	wire [WIDTH*2-1+1:0] tmp01_28_34;
	wire [WIDTH*2-1+1:0] tmp01_28_35;
	wire [WIDTH*2-1+1:0] tmp01_28_36;
	wire [WIDTH*2-1+1:0] tmp01_28_37;
	wire [WIDTH*2-1+1:0] tmp01_28_38;
	wire [WIDTH*2-1+1:0] tmp01_28_39;
	wire [WIDTH*2-1+1:0] tmp01_28_40;
	wire [WIDTH*2-1+1:0] tmp01_28_41;
	wire [WIDTH*2-1+1:0] tmp01_28_42;
	wire [WIDTH*2-1+1:0] tmp01_28_43;
	wire [WIDTH*2-1+1:0] tmp01_28_44;
	wire [WIDTH*2-1+1:0] tmp01_28_45;
	wire [WIDTH*2-1+1:0] tmp01_28_46;
	wire [WIDTH*2-1+1:0] tmp01_28_47;
	wire [WIDTH*2-1+1:0] tmp01_28_48;
	wire [WIDTH*2-1+1:0] tmp01_28_49;
	wire [WIDTH*2-1+1:0] tmp01_28_50;
	wire [WIDTH*2-1+1:0] tmp01_28_51;
	wire [WIDTH*2-1+1:0] tmp01_28_52;
	wire [WIDTH*2-1+1:0] tmp01_28_53;
	wire [WIDTH*2-1+1:0] tmp01_28_54;
	wire [WIDTH*2-1+1:0] tmp01_28_55;
	wire [WIDTH*2-1+1:0] tmp01_28_56;
	wire [WIDTH*2-1+1:0] tmp01_28_57;
	wire [WIDTH*2-1+1:0] tmp01_28_58;
	wire [WIDTH*2-1+1:0] tmp01_28_59;
	wire [WIDTH*2-1+1:0] tmp01_28_60;
	wire [WIDTH*2-1+1:0] tmp01_28_61;
	wire [WIDTH*2-1+1:0] tmp01_28_62;
	wire [WIDTH*2-1+1:0] tmp01_28_63;
	wire [WIDTH*2-1+1:0] tmp01_28_64;
	wire [WIDTH*2-1+1:0] tmp01_28_65;
	wire [WIDTH*2-1+1:0] tmp01_28_66;
	wire [WIDTH*2-1+1:0] tmp01_28_67;
	wire [WIDTH*2-1+1:0] tmp01_28_68;
	wire [WIDTH*2-1+1:0] tmp01_28_69;
	wire [WIDTH*2-1+1:0] tmp01_28_70;
	wire [WIDTH*2-1+1:0] tmp01_28_71;
	wire [WIDTH*2-1+1:0] tmp01_28_72;
	wire [WIDTH*2-1+1:0] tmp01_28_73;
	wire [WIDTH*2-1+1:0] tmp01_28_74;
	wire [WIDTH*2-1+1:0] tmp01_28_75;
	wire [WIDTH*2-1+1:0] tmp01_28_76;
	wire [WIDTH*2-1+1:0] tmp01_28_77;
	wire [WIDTH*2-1+1:0] tmp01_28_78;
	wire [WIDTH*2-1+1:0] tmp01_28_79;
	wire [WIDTH*2-1+1:0] tmp01_28_80;
	wire [WIDTH*2-1+1:0] tmp01_28_81;
	wire [WIDTH*2-1+1:0] tmp01_28_82;
	wire [WIDTH*2-1+1:0] tmp01_28_83;
	wire [WIDTH*2-1+1:0] tmp01_29_0;
	wire [WIDTH*2-1+1:0] tmp01_29_1;
	wire [WIDTH*2-1+1:0] tmp01_29_2;
	wire [WIDTH*2-1+1:0] tmp01_29_3;
	wire [WIDTH*2-1+1:0] tmp01_29_4;
	wire [WIDTH*2-1+1:0] tmp01_29_5;
	wire [WIDTH*2-1+1:0] tmp01_29_6;
	wire [WIDTH*2-1+1:0] tmp01_29_7;
	wire [WIDTH*2-1+1:0] tmp01_29_8;
	wire [WIDTH*2-1+1:0] tmp01_29_9;
	wire [WIDTH*2-1+1:0] tmp01_29_10;
	wire [WIDTH*2-1+1:0] tmp01_29_11;
	wire [WIDTH*2-1+1:0] tmp01_29_12;
	wire [WIDTH*2-1+1:0] tmp01_29_13;
	wire [WIDTH*2-1+1:0] tmp01_29_14;
	wire [WIDTH*2-1+1:0] tmp01_29_15;
	wire [WIDTH*2-1+1:0] tmp01_29_16;
	wire [WIDTH*2-1+1:0] tmp01_29_17;
	wire [WIDTH*2-1+1:0] tmp01_29_18;
	wire [WIDTH*2-1+1:0] tmp01_29_19;
	wire [WIDTH*2-1+1:0] tmp01_29_20;
	wire [WIDTH*2-1+1:0] tmp01_29_21;
	wire [WIDTH*2-1+1:0] tmp01_29_22;
	wire [WIDTH*2-1+1:0] tmp01_29_23;
	wire [WIDTH*2-1+1:0] tmp01_29_24;
	wire [WIDTH*2-1+1:0] tmp01_29_25;
	wire [WIDTH*2-1+1:0] tmp01_29_26;
	wire [WIDTH*2-1+1:0] tmp01_29_27;
	wire [WIDTH*2-1+1:0] tmp01_29_28;
	wire [WIDTH*2-1+1:0] tmp01_29_29;
	wire [WIDTH*2-1+1:0] tmp01_29_30;
	wire [WIDTH*2-1+1:0] tmp01_29_31;
	wire [WIDTH*2-1+1:0] tmp01_29_32;
	wire [WIDTH*2-1+1:0] tmp01_29_33;
	wire [WIDTH*2-1+1:0] tmp01_29_34;
	wire [WIDTH*2-1+1:0] tmp01_29_35;
	wire [WIDTH*2-1+1:0] tmp01_29_36;
	wire [WIDTH*2-1+1:0] tmp01_29_37;
	wire [WIDTH*2-1+1:0] tmp01_29_38;
	wire [WIDTH*2-1+1:0] tmp01_29_39;
	wire [WIDTH*2-1+1:0] tmp01_29_40;
	wire [WIDTH*2-1+1:0] tmp01_29_41;
	wire [WIDTH*2-1+1:0] tmp01_29_42;
	wire [WIDTH*2-1+1:0] tmp01_29_43;
	wire [WIDTH*2-1+1:0] tmp01_29_44;
	wire [WIDTH*2-1+1:0] tmp01_29_45;
	wire [WIDTH*2-1+1:0] tmp01_29_46;
	wire [WIDTH*2-1+1:0] tmp01_29_47;
	wire [WIDTH*2-1+1:0] tmp01_29_48;
	wire [WIDTH*2-1+1:0] tmp01_29_49;
	wire [WIDTH*2-1+1:0] tmp01_29_50;
	wire [WIDTH*2-1+1:0] tmp01_29_51;
	wire [WIDTH*2-1+1:0] tmp01_29_52;
	wire [WIDTH*2-1+1:0] tmp01_29_53;
	wire [WIDTH*2-1+1:0] tmp01_29_54;
	wire [WIDTH*2-1+1:0] tmp01_29_55;
	wire [WIDTH*2-1+1:0] tmp01_29_56;
	wire [WIDTH*2-1+1:0] tmp01_29_57;
	wire [WIDTH*2-1+1:0] tmp01_29_58;
	wire [WIDTH*2-1+1:0] tmp01_29_59;
	wire [WIDTH*2-1+1:0] tmp01_29_60;
	wire [WIDTH*2-1+1:0] tmp01_29_61;
	wire [WIDTH*2-1+1:0] tmp01_29_62;
	wire [WIDTH*2-1+1:0] tmp01_29_63;
	wire [WIDTH*2-1+1:0] tmp01_29_64;
	wire [WIDTH*2-1+1:0] tmp01_29_65;
	wire [WIDTH*2-1+1:0] tmp01_29_66;
	wire [WIDTH*2-1+1:0] tmp01_29_67;
	wire [WIDTH*2-1+1:0] tmp01_29_68;
	wire [WIDTH*2-1+1:0] tmp01_29_69;
	wire [WIDTH*2-1+1:0] tmp01_29_70;
	wire [WIDTH*2-1+1:0] tmp01_29_71;
	wire [WIDTH*2-1+1:0] tmp01_29_72;
	wire [WIDTH*2-1+1:0] tmp01_29_73;
	wire [WIDTH*2-1+1:0] tmp01_29_74;
	wire [WIDTH*2-1+1:0] tmp01_29_75;
	wire [WIDTH*2-1+1:0] tmp01_29_76;
	wire [WIDTH*2-1+1:0] tmp01_29_77;
	wire [WIDTH*2-1+1:0] tmp01_29_78;
	wire [WIDTH*2-1+1:0] tmp01_29_79;
	wire [WIDTH*2-1+1:0] tmp01_29_80;
	wire [WIDTH*2-1+1:0] tmp01_29_81;
	wire [WIDTH*2-1+1:0] tmp01_29_82;
	wire [WIDTH*2-1+1:0] tmp01_29_83;
	wire [WIDTH*2-1+1:0] tmp01_30_0;
	wire [WIDTH*2-1+1:0] tmp01_30_1;
	wire [WIDTH*2-1+1:0] tmp01_30_2;
	wire [WIDTH*2-1+1:0] tmp01_30_3;
	wire [WIDTH*2-1+1:0] tmp01_30_4;
	wire [WIDTH*2-1+1:0] tmp01_30_5;
	wire [WIDTH*2-1+1:0] tmp01_30_6;
	wire [WIDTH*2-1+1:0] tmp01_30_7;
	wire [WIDTH*2-1+1:0] tmp01_30_8;
	wire [WIDTH*2-1+1:0] tmp01_30_9;
	wire [WIDTH*2-1+1:0] tmp01_30_10;
	wire [WIDTH*2-1+1:0] tmp01_30_11;
	wire [WIDTH*2-1+1:0] tmp01_30_12;
	wire [WIDTH*2-1+1:0] tmp01_30_13;
	wire [WIDTH*2-1+1:0] tmp01_30_14;
	wire [WIDTH*2-1+1:0] tmp01_30_15;
	wire [WIDTH*2-1+1:0] tmp01_30_16;
	wire [WIDTH*2-1+1:0] tmp01_30_17;
	wire [WIDTH*2-1+1:0] tmp01_30_18;
	wire [WIDTH*2-1+1:0] tmp01_30_19;
	wire [WIDTH*2-1+1:0] tmp01_30_20;
	wire [WIDTH*2-1+1:0] tmp01_30_21;
	wire [WIDTH*2-1+1:0] tmp01_30_22;
	wire [WIDTH*2-1+1:0] tmp01_30_23;
	wire [WIDTH*2-1+1:0] tmp01_30_24;
	wire [WIDTH*2-1+1:0] tmp01_30_25;
	wire [WIDTH*2-1+1:0] tmp01_30_26;
	wire [WIDTH*2-1+1:0] tmp01_30_27;
	wire [WIDTH*2-1+1:0] tmp01_30_28;
	wire [WIDTH*2-1+1:0] tmp01_30_29;
	wire [WIDTH*2-1+1:0] tmp01_30_30;
	wire [WIDTH*2-1+1:0] tmp01_30_31;
	wire [WIDTH*2-1+1:0] tmp01_30_32;
	wire [WIDTH*2-1+1:0] tmp01_30_33;
	wire [WIDTH*2-1+1:0] tmp01_30_34;
	wire [WIDTH*2-1+1:0] tmp01_30_35;
	wire [WIDTH*2-1+1:0] tmp01_30_36;
	wire [WIDTH*2-1+1:0] tmp01_30_37;
	wire [WIDTH*2-1+1:0] tmp01_30_38;
	wire [WIDTH*2-1+1:0] tmp01_30_39;
	wire [WIDTH*2-1+1:0] tmp01_30_40;
	wire [WIDTH*2-1+1:0] tmp01_30_41;
	wire [WIDTH*2-1+1:0] tmp01_30_42;
	wire [WIDTH*2-1+1:0] tmp01_30_43;
	wire [WIDTH*2-1+1:0] tmp01_30_44;
	wire [WIDTH*2-1+1:0] tmp01_30_45;
	wire [WIDTH*2-1+1:0] tmp01_30_46;
	wire [WIDTH*2-1+1:0] tmp01_30_47;
	wire [WIDTH*2-1+1:0] tmp01_30_48;
	wire [WIDTH*2-1+1:0] tmp01_30_49;
	wire [WIDTH*2-1+1:0] tmp01_30_50;
	wire [WIDTH*2-1+1:0] tmp01_30_51;
	wire [WIDTH*2-1+1:0] tmp01_30_52;
	wire [WIDTH*2-1+1:0] tmp01_30_53;
	wire [WIDTH*2-1+1:0] tmp01_30_54;
	wire [WIDTH*2-1+1:0] tmp01_30_55;
	wire [WIDTH*2-1+1:0] tmp01_30_56;
	wire [WIDTH*2-1+1:0] tmp01_30_57;
	wire [WIDTH*2-1+1:0] tmp01_30_58;
	wire [WIDTH*2-1+1:0] tmp01_30_59;
	wire [WIDTH*2-1+1:0] tmp01_30_60;
	wire [WIDTH*2-1+1:0] tmp01_30_61;
	wire [WIDTH*2-1+1:0] tmp01_30_62;
	wire [WIDTH*2-1+1:0] tmp01_30_63;
	wire [WIDTH*2-1+1:0] tmp01_30_64;
	wire [WIDTH*2-1+1:0] tmp01_30_65;
	wire [WIDTH*2-1+1:0] tmp01_30_66;
	wire [WIDTH*2-1+1:0] tmp01_30_67;
	wire [WIDTH*2-1+1:0] tmp01_30_68;
	wire [WIDTH*2-1+1:0] tmp01_30_69;
	wire [WIDTH*2-1+1:0] tmp01_30_70;
	wire [WIDTH*2-1+1:0] tmp01_30_71;
	wire [WIDTH*2-1+1:0] tmp01_30_72;
	wire [WIDTH*2-1+1:0] tmp01_30_73;
	wire [WIDTH*2-1+1:0] tmp01_30_74;
	wire [WIDTH*2-1+1:0] tmp01_30_75;
	wire [WIDTH*2-1+1:0] tmp01_30_76;
	wire [WIDTH*2-1+1:0] tmp01_30_77;
	wire [WIDTH*2-1+1:0] tmp01_30_78;
	wire [WIDTH*2-1+1:0] tmp01_30_79;
	wire [WIDTH*2-1+1:0] tmp01_30_80;
	wire [WIDTH*2-1+1:0] tmp01_30_81;
	wire [WIDTH*2-1+1:0] tmp01_30_82;
	wire [WIDTH*2-1+1:0] tmp01_30_83;
	wire [WIDTH*2-1+1:0] tmp01_31_0;
	wire [WIDTH*2-1+1:0] tmp01_31_1;
	wire [WIDTH*2-1+1:0] tmp01_31_2;
	wire [WIDTH*2-1+1:0] tmp01_31_3;
	wire [WIDTH*2-1+1:0] tmp01_31_4;
	wire [WIDTH*2-1+1:0] tmp01_31_5;
	wire [WIDTH*2-1+1:0] tmp01_31_6;
	wire [WIDTH*2-1+1:0] tmp01_31_7;
	wire [WIDTH*2-1+1:0] tmp01_31_8;
	wire [WIDTH*2-1+1:0] tmp01_31_9;
	wire [WIDTH*2-1+1:0] tmp01_31_10;
	wire [WIDTH*2-1+1:0] tmp01_31_11;
	wire [WIDTH*2-1+1:0] tmp01_31_12;
	wire [WIDTH*2-1+1:0] tmp01_31_13;
	wire [WIDTH*2-1+1:0] tmp01_31_14;
	wire [WIDTH*2-1+1:0] tmp01_31_15;
	wire [WIDTH*2-1+1:0] tmp01_31_16;
	wire [WIDTH*2-1+1:0] tmp01_31_17;
	wire [WIDTH*2-1+1:0] tmp01_31_18;
	wire [WIDTH*2-1+1:0] tmp01_31_19;
	wire [WIDTH*2-1+1:0] tmp01_31_20;
	wire [WIDTH*2-1+1:0] tmp01_31_21;
	wire [WIDTH*2-1+1:0] tmp01_31_22;
	wire [WIDTH*2-1+1:0] tmp01_31_23;
	wire [WIDTH*2-1+1:0] tmp01_31_24;
	wire [WIDTH*2-1+1:0] tmp01_31_25;
	wire [WIDTH*2-1+1:0] tmp01_31_26;
	wire [WIDTH*2-1+1:0] tmp01_31_27;
	wire [WIDTH*2-1+1:0] tmp01_31_28;
	wire [WIDTH*2-1+1:0] tmp01_31_29;
	wire [WIDTH*2-1+1:0] tmp01_31_30;
	wire [WIDTH*2-1+1:0] tmp01_31_31;
	wire [WIDTH*2-1+1:0] tmp01_31_32;
	wire [WIDTH*2-1+1:0] tmp01_31_33;
	wire [WIDTH*2-1+1:0] tmp01_31_34;
	wire [WIDTH*2-1+1:0] tmp01_31_35;
	wire [WIDTH*2-1+1:0] tmp01_31_36;
	wire [WIDTH*2-1+1:0] tmp01_31_37;
	wire [WIDTH*2-1+1:0] tmp01_31_38;
	wire [WIDTH*2-1+1:0] tmp01_31_39;
	wire [WIDTH*2-1+1:0] tmp01_31_40;
	wire [WIDTH*2-1+1:0] tmp01_31_41;
	wire [WIDTH*2-1+1:0] tmp01_31_42;
	wire [WIDTH*2-1+1:0] tmp01_31_43;
	wire [WIDTH*2-1+1:0] tmp01_31_44;
	wire [WIDTH*2-1+1:0] tmp01_31_45;
	wire [WIDTH*2-1+1:0] tmp01_31_46;
	wire [WIDTH*2-1+1:0] tmp01_31_47;
	wire [WIDTH*2-1+1:0] tmp01_31_48;
	wire [WIDTH*2-1+1:0] tmp01_31_49;
	wire [WIDTH*2-1+1:0] tmp01_31_50;
	wire [WIDTH*2-1+1:0] tmp01_31_51;
	wire [WIDTH*2-1+1:0] tmp01_31_52;
	wire [WIDTH*2-1+1:0] tmp01_31_53;
	wire [WIDTH*2-1+1:0] tmp01_31_54;
	wire [WIDTH*2-1+1:0] tmp01_31_55;
	wire [WIDTH*2-1+1:0] tmp01_31_56;
	wire [WIDTH*2-1+1:0] tmp01_31_57;
	wire [WIDTH*2-1+1:0] tmp01_31_58;
	wire [WIDTH*2-1+1:0] tmp01_31_59;
	wire [WIDTH*2-1+1:0] tmp01_31_60;
	wire [WIDTH*2-1+1:0] tmp01_31_61;
	wire [WIDTH*2-1+1:0] tmp01_31_62;
	wire [WIDTH*2-1+1:0] tmp01_31_63;
	wire [WIDTH*2-1+1:0] tmp01_31_64;
	wire [WIDTH*2-1+1:0] tmp01_31_65;
	wire [WIDTH*2-1+1:0] tmp01_31_66;
	wire [WIDTH*2-1+1:0] tmp01_31_67;
	wire [WIDTH*2-1+1:0] tmp01_31_68;
	wire [WIDTH*2-1+1:0] tmp01_31_69;
	wire [WIDTH*2-1+1:0] tmp01_31_70;
	wire [WIDTH*2-1+1:0] tmp01_31_71;
	wire [WIDTH*2-1+1:0] tmp01_31_72;
	wire [WIDTH*2-1+1:0] tmp01_31_73;
	wire [WIDTH*2-1+1:0] tmp01_31_74;
	wire [WIDTH*2-1+1:0] tmp01_31_75;
	wire [WIDTH*2-1+1:0] tmp01_31_76;
	wire [WIDTH*2-1+1:0] tmp01_31_77;
	wire [WIDTH*2-1+1:0] tmp01_31_78;
	wire [WIDTH*2-1+1:0] tmp01_31_79;
	wire [WIDTH*2-1+1:0] tmp01_31_80;
	wire [WIDTH*2-1+1:0] tmp01_31_81;
	wire [WIDTH*2-1+1:0] tmp01_31_82;
	wire [WIDTH*2-1+1:0] tmp01_31_83;
	wire [WIDTH*2-1+1:0] tmp01_32_0;
	wire [WIDTH*2-1+1:0] tmp01_32_1;
	wire [WIDTH*2-1+1:0] tmp01_32_2;
	wire [WIDTH*2-1+1:0] tmp01_32_3;
	wire [WIDTH*2-1+1:0] tmp01_32_4;
	wire [WIDTH*2-1+1:0] tmp01_32_5;
	wire [WIDTH*2-1+1:0] tmp01_32_6;
	wire [WIDTH*2-1+1:0] tmp01_32_7;
	wire [WIDTH*2-1+1:0] tmp01_32_8;
	wire [WIDTH*2-1+1:0] tmp01_32_9;
	wire [WIDTH*2-1+1:0] tmp01_32_10;
	wire [WIDTH*2-1+1:0] tmp01_32_11;
	wire [WIDTH*2-1+1:0] tmp01_32_12;
	wire [WIDTH*2-1+1:0] tmp01_32_13;
	wire [WIDTH*2-1+1:0] tmp01_32_14;
	wire [WIDTH*2-1+1:0] tmp01_32_15;
	wire [WIDTH*2-1+1:0] tmp01_32_16;
	wire [WIDTH*2-1+1:0] tmp01_32_17;
	wire [WIDTH*2-1+1:0] tmp01_32_18;
	wire [WIDTH*2-1+1:0] tmp01_32_19;
	wire [WIDTH*2-1+1:0] tmp01_32_20;
	wire [WIDTH*2-1+1:0] tmp01_32_21;
	wire [WIDTH*2-1+1:0] tmp01_32_22;
	wire [WIDTH*2-1+1:0] tmp01_32_23;
	wire [WIDTH*2-1+1:0] tmp01_32_24;
	wire [WIDTH*2-1+1:0] tmp01_32_25;
	wire [WIDTH*2-1+1:0] tmp01_32_26;
	wire [WIDTH*2-1+1:0] tmp01_32_27;
	wire [WIDTH*2-1+1:0] tmp01_32_28;
	wire [WIDTH*2-1+1:0] tmp01_32_29;
	wire [WIDTH*2-1+1:0] tmp01_32_30;
	wire [WIDTH*2-1+1:0] tmp01_32_31;
	wire [WIDTH*2-1+1:0] tmp01_32_32;
	wire [WIDTH*2-1+1:0] tmp01_32_33;
	wire [WIDTH*2-1+1:0] tmp01_32_34;
	wire [WIDTH*2-1+1:0] tmp01_32_35;
	wire [WIDTH*2-1+1:0] tmp01_32_36;
	wire [WIDTH*2-1+1:0] tmp01_32_37;
	wire [WIDTH*2-1+1:0] tmp01_32_38;
	wire [WIDTH*2-1+1:0] tmp01_32_39;
	wire [WIDTH*2-1+1:0] tmp01_32_40;
	wire [WIDTH*2-1+1:0] tmp01_32_41;
	wire [WIDTH*2-1+1:0] tmp01_32_42;
	wire [WIDTH*2-1+1:0] tmp01_32_43;
	wire [WIDTH*2-1+1:0] tmp01_32_44;
	wire [WIDTH*2-1+1:0] tmp01_32_45;
	wire [WIDTH*2-1+1:0] tmp01_32_46;
	wire [WIDTH*2-1+1:0] tmp01_32_47;
	wire [WIDTH*2-1+1:0] tmp01_32_48;
	wire [WIDTH*2-1+1:0] tmp01_32_49;
	wire [WIDTH*2-1+1:0] tmp01_32_50;
	wire [WIDTH*2-1+1:0] tmp01_32_51;
	wire [WIDTH*2-1+1:0] tmp01_32_52;
	wire [WIDTH*2-1+1:0] tmp01_32_53;
	wire [WIDTH*2-1+1:0] tmp01_32_54;
	wire [WIDTH*2-1+1:0] tmp01_32_55;
	wire [WIDTH*2-1+1:0] tmp01_32_56;
	wire [WIDTH*2-1+1:0] tmp01_32_57;
	wire [WIDTH*2-1+1:0] tmp01_32_58;
	wire [WIDTH*2-1+1:0] tmp01_32_59;
	wire [WIDTH*2-1+1:0] tmp01_32_60;
	wire [WIDTH*2-1+1:0] tmp01_32_61;
	wire [WIDTH*2-1+1:0] tmp01_32_62;
	wire [WIDTH*2-1+1:0] tmp01_32_63;
	wire [WIDTH*2-1+1:0] tmp01_32_64;
	wire [WIDTH*2-1+1:0] tmp01_32_65;
	wire [WIDTH*2-1+1:0] tmp01_32_66;
	wire [WIDTH*2-1+1:0] tmp01_32_67;
	wire [WIDTH*2-1+1:0] tmp01_32_68;
	wire [WIDTH*2-1+1:0] tmp01_32_69;
	wire [WIDTH*2-1+1:0] tmp01_32_70;
	wire [WIDTH*2-1+1:0] tmp01_32_71;
	wire [WIDTH*2-1+1:0] tmp01_32_72;
	wire [WIDTH*2-1+1:0] tmp01_32_73;
	wire [WIDTH*2-1+1:0] tmp01_32_74;
	wire [WIDTH*2-1+1:0] tmp01_32_75;
	wire [WIDTH*2-1+1:0] tmp01_32_76;
	wire [WIDTH*2-1+1:0] tmp01_32_77;
	wire [WIDTH*2-1+1:0] tmp01_32_78;
	wire [WIDTH*2-1+1:0] tmp01_32_79;
	wire [WIDTH*2-1+1:0] tmp01_32_80;
	wire [WIDTH*2-1+1:0] tmp01_32_81;
	wire [WIDTH*2-1+1:0] tmp01_32_82;
	wire [WIDTH*2-1+1:0] tmp01_32_83;
	wire [WIDTH*2-1+1:0] tmp01_33_0;
	wire [WIDTH*2-1+1:0] tmp01_33_1;
	wire [WIDTH*2-1+1:0] tmp01_33_2;
	wire [WIDTH*2-1+1:0] tmp01_33_3;
	wire [WIDTH*2-1+1:0] tmp01_33_4;
	wire [WIDTH*2-1+1:0] tmp01_33_5;
	wire [WIDTH*2-1+1:0] tmp01_33_6;
	wire [WIDTH*2-1+1:0] tmp01_33_7;
	wire [WIDTH*2-1+1:0] tmp01_33_8;
	wire [WIDTH*2-1+1:0] tmp01_33_9;
	wire [WIDTH*2-1+1:0] tmp01_33_10;
	wire [WIDTH*2-1+1:0] tmp01_33_11;
	wire [WIDTH*2-1+1:0] tmp01_33_12;
	wire [WIDTH*2-1+1:0] tmp01_33_13;
	wire [WIDTH*2-1+1:0] tmp01_33_14;
	wire [WIDTH*2-1+1:0] tmp01_33_15;
	wire [WIDTH*2-1+1:0] tmp01_33_16;
	wire [WIDTH*2-1+1:0] tmp01_33_17;
	wire [WIDTH*2-1+1:0] tmp01_33_18;
	wire [WIDTH*2-1+1:0] tmp01_33_19;
	wire [WIDTH*2-1+1:0] tmp01_33_20;
	wire [WIDTH*2-1+1:0] tmp01_33_21;
	wire [WIDTH*2-1+1:0] tmp01_33_22;
	wire [WIDTH*2-1+1:0] tmp01_33_23;
	wire [WIDTH*2-1+1:0] tmp01_33_24;
	wire [WIDTH*2-1+1:0] tmp01_33_25;
	wire [WIDTH*2-1+1:0] tmp01_33_26;
	wire [WIDTH*2-1+1:0] tmp01_33_27;
	wire [WIDTH*2-1+1:0] tmp01_33_28;
	wire [WIDTH*2-1+1:0] tmp01_33_29;
	wire [WIDTH*2-1+1:0] tmp01_33_30;
	wire [WIDTH*2-1+1:0] tmp01_33_31;
	wire [WIDTH*2-1+1:0] tmp01_33_32;
	wire [WIDTH*2-1+1:0] tmp01_33_33;
	wire [WIDTH*2-1+1:0] tmp01_33_34;
	wire [WIDTH*2-1+1:0] tmp01_33_35;
	wire [WIDTH*2-1+1:0] tmp01_33_36;
	wire [WIDTH*2-1+1:0] tmp01_33_37;
	wire [WIDTH*2-1+1:0] tmp01_33_38;
	wire [WIDTH*2-1+1:0] tmp01_33_39;
	wire [WIDTH*2-1+1:0] tmp01_33_40;
	wire [WIDTH*2-1+1:0] tmp01_33_41;
	wire [WIDTH*2-1+1:0] tmp01_33_42;
	wire [WIDTH*2-1+1:0] tmp01_33_43;
	wire [WIDTH*2-1+1:0] tmp01_33_44;
	wire [WIDTH*2-1+1:0] tmp01_33_45;
	wire [WIDTH*2-1+1:0] tmp01_33_46;
	wire [WIDTH*2-1+1:0] tmp01_33_47;
	wire [WIDTH*2-1+1:0] tmp01_33_48;
	wire [WIDTH*2-1+1:0] tmp01_33_49;
	wire [WIDTH*2-1+1:0] tmp01_33_50;
	wire [WIDTH*2-1+1:0] tmp01_33_51;
	wire [WIDTH*2-1+1:0] tmp01_33_52;
	wire [WIDTH*2-1+1:0] tmp01_33_53;
	wire [WIDTH*2-1+1:0] tmp01_33_54;
	wire [WIDTH*2-1+1:0] tmp01_33_55;
	wire [WIDTH*2-1+1:0] tmp01_33_56;
	wire [WIDTH*2-1+1:0] tmp01_33_57;
	wire [WIDTH*2-1+1:0] tmp01_33_58;
	wire [WIDTH*2-1+1:0] tmp01_33_59;
	wire [WIDTH*2-1+1:0] tmp01_33_60;
	wire [WIDTH*2-1+1:0] tmp01_33_61;
	wire [WIDTH*2-1+1:0] tmp01_33_62;
	wire [WIDTH*2-1+1:0] tmp01_33_63;
	wire [WIDTH*2-1+1:0] tmp01_33_64;
	wire [WIDTH*2-1+1:0] tmp01_33_65;
	wire [WIDTH*2-1+1:0] tmp01_33_66;
	wire [WIDTH*2-1+1:0] tmp01_33_67;
	wire [WIDTH*2-1+1:0] tmp01_33_68;
	wire [WIDTH*2-1+1:0] tmp01_33_69;
	wire [WIDTH*2-1+1:0] tmp01_33_70;
	wire [WIDTH*2-1+1:0] tmp01_33_71;
	wire [WIDTH*2-1+1:0] tmp01_33_72;
	wire [WIDTH*2-1+1:0] tmp01_33_73;
	wire [WIDTH*2-1+1:0] tmp01_33_74;
	wire [WIDTH*2-1+1:0] tmp01_33_75;
	wire [WIDTH*2-1+1:0] tmp01_33_76;
	wire [WIDTH*2-1+1:0] tmp01_33_77;
	wire [WIDTH*2-1+1:0] tmp01_33_78;
	wire [WIDTH*2-1+1:0] tmp01_33_79;
	wire [WIDTH*2-1+1:0] tmp01_33_80;
	wire [WIDTH*2-1+1:0] tmp01_33_81;
	wire [WIDTH*2-1+1:0] tmp01_33_82;
	wire [WIDTH*2-1+1:0] tmp01_33_83;
	wire [WIDTH*2-1+1:0] tmp01_34_0;
	wire [WIDTH*2-1+1:0] tmp01_34_1;
	wire [WIDTH*2-1+1:0] tmp01_34_2;
	wire [WIDTH*2-1+1:0] tmp01_34_3;
	wire [WIDTH*2-1+1:0] tmp01_34_4;
	wire [WIDTH*2-1+1:0] tmp01_34_5;
	wire [WIDTH*2-1+1:0] tmp01_34_6;
	wire [WIDTH*2-1+1:0] tmp01_34_7;
	wire [WIDTH*2-1+1:0] tmp01_34_8;
	wire [WIDTH*2-1+1:0] tmp01_34_9;
	wire [WIDTH*2-1+1:0] tmp01_34_10;
	wire [WIDTH*2-1+1:0] tmp01_34_11;
	wire [WIDTH*2-1+1:0] tmp01_34_12;
	wire [WIDTH*2-1+1:0] tmp01_34_13;
	wire [WIDTH*2-1+1:0] tmp01_34_14;
	wire [WIDTH*2-1+1:0] tmp01_34_15;
	wire [WIDTH*2-1+1:0] tmp01_34_16;
	wire [WIDTH*2-1+1:0] tmp01_34_17;
	wire [WIDTH*2-1+1:0] tmp01_34_18;
	wire [WIDTH*2-1+1:0] tmp01_34_19;
	wire [WIDTH*2-1+1:0] tmp01_34_20;
	wire [WIDTH*2-1+1:0] tmp01_34_21;
	wire [WIDTH*2-1+1:0] tmp01_34_22;
	wire [WIDTH*2-1+1:0] tmp01_34_23;
	wire [WIDTH*2-1+1:0] tmp01_34_24;
	wire [WIDTH*2-1+1:0] tmp01_34_25;
	wire [WIDTH*2-1+1:0] tmp01_34_26;
	wire [WIDTH*2-1+1:0] tmp01_34_27;
	wire [WIDTH*2-1+1:0] tmp01_34_28;
	wire [WIDTH*2-1+1:0] tmp01_34_29;
	wire [WIDTH*2-1+1:0] tmp01_34_30;
	wire [WIDTH*2-1+1:0] tmp01_34_31;
	wire [WIDTH*2-1+1:0] tmp01_34_32;
	wire [WIDTH*2-1+1:0] tmp01_34_33;
	wire [WIDTH*2-1+1:0] tmp01_34_34;
	wire [WIDTH*2-1+1:0] tmp01_34_35;
	wire [WIDTH*2-1+1:0] tmp01_34_36;
	wire [WIDTH*2-1+1:0] tmp01_34_37;
	wire [WIDTH*2-1+1:0] tmp01_34_38;
	wire [WIDTH*2-1+1:0] tmp01_34_39;
	wire [WIDTH*2-1+1:0] tmp01_34_40;
	wire [WIDTH*2-1+1:0] tmp01_34_41;
	wire [WIDTH*2-1+1:0] tmp01_34_42;
	wire [WIDTH*2-1+1:0] tmp01_34_43;
	wire [WIDTH*2-1+1:0] tmp01_34_44;
	wire [WIDTH*2-1+1:0] tmp01_34_45;
	wire [WIDTH*2-1+1:0] tmp01_34_46;
	wire [WIDTH*2-1+1:0] tmp01_34_47;
	wire [WIDTH*2-1+1:0] tmp01_34_48;
	wire [WIDTH*2-1+1:0] tmp01_34_49;
	wire [WIDTH*2-1+1:0] tmp01_34_50;
	wire [WIDTH*2-1+1:0] tmp01_34_51;
	wire [WIDTH*2-1+1:0] tmp01_34_52;
	wire [WIDTH*2-1+1:0] tmp01_34_53;
	wire [WIDTH*2-1+1:0] tmp01_34_54;
	wire [WIDTH*2-1+1:0] tmp01_34_55;
	wire [WIDTH*2-1+1:0] tmp01_34_56;
	wire [WIDTH*2-1+1:0] tmp01_34_57;
	wire [WIDTH*2-1+1:0] tmp01_34_58;
	wire [WIDTH*2-1+1:0] tmp01_34_59;
	wire [WIDTH*2-1+1:0] tmp01_34_60;
	wire [WIDTH*2-1+1:0] tmp01_34_61;
	wire [WIDTH*2-1+1:0] tmp01_34_62;
	wire [WIDTH*2-1+1:0] tmp01_34_63;
	wire [WIDTH*2-1+1:0] tmp01_34_64;
	wire [WIDTH*2-1+1:0] tmp01_34_65;
	wire [WIDTH*2-1+1:0] tmp01_34_66;
	wire [WIDTH*2-1+1:0] tmp01_34_67;
	wire [WIDTH*2-1+1:0] tmp01_34_68;
	wire [WIDTH*2-1+1:0] tmp01_34_69;
	wire [WIDTH*2-1+1:0] tmp01_34_70;
	wire [WIDTH*2-1+1:0] tmp01_34_71;
	wire [WIDTH*2-1+1:0] tmp01_34_72;
	wire [WIDTH*2-1+1:0] tmp01_34_73;
	wire [WIDTH*2-1+1:0] tmp01_34_74;
	wire [WIDTH*2-1+1:0] tmp01_34_75;
	wire [WIDTH*2-1+1:0] tmp01_34_76;
	wire [WIDTH*2-1+1:0] tmp01_34_77;
	wire [WIDTH*2-1+1:0] tmp01_34_78;
	wire [WIDTH*2-1+1:0] tmp01_34_79;
	wire [WIDTH*2-1+1:0] tmp01_34_80;
	wire [WIDTH*2-1+1:0] tmp01_34_81;
	wire [WIDTH*2-1+1:0] tmp01_34_82;
	wire [WIDTH*2-1+1:0] tmp01_34_83;
	wire [WIDTH*2-1+1:0] tmp01_35_0;
	wire [WIDTH*2-1+1:0] tmp01_35_1;
	wire [WIDTH*2-1+1:0] tmp01_35_2;
	wire [WIDTH*2-1+1:0] tmp01_35_3;
	wire [WIDTH*2-1+1:0] tmp01_35_4;
	wire [WIDTH*2-1+1:0] tmp01_35_5;
	wire [WIDTH*2-1+1:0] tmp01_35_6;
	wire [WIDTH*2-1+1:0] tmp01_35_7;
	wire [WIDTH*2-1+1:0] tmp01_35_8;
	wire [WIDTH*2-1+1:0] tmp01_35_9;
	wire [WIDTH*2-1+1:0] tmp01_35_10;
	wire [WIDTH*2-1+1:0] tmp01_35_11;
	wire [WIDTH*2-1+1:0] tmp01_35_12;
	wire [WIDTH*2-1+1:0] tmp01_35_13;
	wire [WIDTH*2-1+1:0] tmp01_35_14;
	wire [WIDTH*2-1+1:0] tmp01_35_15;
	wire [WIDTH*2-1+1:0] tmp01_35_16;
	wire [WIDTH*2-1+1:0] tmp01_35_17;
	wire [WIDTH*2-1+1:0] tmp01_35_18;
	wire [WIDTH*2-1+1:0] tmp01_35_19;
	wire [WIDTH*2-1+1:0] tmp01_35_20;
	wire [WIDTH*2-1+1:0] tmp01_35_21;
	wire [WIDTH*2-1+1:0] tmp01_35_22;
	wire [WIDTH*2-1+1:0] tmp01_35_23;
	wire [WIDTH*2-1+1:0] tmp01_35_24;
	wire [WIDTH*2-1+1:0] tmp01_35_25;
	wire [WIDTH*2-1+1:0] tmp01_35_26;
	wire [WIDTH*2-1+1:0] tmp01_35_27;
	wire [WIDTH*2-1+1:0] tmp01_35_28;
	wire [WIDTH*2-1+1:0] tmp01_35_29;
	wire [WIDTH*2-1+1:0] tmp01_35_30;
	wire [WIDTH*2-1+1:0] tmp01_35_31;
	wire [WIDTH*2-1+1:0] tmp01_35_32;
	wire [WIDTH*2-1+1:0] tmp01_35_33;
	wire [WIDTH*2-1+1:0] tmp01_35_34;
	wire [WIDTH*2-1+1:0] tmp01_35_35;
	wire [WIDTH*2-1+1:0] tmp01_35_36;
	wire [WIDTH*2-1+1:0] tmp01_35_37;
	wire [WIDTH*2-1+1:0] tmp01_35_38;
	wire [WIDTH*2-1+1:0] tmp01_35_39;
	wire [WIDTH*2-1+1:0] tmp01_35_40;
	wire [WIDTH*2-1+1:0] tmp01_35_41;
	wire [WIDTH*2-1+1:0] tmp01_35_42;
	wire [WIDTH*2-1+1:0] tmp01_35_43;
	wire [WIDTH*2-1+1:0] tmp01_35_44;
	wire [WIDTH*2-1+1:0] tmp01_35_45;
	wire [WIDTH*2-1+1:0] tmp01_35_46;
	wire [WIDTH*2-1+1:0] tmp01_35_47;
	wire [WIDTH*2-1+1:0] tmp01_35_48;
	wire [WIDTH*2-1+1:0] tmp01_35_49;
	wire [WIDTH*2-1+1:0] tmp01_35_50;
	wire [WIDTH*2-1+1:0] tmp01_35_51;
	wire [WIDTH*2-1+1:0] tmp01_35_52;
	wire [WIDTH*2-1+1:0] tmp01_35_53;
	wire [WIDTH*2-1+1:0] tmp01_35_54;
	wire [WIDTH*2-1+1:0] tmp01_35_55;
	wire [WIDTH*2-1+1:0] tmp01_35_56;
	wire [WIDTH*2-1+1:0] tmp01_35_57;
	wire [WIDTH*2-1+1:0] tmp01_35_58;
	wire [WIDTH*2-1+1:0] tmp01_35_59;
	wire [WIDTH*2-1+1:0] tmp01_35_60;
	wire [WIDTH*2-1+1:0] tmp01_35_61;
	wire [WIDTH*2-1+1:0] tmp01_35_62;
	wire [WIDTH*2-1+1:0] tmp01_35_63;
	wire [WIDTH*2-1+1:0] tmp01_35_64;
	wire [WIDTH*2-1+1:0] tmp01_35_65;
	wire [WIDTH*2-1+1:0] tmp01_35_66;
	wire [WIDTH*2-1+1:0] tmp01_35_67;
	wire [WIDTH*2-1+1:0] tmp01_35_68;
	wire [WIDTH*2-1+1:0] tmp01_35_69;
	wire [WIDTH*2-1+1:0] tmp01_35_70;
	wire [WIDTH*2-1+1:0] tmp01_35_71;
	wire [WIDTH*2-1+1:0] tmp01_35_72;
	wire [WIDTH*2-1+1:0] tmp01_35_73;
	wire [WIDTH*2-1+1:0] tmp01_35_74;
	wire [WIDTH*2-1+1:0] tmp01_35_75;
	wire [WIDTH*2-1+1:0] tmp01_35_76;
	wire [WIDTH*2-1+1:0] tmp01_35_77;
	wire [WIDTH*2-1+1:0] tmp01_35_78;
	wire [WIDTH*2-1+1:0] tmp01_35_79;
	wire [WIDTH*2-1+1:0] tmp01_35_80;
	wire [WIDTH*2-1+1:0] tmp01_35_81;
	wire [WIDTH*2-1+1:0] tmp01_35_82;
	wire [WIDTH*2-1+1:0] tmp01_35_83;
	wire [WIDTH*2-1+1:0] tmp01_36_0;
	wire [WIDTH*2-1+1:0] tmp01_36_1;
	wire [WIDTH*2-1+1:0] tmp01_36_2;
	wire [WIDTH*2-1+1:0] tmp01_36_3;
	wire [WIDTH*2-1+1:0] tmp01_36_4;
	wire [WIDTH*2-1+1:0] tmp01_36_5;
	wire [WIDTH*2-1+1:0] tmp01_36_6;
	wire [WIDTH*2-1+1:0] tmp01_36_7;
	wire [WIDTH*2-1+1:0] tmp01_36_8;
	wire [WIDTH*2-1+1:0] tmp01_36_9;
	wire [WIDTH*2-1+1:0] tmp01_36_10;
	wire [WIDTH*2-1+1:0] tmp01_36_11;
	wire [WIDTH*2-1+1:0] tmp01_36_12;
	wire [WIDTH*2-1+1:0] tmp01_36_13;
	wire [WIDTH*2-1+1:0] tmp01_36_14;
	wire [WIDTH*2-1+1:0] tmp01_36_15;
	wire [WIDTH*2-1+1:0] tmp01_36_16;
	wire [WIDTH*2-1+1:0] tmp01_36_17;
	wire [WIDTH*2-1+1:0] tmp01_36_18;
	wire [WIDTH*2-1+1:0] tmp01_36_19;
	wire [WIDTH*2-1+1:0] tmp01_36_20;
	wire [WIDTH*2-1+1:0] tmp01_36_21;
	wire [WIDTH*2-1+1:0] tmp01_36_22;
	wire [WIDTH*2-1+1:0] tmp01_36_23;
	wire [WIDTH*2-1+1:0] tmp01_36_24;
	wire [WIDTH*2-1+1:0] tmp01_36_25;
	wire [WIDTH*2-1+1:0] tmp01_36_26;
	wire [WIDTH*2-1+1:0] tmp01_36_27;
	wire [WIDTH*2-1+1:0] tmp01_36_28;
	wire [WIDTH*2-1+1:0] tmp01_36_29;
	wire [WIDTH*2-1+1:0] tmp01_36_30;
	wire [WIDTH*2-1+1:0] tmp01_36_31;
	wire [WIDTH*2-1+1:0] tmp01_36_32;
	wire [WIDTH*2-1+1:0] tmp01_36_33;
	wire [WIDTH*2-1+1:0] tmp01_36_34;
	wire [WIDTH*2-1+1:0] tmp01_36_35;
	wire [WIDTH*2-1+1:0] tmp01_36_36;
	wire [WIDTH*2-1+1:0] tmp01_36_37;
	wire [WIDTH*2-1+1:0] tmp01_36_38;
	wire [WIDTH*2-1+1:0] tmp01_36_39;
	wire [WIDTH*2-1+1:0] tmp01_36_40;
	wire [WIDTH*2-1+1:0] tmp01_36_41;
	wire [WIDTH*2-1+1:0] tmp01_36_42;
	wire [WIDTH*2-1+1:0] tmp01_36_43;
	wire [WIDTH*2-1+1:0] tmp01_36_44;
	wire [WIDTH*2-1+1:0] tmp01_36_45;
	wire [WIDTH*2-1+1:0] tmp01_36_46;
	wire [WIDTH*2-1+1:0] tmp01_36_47;
	wire [WIDTH*2-1+1:0] tmp01_36_48;
	wire [WIDTH*2-1+1:0] tmp01_36_49;
	wire [WIDTH*2-1+1:0] tmp01_36_50;
	wire [WIDTH*2-1+1:0] tmp01_36_51;
	wire [WIDTH*2-1+1:0] tmp01_36_52;
	wire [WIDTH*2-1+1:0] tmp01_36_53;
	wire [WIDTH*2-1+1:0] tmp01_36_54;
	wire [WIDTH*2-1+1:0] tmp01_36_55;
	wire [WIDTH*2-1+1:0] tmp01_36_56;
	wire [WIDTH*2-1+1:0] tmp01_36_57;
	wire [WIDTH*2-1+1:0] tmp01_36_58;
	wire [WIDTH*2-1+1:0] tmp01_36_59;
	wire [WIDTH*2-1+1:0] tmp01_36_60;
	wire [WIDTH*2-1+1:0] tmp01_36_61;
	wire [WIDTH*2-1+1:0] tmp01_36_62;
	wire [WIDTH*2-1+1:0] tmp01_36_63;
	wire [WIDTH*2-1+1:0] tmp01_36_64;
	wire [WIDTH*2-1+1:0] tmp01_36_65;
	wire [WIDTH*2-1+1:0] tmp01_36_66;
	wire [WIDTH*2-1+1:0] tmp01_36_67;
	wire [WIDTH*2-1+1:0] tmp01_36_68;
	wire [WIDTH*2-1+1:0] tmp01_36_69;
	wire [WIDTH*2-1+1:0] tmp01_36_70;
	wire [WIDTH*2-1+1:0] tmp01_36_71;
	wire [WIDTH*2-1+1:0] tmp01_36_72;
	wire [WIDTH*2-1+1:0] tmp01_36_73;
	wire [WIDTH*2-1+1:0] tmp01_36_74;
	wire [WIDTH*2-1+1:0] tmp01_36_75;
	wire [WIDTH*2-1+1:0] tmp01_36_76;
	wire [WIDTH*2-1+1:0] tmp01_36_77;
	wire [WIDTH*2-1+1:0] tmp01_36_78;
	wire [WIDTH*2-1+1:0] tmp01_36_79;
	wire [WIDTH*2-1+1:0] tmp01_36_80;
	wire [WIDTH*2-1+1:0] tmp01_36_81;
	wire [WIDTH*2-1+1:0] tmp01_36_82;
	wire [WIDTH*2-1+1:0] tmp01_36_83;
	wire [WIDTH*2-1+1:0] tmp01_37_0;
	wire [WIDTH*2-1+1:0] tmp01_37_1;
	wire [WIDTH*2-1+1:0] tmp01_37_2;
	wire [WIDTH*2-1+1:0] tmp01_37_3;
	wire [WIDTH*2-1+1:0] tmp01_37_4;
	wire [WIDTH*2-1+1:0] tmp01_37_5;
	wire [WIDTH*2-1+1:0] tmp01_37_6;
	wire [WIDTH*2-1+1:0] tmp01_37_7;
	wire [WIDTH*2-1+1:0] tmp01_37_8;
	wire [WIDTH*2-1+1:0] tmp01_37_9;
	wire [WIDTH*2-1+1:0] tmp01_37_10;
	wire [WIDTH*2-1+1:0] tmp01_37_11;
	wire [WIDTH*2-1+1:0] tmp01_37_12;
	wire [WIDTH*2-1+1:0] tmp01_37_13;
	wire [WIDTH*2-1+1:0] tmp01_37_14;
	wire [WIDTH*2-1+1:0] tmp01_37_15;
	wire [WIDTH*2-1+1:0] tmp01_37_16;
	wire [WIDTH*2-1+1:0] tmp01_37_17;
	wire [WIDTH*2-1+1:0] tmp01_37_18;
	wire [WIDTH*2-1+1:0] tmp01_37_19;
	wire [WIDTH*2-1+1:0] tmp01_37_20;
	wire [WIDTH*2-1+1:0] tmp01_37_21;
	wire [WIDTH*2-1+1:0] tmp01_37_22;
	wire [WIDTH*2-1+1:0] tmp01_37_23;
	wire [WIDTH*2-1+1:0] tmp01_37_24;
	wire [WIDTH*2-1+1:0] tmp01_37_25;
	wire [WIDTH*2-1+1:0] tmp01_37_26;
	wire [WIDTH*2-1+1:0] tmp01_37_27;
	wire [WIDTH*2-1+1:0] tmp01_37_28;
	wire [WIDTH*2-1+1:0] tmp01_37_29;
	wire [WIDTH*2-1+1:0] tmp01_37_30;
	wire [WIDTH*2-1+1:0] tmp01_37_31;
	wire [WIDTH*2-1+1:0] tmp01_37_32;
	wire [WIDTH*2-1+1:0] tmp01_37_33;
	wire [WIDTH*2-1+1:0] tmp01_37_34;
	wire [WIDTH*2-1+1:0] tmp01_37_35;
	wire [WIDTH*2-1+1:0] tmp01_37_36;
	wire [WIDTH*2-1+1:0] tmp01_37_37;
	wire [WIDTH*2-1+1:0] tmp01_37_38;
	wire [WIDTH*2-1+1:0] tmp01_37_39;
	wire [WIDTH*2-1+1:0] tmp01_37_40;
	wire [WIDTH*2-1+1:0] tmp01_37_41;
	wire [WIDTH*2-1+1:0] tmp01_37_42;
	wire [WIDTH*2-1+1:0] tmp01_37_43;
	wire [WIDTH*2-1+1:0] tmp01_37_44;
	wire [WIDTH*2-1+1:0] tmp01_37_45;
	wire [WIDTH*2-1+1:0] tmp01_37_46;
	wire [WIDTH*2-1+1:0] tmp01_37_47;
	wire [WIDTH*2-1+1:0] tmp01_37_48;
	wire [WIDTH*2-1+1:0] tmp01_37_49;
	wire [WIDTH*2-1+1:0] tmp01_37_50;
	wire [WIDTH*2-1+1:0] tmp01_37_51;
	wire [WIDTH*2-1+1:0] tmp01_37_52;
	wire [WIDTH*2-1+1:0] tmp01_37_53;
	wire [WIDTH*2-1+1:0] tmp01_37_54;
	wire [WIDTH*2-1+1:0] tmp01_37_55;
	wire [WIDTH*2-1+1:0] tmp01_37_56;
	wire [WIDTH*2-1+1:0] tmp01_37_57;
	wire [WIDTH*2-1+1:0] tmp01_37_58;
	wire [WIDTH*2-1+1:0] tmp01_37_59;
	wire [WIDTH*2-1+1:0] tmp01_37_60;
	wire [WIDTH*2-1+1:0] tmp01_37_61;
	wire [WIDTH*2-1+1:0] tmp01_37_62;
	wire [WIDTH*2-1+1:0] tmp01_37_63;
	wire [WIDTH*2-1+1:0] tmp01_37_64;
	wire [WIDTH*2-1+1:0] tmp01_37_65;
	wire [WIDTH*2-1+1:0] tmp01_37_66;
	wire [WIDTH*2-1+1:0] tmp01_37_67;
	wire [WIDTH*2-1+1:0] tmp01_37_68;
	wire [WIDTH*2-1+1:0] tmp01_37_69;
	wire [WIDTH*2-1+1:0] tmp01_37_70;
	wire [WIDTH*2-1+1:0] tmp01_37_71;
	wire [WIDTH*2-1+1:0] tmp01_37_72;
	wire [WIDTH*2-1+1:0] tmp01_37_73;
	wire [WIDTH*2-1+1:0] tmp01_37_74;
	wire [WIDTH*2-1+1:0] tmp01_37_75;
	wire [WIDTH*2-1+1:0] tmp01_37_76;
	wire [WIDTH*2-1+1:0] tmp01_37_77;
	wire [WIDTH*2-1+1:0] tmp01_37_78;
	wire [WIDTH*2-1+1:0] tmp01_37_79;
	wire [WIDTH*2-1+1:0] tmp01_37_80;
	wire [WIDTH*2-1+1:0] tmp01_37_81;
	wire [WIDTH*2-1+1:0] tmp01_37_82;
	wire [WIDTH*2-1+1:0] tmp01_37_83;
	wire [WIDTH*2-1+1:0] tmp01_38_0;
	wire [WIDTH*2-1+1:0] tmp01_38_1;
	wire [WIDTH*2-1+1:0] tmp01_38_2;
	wire [WIDTH*2-1+1:0] tmp01_38_3;
	wire [WIDTH*2-1+1:0] tmp01_38_4;
	wire [WIDTH*2-1+1:0] tmp01_38_5;
	wire [WIDTH*2-1+1:0] tmp01_38_6;
	wire [WIDTH*2-1+1:0] tmp01_38_7;
	wire [WIDTH*2-1+1:0] tmp01_38_8;
	wire [WIDTH*2-1+1:0] tmp01_38_9;
	wire [WIDTH*2-1+1:0] tmp01_38_10;
	wire [WIDTH*2-1+1:0] tmp01_38_11;
	wire [WIDTH*2-1+1:0] tmp01_38_12;
	wire [WIDTH*2-1+1:0] tmp01_38_13;
	wire [WIDTH*2-1+1:0] tmp01_38_14;
	wire [WIDTH*2-1+1:0] tmp01_38_15;
	wire [WIDTH*2-1+1:0] tmp01_38_16;
	wire [WIDTH*2-1+1:0] tmp01_38_17;
	wire [WIDTH*2-1+1:0] tmp01_38_18;
	wire [WIDTH*2-1+1:0] tmp01_38_19;
	wire [WIDTH*2-1+1:0] tmp01_38_20;
	wire [WIDTH*2-1+1:0] tmp01_38_21;
	wire [WIDTH*2-1+1:0] tmp01_38_22;
	wire [WIDTH*2-1+1:0] tmp01_38_23;
	wire [WIDTH*2-1+1:0] tmp01_38_24;
	wire [WIDTH*2-1+1:0] tmp01_38_25;
	wire [WIDTH*2-1+1:0] tmp01_38_26;
	wire [WIDTH*2-1+1:0] tmp01_38_27;
	wire [WIDTH*2-1+1:0] tmp01_38_28;
	wire [WIDTH*2-1+1:0] tmp01_38_29;
	wire [WIDTH*2-1+1:0] tmp01_38_30;
	wire [WIDTH*2-1+1:0] tmp01_38_31;
	wire [WIDTH*2-1+1:0] tmp01_38_32;
	wire [WIDTH*2-1+1:0] tmp01_38_33;
	wire [WIDTH*2-1+1:0] tmp01_38_34;
	wire [WIDTH*2-1+1:0] tmp01_38_35;
	wire [WIDTH*2-1+1:0] tmp01_38_36;
	wire [WIDTH*2-1+1:0] tmp01_38_37;
	wire [WIDTH*2-1+1:0] tmp01_38_38;
	wire [WIDTH*2-1+1:0] tmp01_38_39;
	wire [WIDTH*2-1+1:0] tmp01_38_40;
	wire [WIDTH*2-1+1:0] tmp01_38_41;
	wire [WIDTH*2-1+1:0] tmp01_38_42;
	wire [WIDTH*2-1+1:0] tmp01_38_43;
	wire [WIDTH*2-1+1:0] tmp01_38_44;
	wire [WIDTH*2-1+1:0] tmp01_38_45;
	wire [WIDTH*2-1+1:0] tmp01_38_46;
	wire [WIDTH*2-1+1:0] tmp01_38_47;
	wire [WIDTH*2-1+1:0] tmp01_38_48;
	wire [WIDTH*2-1+1:0] tmp01_38_49;
	wire [WIDTH*2-1+1:0] tmp01_38_50;
	wire [WIDTH*2-1+1:0] tmp01_38_51;
	wire [WIDTH*2-1+1:0] tmp01_38_52;
	wire [WIDTH*2-1+1:0] tmp01_38_53;
	wire [WIDTH*2-1+1:0] tmp01_38_54;
	wire [WIDTH*2-1+1:0] tmp01_38_55;
	wire [WIDTH*2-1+1:0] tmp01_38_56;
	wire [WIDTH*2-1+1:0] tmp01_38_57;
	wire [WIDTH*2-1+1:0] tmp01_38_58;
	wire [WIDTH*2-1+1:0] tmp01_38_59;
	wire [WIDTH*2-1+1:0] tmp01_38_60;
	wire [WIDTH*2-1+1:0] tmp01_38_61;
	wire [WIDTH*2-1+1:0] tmp01_38_62;
	wire [WIDTH*2-1+1:0] tmp01_38_63;
	wire [WIDTH*2-1+1:0] tmp01_38_64;
	wire [WIDTH*2-1+1:0] tmp01_38_65;
	wire [WIDTH*2-1+1:0] tmp01_38_66;
	wire [WIDTH*2-1+1:0] tmp01_38_67;
	wire [WIDTH*2-1+1:0] tmp01_38_68;
	wire [WIDTH*2-1+1:0] tmp01_38_69;
	wire [WIDTH*2-1+1:0] tmp01_38_70;
	wire [WIDTH*2-1+1:0] tmp01_38_71;
	wire [WIDTH*2-1+1:0] tmp01_38_72;
	wire [WIDTH*2-1+1:0] tmp01_38_73;
	wire [WIDTH*2-1+1:0] tmp01_38_74;
	wire [WIDTH*2-1+1:0] tmp01_38_75;
	wire [WIDTH*2-1+1:0] tmp01_38_76;
	wire [WIDTH*2-1+1:0] tmp01_38_77;
	wire [WIDTH*2-1+1:0] tmp01_38_78;
	wire [WIDTH*2-1+1:0] tmp01_38_79;
	wire [WIDTH*2-1+1:0] tmp01_38_80;
	wire [WIDTH*2-1+1:0] tmp01_38_81;
	wire [WIDTH*2-1+1:0] tmp01_38_82;
	wire [WIDTH*2-1+1:0] tmp01_38_83;
	wire [WIDTH*2-1+1:0] tmp01_39_0;
	wire [WIDTH*2-1+1:0] tmp01_39_1;
	wire [WIDTH*2-1+1:0] tmp01_39_2;
	wire [WIDTH*2-1+1:0] tmp01_39_3;
	wire [WIDTH*2-1+1:0] tmp01_39_4;
	wire [WIDTH*2-1+1:0] tmp01_39_5;
	wire [WIDTH*2-1+1:0] tmp01_39_6;
	wire [WIDTH*2-1+1:0] tmp01_39_7;
	wire [WIDTH*2-1+1:0] tmp01_39_8;
	wire [WIDTH*2-1+1:0] tmp01_39_9;
	wire [WIDTH*2-1+1:0] tmp01_39_10;
	wire [WIDTH*2-1+1:0] tmp01_39_11;
	wire [WIDTH*2-1+1:0] tmp01_39_12;
	wire [WIDTH*2-1+1:0] tmp01_39_13;
	wire [WIDTH*2-1+1:0] tmp01_39_14;
	wire [WIDTH*2-1+1:0] tmp01_39_15;
	wire [WIDTH*2-1+1:0] tmp01_39_16;
	wire [WIDTH*2-1+1:0] tmp01_39_17;
	wire [WIDTH*2-1+1:0] tmp01_39_18;
	wire [WIDTH*2-1+1:0] tmp01_39_19;
	wire [WIDTH*2-1+1:0] tmp01_39_20;
	wire [WIDTH*2-1+1:0] tmp01_39_21;
	wire [WIDTH*2-1+1:0] tmp01_39_22;
	wire [WIDTH*2-1+1:0] tmp01_39_23;
	wire [WIDTH*2-1+1:0] tmp01_39_24;
	wire [WIDTH*2-1+1:0] tmp01_39_25;
	wire [WIDTH*2-1+1:0] tmp01_39_26;
	wire [WIDTH*2-1+1:0] tmp01_39_27;
	wire [WIDTH*2-1+1:0] tmp01_39_28;
	wire [WIDTH*2-1+1:0] tmp01_39_29;
	wire [WIDTH*2-1+1:0] tmp01_39_30;
	wire [WIDTH*2-1+1:0] tmp01_39_31;
	wire [WIDTH*2-1+1:0] tmp01_39_32;
	wire [WIDTH*2-1+1:0] tmp01_39_33;
	wire [WIDTH*2-1+1:0] tmp01_39_34;
	wire [WIDTH*2-1+1:0] tmp01_39_35;
	wire [WIDTH*2-1+1:0] tmp01_39_36;
	wire [WIDTH*2-1+1:0] tmp01_39_37;
	wire [WIDTH*2-1+1:0] tmp01_39_38;
	wire [WIDTH*2-1+1:0] tmp01_39_39;
	wire [WIDTH*2-1+1:0] tmp01_39_40;
	wire [WIDTH*2-1+1:0] tmp01_39_41;
	wire [WIDTH*2-1+1:0] tmp01_39_42;
	wire [WIDTH*2-1+1:0] tmp01_39_43;
	wire [WIDTH*2-1+1:0] tmp01_39_44;
	wire [WIDTH*2-1+1:0] tmp01_39_45;
	wire [WIDTH*2-1+1:0] tmp01_39_46;
	wire [WIDTH*2-1+1:0] tmp01_39_47;
	wire [WIDTH*2-1+1:0] tmp01_39_48;
	wire [WIDTH*2-1+1:0] tmp01_39_49;
	wire [WIDTH*2-1+1:0] tmp01_39_50;
	wire [WIDTH*2-1+1:0] tmp01_39_51;
	wire [WIDTH*2-1+1:0] tmp01_39_52;
	wire [WIDTH*2-1+1:0] tmp01_39_53;
	wire [WIDTH*2-1+1:0] tmp01_39_54;
	wire [WIDTH*2-1+1:0] tmp01_39_55;
	wire [WIDTH*2-1+1:0] tmp01_39_56;
	wire [WIDTH*2-1+1:0] tmp01_39_57;
	wire [WIDTH*2-1+1:0] tmp01_39_58;
	wire [WIDTH*2-1+1:0] tmp01_39_59;
	wire [WIDTH*2-1+1:0] tmp01_39_60;
	wire [WIDTH*2-1+1:0] tmp01_39_61;
	wire [WIDTH*2-1+1:0] tmp01_39_62;
	wire [WIDTH*2-1+1:0] tmp01_39_63;
	wire [WIDTH*2-1+1:0] tmp01_39_64;
	wire [WIDTH*2-1+1:0] tmp01_39_65;
	wire [WIDTH*2-1+1:0] tmp01_39_66;
	wire [WIDTH*2-1+1:0] tmp01_39_67;
	wire [WIDTH*2-1+1:0] tmp01_39_68;
	wire [WIDTH*2-1+1:0] tmp01_39_69;
	wire [WIDTH*2-1+1:0] tmp01_39_70;
	wire [WIDTH*2-1+1:0] tmp01_39_71;
	wire [WIDTH*2-1+1:0] tmp01_39_72;
	wire [WIDTH*2-1+1:0] tmp01_39_73;
	wire [WIDTH*2-1+1:0] tmp01_39_74;
	wire [WIDTH*2-1+1:0] tmp01_39_75;
	wire [WIDTH*2-1+1:0] tmp01_39_76;
	wire [WIDTH*2-1+1:0] tmp01_39_77;
	wire [WIDTH*2-1+1:0] tmp01_39_78;
	wire [WIDTH*2-1+1:0] tmp01_39_79;
	wire [WIDTH*2-1+1:0] tmp01_39_80;
	wire [WIDTH*2-1+1:0] tmp01_39_81;
	wire [WIDTH*2-1+1:0] tmp01_39_82;
	wire [WIDTH*2-1+1:0] tmp01_39_83;
	wire [WIDTH*2-1+1:0] tmp01_40_0;
	wire [WIDTH*2-1+1:0] tmp01_40_1;
	wire [WIDTH*2-1+1:0] tmp01_40_2;
	wire [WIDTH*2-1+1:0] tmp01_40_3;
	wire [WIDTH*2-1+1:0] tmp01_40_4;
	wire [WIDTH*2-1+1:0] tmp01_40_5;
	wire [WIDTH*2-1+1:0] tmp01_40_6;
	wire [WIDTH*2-1+1:0] tmp01_40_7;
	wire [WIDTH*2-1+1:0] tmp01_40_8;
	wire [WIDTH*2-1+1:0] tmp01_40_9;
	wire [WIDTH*2-1+1:0] tmp01_40_10;
	wire [WIDTH*2-1+1:0] tmp01_40_11;
	wire [WIDTH*2-1+1:0] tmp01_40_12;
	wire [WIDTH*2-1+1:0] tmp01_40_13;
	wire [WIDTH*2-1+1:0] tmp01_40_14;
	wire [WIDTH*2-1+1:0] tmp01_40_15;
	wire [WIDTH*2-1+1:0] tmp01_40_16;
	wire [WIDTH*2-1+1:0] tmp01_40_17;
	wire [WIDTH*2-1+1:0] tmp01_40_18;
	wire [WIDTH*2-1+1:0] tmp01_40_19;
	wire [WIDTH*2-1+1:0] tmp01_40_20;
	wire [WIDTH*2-1+1:0] tmp01_40_21;
	wire [WIDTH*2-1+1:0] tmp01_40_22;
	wire [WIDTH*2-1+1:0] tmp01_40_23;
	wire [WIDTH*2-1+1:0] tmp01_40_24;
	wire [WIDTH*2-1+1:0] tmp01_40_25;
	wire [WIDTH*2-1+1:0] tmp01_40_26;
	wire [WIDTH*2-1+1:0] tmp01_40_27;
	wire [WIDTH*2-1+1:0] tmp01_40_28;
	wire [WIDTH*2-1+1:0] tmp01_40_29;
	wire [WIDTH*2-1+1:0] tmp01_40_30;
	wire [WIDTH*2-1+1:0] tmp01_40_31;
	wire [WIDTH*2-1+1:0] tmp01_40_32;
	wire [WIDTH*2-1+1:0] tmp01_40_33;
	wire [WIDTH*2-1+1:0] tmp01_40_34;
	wire [WIDTH*2-1+1:0] tmp01_40_35;
	wire [WIDTH*2-1+1:0] tmp01_40_36;
	wire [WIDTH*2-1+1:0] tmp01_40_37;
	wire [WIDTH*2-1+1:0] tmp01_40_38;
	wire [WIDTH*2-1+1:0] tmp01_40_39;
	wire [WIDTH*2-1+1:0] tmp01_40_40;
	wire [WIDTH*2-1+1:0] tmp01_40_41;
	wire [WIDTH*2-1+1:0] tmp01_40_42;
	wire [WIDTH*2-1+1:0] tmp01_40_43;
	wire [WIDTH*2-1+1:0] tmp01_40_44;
	wire [WIDTH*2-1+1:0] tmp01_40_45;
	wire [WIDTH*2-1+1:0] tmp01_40_46;
	wire [WIDTH*2-1+1:0] tmp01_40_47;
	wire [WIDTH*2-1+1:0] tmp01_40_48;
	wire [WIDTH*2-1+1:0] tmp01_40_49;
	wire [WIDTH*2-1+1:0] tmp01_40_50;
	wire [WIDTH*2-1+1:0] tmp01_40_51;
	wire [WIDTH*2-1+1:0] tmp01_40_52;
	wire [WIDTH*2-1+1:0] tmp01_40_53;
	wire [WIDTH*2-1+1:0] tmp01_40_54;
	wire [WIDTH*2-1+1:0] tmp01_40_55;
	wire [WIDTH*2-1+1:0] tmp01_40_56;
	wire [WIDTH*2-1+1:0] tmp01_40_57;
	wire [WIDTH*2-1+1:0] tmp01_40_58;
	wire [WIDTH*2-1+1:0] tmp01_40_59;
	wire [WIDTH*2-1+1:0] tmp01_40_60;
	wire [WIDTH*2-1+1:0] tmp01_40_61;
	wire [WIDTH*2-1+1:0] tmp01_40_62;
	wire [WIDTH*2-1+1:0] tmp01_40_63;
	wire [WIDTH*2-1+1:0] tmp01_40_64;
	wire [WIDTH*2-1+1:0] tmp01_40_65;
	wire [WIDTH*2-1+1:0] tmp01_40_66;
	wire [WIDTH*2-1+1:0] tmp01_40_67;
	wire [WIDTH*2-1+1:0] tmp01_40_68;
	wire [WIDTH*2-1+1:0] tmp01_40_69;
	wire [WIDTH*2-1+1:0] tmp01_40_70;
	wire [WIDTH*2-1+1:0] tmp01_40_71;
	wire [WIDTH*2-1+1:0] tmp01_40_72;
	wire [WIDTH*2-1+1:0] tmp01_40_73;
	wire [WIDTH*2-1+1:0] tmp01_40_74;
	wire [WIDTH*2-1+1:0] tmp01_40_75;
	wire [WIDTH*2-1+1:0] tmp01_40_76;
	wire [WIDTH*2-1+1:0] tmp01_40_77;
	wire [WIDTH*2-1+1:0] tmp01_40_78;
	wire [WIDTH*2-1+1:0] tmp01_40_79;
	wire [WIDTH*2-1+1:0] tmp01_40_80;
	wire [WIDTH*2-1+1:0] tmp01_40_81;
	wire [WIDTH*2-1+1:0] tmp01_40_82;
	wire [WIDTH*2-1+1:0] tmp01_40_83;
	wire [WIDTH*2-1+1:0] tmp01_41_0;
	wire [WIDTH*2-1+1:0] tmp01_41_1;
	wire [WIDTH*2-1+1:0] tmp01_41_2;
	wire [WIDTH*2-1+1:0] tmp01_41_3;
	wire [WIDTH*2-1+1:0] tmp01_41_4;
	wire [WIDTH*2-1+1:0] tmp01_41_5;
	wire [WIDTH*2-1+1:0] tmp01_41_6;
	wire [WIDTH*2-1+1:0] tmp01_41_7;
	wire [WIDTH*2-1+1:0] tmp01_41_8;
	wire [WIDTH*2-1+1:0] tmp01_41_9;
	wire [WIDTH*2-1+1:0] tmp01_41_10;
	wire [WIDTH*2-1+1:0] tmp01_41_11;
	wire [WIDTH*2-1+1:0] tmp01_41_12;
	wire [WIDTH*2-1+1:0] tmp01_41_13;
	wire [WIDTH*2-1+1:0] tmp01_41_14;
	wire [WIDTH*2-1+1:0] tmp01_41_15;
	wire [WIDTH*2-1+1:0] tmp01_41_16;
	wire [WIDTH*2-1+1:0] tmp01_41_17;
	wire [WIDTH*2-1+1:0] tmp01_41_18;
	wire [WIDTH*2-1+1:0] tmp01_41_19;
	wire [WIDTH*2-1+1:0] tmp01_41_20;
	wire [WIDTH*2-1+1:0] tmp01_41_21;
	wire [WIDTH*2-1+1:0] tmp01_41_22;
	wire [WIDTH*2-1+1:0] tmp01_41_23;
	wire [WIDTH*2-1+1:0] tmp01_41_24;
	wire [WIDTH*2-1+1:0] tmp01_41_25;
	wire [WIDTH*2-1+1:0] tmp01_41_26;
	wire [WIDTH*2-1+1:0] tmp01_41_27;
	wire [WIDTH*2-1+1:0] tmp01_41_28;
	wire [WIDTH*2-1+1:0] tmp01_41_29;
	wire [WIDTH*2-1+1:0] tmp01_41_30;
	wire [WIDTH*2-1+1:0] tmp01_41_31;
	wire [WIDTH*2-1+1:0] tmp01_41_32;
	wire [WIDTH*2-1+1:0] tmp01_41_33;
	wire [WIDTH*2-1+1:0] tmp01_41_34;
	wire [WIDTH*2-1+1:0] tmp01_41_35;
	wire [WIDTH*2-1+1:0] tmp01_41_36;
	wire [WIDTH*2-1+1:0] tmp01_41_37;
	wire [WIDTH*2-1+1:0] tmp01_41_38;
	wire [WIDTH*2-1+1:0] tmp01_41_39;
	wire [WIDTH*2-1+1:0] tmp01_41_40;
	wire [WIDTH*2-1+1:0] tmp01_41_41;
	wire [WIDTH*2-1+1:0] tmp01_41_42;
	wire [WIDTH*2-1+1:0] tmp01_41_43;
	wire [WIDTH*2-1+1:0] tmp01_41_44;
	wire [WIDTH*2-1+1:0] tmp01_41_45;
	wire [WIDTH*2-1+1:0] tmp01_41_46;
	wire [WIDTH*2-1+1:0] tmp01_41_47;
	wire [WIDTH*2-1+1:0] tmp01_41_48;
	wire [WIDTH*2-1+1:0] tmp01_41_49;
	wire [WIDTH*2-1+1:0] tmp01_41_50;
	wire [WIDTH*2-1+1:0] tmp01_41_51;
	wire [WIDTH*2-1+1:0] tmp01_41_52;
	wire [WIDTH*2-1+1:0] tmp01_41_53;
	wire [WIDTH*2-1+1:0] tmp01_41_54;
	wire [WIDTH*2-1+1:0] tmp01_41_55;
	wire [WIDTH*2-1+1:0] tmp01_41_56;
	wire [WIDTH*2-1+1:0] tmp01_41_57;
	wire [WIDTH*2-1+1:0] tmp01_41_58;
	wire [WIDTH*2-1+1:0] tmp01_41_59;
	wire [WIDTH*2-1+1:0] tmp01_41_60;
	wire [WIDTH*2-1+1:0] tmp01_41_61;
	wire [WIDTH*2-1+1:0] tmp01_41_62;
	wire [WIDTH*2-1+1:0] tmp01_41_63;
	wire [WIDTH*2-1+1:0] tmp01_41_64;
	wire [WIDTH*2-1+1:0] tmp01_41_65;
	wire [WIDTH*2-1+1:0] tmp01_41_66;
	wire [WIDTH*2-1+1:0] tmp01_41_67;
	wire [WIDTH*2-1+1:0] tmp01_41_68;
	wire [WIDTH*2-1+1:0] tmp01_41_69;
	wire [WIDTH*2-1+1:0] tmp01_41_70;
	wire [WIDTH*2-1+1:0] tmp01_41_71;
	wire [WIDTH*2-1+1:0] tmp01_41_72;
	wire [WIDTH*2-1+1:0] tmp01_41_73;
	wire [WIDTH*2-1+1:0] tmp01_41_74;
	wire [WIDTH*2-1+1:0] tmp01_41_75;
	wire [WIDTH*2-1+1:0] tmp01_41_76;
	wire [WIDTH*2-1+1:0] tmp01_41_77;
	wire [WIDTH*2-1+1:0] tmp01_41_78;
	wire [WIDTH*2-1+1:0] tmp01_41_79;
	wire [WIDTH*2-1+1:0] tmp01_41_80;
	wire [WIDTH*2-1+1:0] tmp01_41_81;
	wire [WIDTH*2-1+1:0] tmp01_41_82;
	wire [WIDTH*2-1+1:0] tmp01_41_83;
	wire [WIDTH*2-1+1:0] tmp01_42_0;
	wire [WIDTH*2-1+1:0] tmp01_42_1;
	wire [WIDTH*2-1+1:0] tmp01_42_2;
	wire [WIDTH*2-1+1:0] tmp01_42_3;
	wire [WIDTH*2-1+1:0] tmp01_42_4;
	wire [WIDTH*2-1+1:0] tmp01_42_5;
	wire [WIDTH*2-1+1:0] tmp01_42_6;
	wire [WIDTH*2-1+1:0] tmp01_42_7;
	wire [WIDTH*2-1+1:0] tmp01_42_8;
	wire [WIDTH*2-1+1:0] tmp01_42_9;
	wire [WIDTH*2-1+1:0] tmp01_42_10;
	wire [WIDTH*2-1+1:0] tmp01_42_11;
	wire [WIDTH*2-1+1:0] tmp01_42_12;
	wire [WIDTH*2-1+1:0] tmp01_42_13;
	wire [WIDTH*2-1+1:0] tmp01_42_14;
	wire [WIDTH*2-1+1:0] tmp01_42_15;
	wire [WIDTH*2-1+1:0] tmp01_42_16;
	wire [WIDTH*2-1+1:0] tmp01_42_17;
	wire [WIDTH*2-1+1:0] tmp01_42_18;
	wire [WIDTH*2-1+1:0] tmp01_42_19;
	wire [WIDTH*2-1+1:0] tmp01_42_20;
	wire [WIDTH*2-1+1:0] tmp01_42_21;
	wire [WIDTH*2-1+1:0] tmp01_42_22;
	wire [WIDTH*2-1+1:0] tmp01_42_23;
	wire [WIDTH*2-1+1:0] tmp01_42_24;
	wire [WIDTH*2-1+1:0] tmp01_42_25;
	wire [WIDTH*2-1+1:0] tmp01_42_26;
	wire [WIDTH*2-1+1:0] tmp01_42_27;
	wire [WIDTH*2-1+1:0] tmp01_42_28;
	wire [WIDTH*2-1+1:0] tmp01_42_29;
	wire [WIDTH*2-1+1:0] tmp01_42_30;
	wire [WIDTH*2-1+1:0] tmp01_42_31;
	wire [WIDTH*2-1+1:0] tmp01_42_32;
	wire [WIDTH*2-1+1:0] tmp01_42_33;
	wire [WIDTH*2-1+1:0] tmp01_42_34;
	wire [WIDTH*2-1+1:0] tmp01_42_35;
	wire [WIDTH*2-1+1:0] tmp01_42_36;
	wire [WIDTH*2-1+1:0] tmp01_42_37;
	wire [WIDTH*2-1+1:0] tmp01_42_38;
	wire [WIDTH*2-1+1:0] tmp01_42_39;
	wire [WIDTH*2-1+1:0] tmp01_42_40;
	wire [WIDTH*2-1+1:0] tmp01_42_41;
	wire [WIDTH*2-1+1:0] tmp01_42_42;
	wire [WIDTH*2-1+1:0] tmp01_42_43;
	wire [WIDTH*2-1+1:0] tmp01_42_44;
	wire [WIDTH*2-1+1:0] tmp01_42_45;
	wire [WIDTH*2-1+1:0] tmp01_42_46;
	wire [WIDTH*2-1+1:0] tmp01_42_47;
	wire [WIDTH*2-1+1:0] tmp01_42_48;
	wire [WIDTH*2-1+1:0] tmp01_42_49;
	wire [WIDTH*2-1+1:0] tmp01_42_50;
	wire [WIDTH*2-1+1:0] tmp01_42_51;
	wire [WIDTH*2-1+1:0] tmp01_42_52;
	wire [WIDTH*2-1+1:0] tmp01_42_53;
	wire [WIDTH*2-1+1:0] tmp01_42_54;
	wire [WIDTH*2-1+1:0] tmp01_42_55;
	wire [WIDTH*2-1+1:0] tmp01_42_56;
	wire [WIDTH*2-1+1:0] tmp01_42_57;
	wire [WIDTH*2-1+1:0] tmp01_42_58;
	wire [WIDTH*2-1+1:0] tmp01_42_59;
	wire [WIDTH*2-1+1:0] tmp01_42_60;
	wire [WIDTH*2-1+1:0] tmp01_42_61;
	wire [WIDTH*2-1+1:0] tmp01_42_62;
	wire [WIDTH*2-1+1:0] tmp01_42_63;
	wire [WIDTH*2-1+1:0] tmp01_42_64;
	wire [WIDTH*2-1+1:0] tmp01_42_65;
	wire [WIDTH*2-1+1:0] tmp01_42_66;
	wire [WIDTH*2-1+1:0] tmp01_42_67;
	wire [WIDTH*2-1+1:0] tmp01_42_68;
	wire [WIDTH*2-1+1:0] tmp01_42_69;
	wire [WIDTH*2-1+1:0] tmp01_42_70;
	wire [WIDTH*2-1+1:0] tmp01_42_71;
	wire [WIDTH*2-1+1:0] tmp01_42_72;
	wire [WIDTH*2-1+1:0] tmp01_42_73;
	wire [WIDTH*2-1+1:0] tmp01_42_74;
	wire [WIDTH*2-1+1:0] tmp01_42_75;
	wire [WIDTH*2-1+1:0] tmp01_42_76;
	wire [WIDTH*2-1+1:0] tmp01_42_77;
	wire [WIDTH*2-1+1:0] tmp01_42_78;
	wire [WIDTH*2-1+1:0] tmp01_42_79;
	wire [WIDTH*2-1+1:0] tmp01_42_80;
	wire [WIDTH*2-1+1:0] tmp01_42_81;
	wire [WIDTH*2-1+1:0] tmp01_42_82;
	wire [WIDTH*2-1+1:0] tmp01_42_83;
	wire [WIDTH*2-1+1:0] tmp01_43_0;
	wire [WIDTH*2-1+1:0] tmp01_43_1;
	wire [WIDTH*2-1+1:0] tmp01_43_2;
	wire [WIDTH*2-1+1:0] tmp01_43_3;
	wire [WIDTH*2-1+1:0] tmp01_43_4;
	wire [WIDTH*2-1+1:0] tmp01_43_5;
	wire [WIDTH*2-1+1:0] tmp01_43_6;
	wire [WIDTH*2-1+1:0] tmp01_43_7;
	wire [WIDTH*2-1+1:0] tmp01_43_8;
	wire [WIDTH*2-1+1:0] tmp01_43_9;
	wire [WIDTH*2-1+1:0] tmp01_43_10;
	wire [WIDTH*2-1+1:0] tmp01_43_11;
	wire [WIDTH*2-1+1:0] tmp01_43_12;
	wire [WIDTH*2-1+1:0] tmp01_43_13;
	wire [WIDTH*2-1+1:0] tmp01_43_14;
	wire [WIDTH*2-1+1:0] tmp01_43_15;
	wire [WIDTH*2-1+1:0] tmp01_43_16;
	wire [WIDTH*2-1+1:0] tmp01_43_17;
	wire [WIDTH*2-1+1:0] tmp01_43_18;
	wire [WIDTH*2-1+1:0] tmp01_43_19;
	wire [WIDTH*2-1+1:0] tmp01_43_20;
	wire [WIDTH*2-1+1:0] tmp01_43_21;
	wire [WIDTH*2-1+1:0] tmp01_43_22;
	wire [WIDTH*2-1+1:0] tmp01_43_23;
	wire [WIDTH*2-1+1:0] tmp01_43_24;
	wire [WIDTH*2-1+1:0] tmp01_43_25;
	wire [WIDTH*2-1+1:0] tmp01_43_26;
	wire [WIDTH*2-1+1:0] tmp01_43_27;
	wire [WIDTH*2-1+1:0] tmp01_43_28;
	wire [WIDTH*2-1+1:0] tmp01_43_29;
	wire [WIDTH*2-1+1:0] tmp01_43_30;
	wire [WIDTH*2-1+1:0] tmp01_43_31;
	wire [WIDTH*2-1+1:0] tmp01_43_32;
	wire [WIDTH*2-1+1:0] tmp01_43_33;
	wire [WIDTH*2-1+1:0] tmp01_43_34;
	wire [WIDTH*2-1+1:0] tmp01_43_35;
	wire [WIDTH*2-1+1:0] tmp01_43_36;
	wire [WIDTH*2-1+1:0] tmp01_43_37;
	wire [WIDTH*2-1+1:0] tmp01_43_38;
	wire [WIDTH*2-1+1:0] tmp01_43_39;
	wire [WIDTH*2-1+1:0] tmp01_43_40;
	wire [WIDTH*2-1+1:0] tmp01_43_41;
	wire [WIDTH*2-1+1:0] tmp01_43_42;
	wire [WIDTH*2-1+1:0] tmp01_43_43;
	wire [WIDTH*2-1+1:0] tmp01_43_44;
	wire [WIDTH*2-1+1:0] tmp01_43_45;
	wire [WIDTH*2-1+1:0] tmp01_43_46;
	wire [WIDTH*2-1+1:0] tmp01_43_47;
	wire [WIDTH*2-1+1:0] tmp01_43_48;
	wire [WIDTH*2-1+1:0] tmp01_43_49;
	wire [WIDTH*2-1+1:0] tmp01_43_50;
	wire [WIDTH*2-1+1:0] tmp01_43_51;
	wire [WIDTH*2-1+1:0] tmp01_43_52;
	wire [WIDTH*2-1+1:0] tmp01_43_53;
	wire [WIDTH*2-1+1:0] tmp01_43_54;
	wire [WIDTH*2-1+1:0] tmp01_43_55;
	wire [WIDTH*2-1+1:0] tmp01_43_56;
	wire [WIDTH*2-1+1:0] tmp01_43_57;
	wire [WIDTH*2-1+1:0] tmp01_43_58;
	wire [WIDTH*2-1+1:0] tmp01_43_59;
	wire [WIDTH*2-1+1:0] tmp01_43_60;
	wire [WIDTH*2-1+1:0] tmp01_43_61;
	wire [WIDTH*2-1+1:0] tmp01_43_62;
	wire [WIDTH*2-1+1:0] tmp01_43_63;
	wire [WIDTH*2-1+1:0] tmp01_43_64;
	wire [WIDTH*2-1+1:0] tmp01_43_65;
	wire [WIDTH*2-1+1:0] tmp01_43_66;
	wire [WIDTH*2-1+1:0] tmp01_43_67;
	wire [WIDTH*2-1+1:0] tmp01_43_68;
	wire [WIDTH*2-1+1:0] tmp01_43_69;
	wire [WIDTH*2-1+1:0] tmp01_43_70;
	wire [WIDTH*2-1+1:0] tmp01_43_71;
	wire [WIDTH*2-1+1:0] tmp01_43_72;
	wire [WIDTH*2-1+1:0] tmp01_43_73;
	wire [WIDTH*2-1+1:0] tmp01_43_74;
	wire [WIDTH*2-1+1:0] tmp01_43_75;
	wire [WIDTH*2-1+1:0] tmp01_43_76;
	wire [WIDTH*2-1+1:0] tmp01_43_77;
	wire [WIDTH*2-1+1:0] tmp01_43_78;
	wire [WIDTH*2-1+1:0] tmp01_43_79;
	wire [WIDTH*2-1+1:0] tmp01_43_80;
	wire [WIDTH*2-1+1:0] tmp01_43_81;
	wire [WIDTH*2-1+1:0] tmp01_43_82;
	wire [WIDTH*2-1+1:0] tmp01_43_83;
	wire [WIDTH*2-1+1:0] tmp01_44_0;
	wire [WIDTH*2-1+1:0] tmp01_44_1;
	wire [WIDTH*2-1+1:0] tmp01_44_2;
	wire [WIDTH*2-1+1:0] tmp01_44_3;
	wire [WIDTH*2-1+1:0] tmp01_44_4;
	wire [WIDTH*2-1+1:0] tmp01_44_5;
	wire [WIDTH*2-1+1:0] tmp01_44_6;
	wire [WIDTH*2-1+1:0] tmp01_44_7;
	wire [WIDTH*2-1+1:0] tmp01_44_8;
	wire [WIDTH*2-1+1:0] tmp01_44_9;
	wire [WIDTH*2-1+1:0] tmp01_44_10;
	wire [WIDTH*2-1+1:0] tmp01_44_11;
	wire [WIDTH*2-1+1:0] tmp01_44_12;
	wire [WIDTH*2-1+1:0] tmp01_44_13;
	wire [WIDTH*2-1+1:0] tmp01_44_14;
	wire [WIDTH*2-1+1:0] tmp01_44_15;
	wire [WIDTH*2-1+1:0] tmp01_44_16;
	wire [WIDTH*2-1+1:0] tmp01_44_17;
	wire [WIDTH*2-1+1:0] tmp01_44_18;
	wire [WIDTH*2-1+1:0] tmp01_44_19;
	wire [WIDTH*2-1+1:0] tmp01_44_20;
	wire [WIDTH*2-1+1:0] tmp01_44_21;
	wire [WIDTH*2-1+1:0] tmp01_44_22;
	wire [WIDTH*2-1+1:0] tmp01_44_23;
	wire [WIDTH*2-1+1:0] tmp01_44_24;
	wire [WIDTH*2-1+1:0] tmp01_44_25;
	wire [WIDTH*2-1+1:0] tmp01_44_26;
	wire [WIDTH*2-1+1:0] tmp01_44_27;
	wire [WIDTH*2-1+1:0] tmp01_44_28;
	wire [WIDTH*2-1+1:0] tmp01_44_29;
	wire [WIDTH*2-1+1:0] tmp01_44_30;
	wire [WIDTH*2-1+1:0] tmp01_44_31;
	wire [WIDTH*2-1+1:0] tmp01_44_32;
	wire [WIDTH*2-1+1:0] tmp01_44_33;
	wire [WIDTH*2-1+1:0] tmp01_44_34;
	wire [WIDTH*2-1+1:0] tmp01_44_35;
	wire [WIDTH*2-1+1:0] tmp01_44_36;
	wire [WIDTH*2-1+1:0] tmp01_44_37;
	wire [WIDTH*2-1+1:0] tmp01_44_38;
	wire [WIDTH*2-1+1:0] tmp01_44_39;
	wire [WIDTH*2-1+1:0] tmp01_44_40;
	wire [WIDTH*2-1+1:0] tmp01_44_41;
	wire [WIDTH*2-1+1:0] tmp01_44_42;
	wire [WIDTH*2-1+1:0] tmp01_44_43;
	wire [WIDTH*2-1+1:0] tmp01_44_44;
	wire [WIDTH*2-1+1:0] tmp01_44_45;
	wire [WIDTH*2-1+1:0] tmp01_44_46;
	wire [WIDTH*2-1+1:0] tmp01_44_47;
	wire [WIDTH*2-1+1:0] tmp01_44_48;
	wire [WIDTH*2-1+1:0] tmp01_44_49;
	wire [WIDTH*2-1+1:0] tmp01_44_50;
	wire [WIDTH*2-1+1:0] tmp01_44_51;
	wire [WIDTH*2-1+1:0] tmp01_44_52;
	wire [WIDTH*2-1+1:0] tmp01_44_53;
	wire [WIDTH*2-1+1:0] tmp01_44_54;
	wire [WIDTH*2-1+1:0] tmp01_44_55;
	wire [WIDTH*2-1+1:0] tmp01_44_56;
	wire [WIDTH*2-1+1:0] tmp01_44_57;
	wire [WIDTH*2-1+1:0] tmp01_44_58;
	wire [WIDTH*2-1+1:0] tmp01_44_59;
	wire [WIDTH*2-1+1:0] tmp01_44_60;
	wire [WIDTH*2-1+1:0] tmp01_44_61;
	wire [WIDTH*2-1+1:0] tmp01_44_62;
	wire [WIDTH*2-1+1:0] tmp01_44_63;
	wire [WIDTH*2-1+1:0] tmp01_44_64;
	wire [WIDTH*2-1+1:0] tmp01_44_65;
	wire [WIDTH*2-1+1:0] tmp01_44_66;
	wire [WIDTH*2-1+1:0] tmp01_44_67;
	wire [WIDTH*2-1+1:0] tmp01_44_68;
	wire [WIDTH*2-1+1:0] tmp01_44_69;
	wire [WIDTH*2-1+1:0] tmp01_44_70;
	wire [WIDTH*2-1+1:0] tmp01_44_71;
	wire [WIDTH*2-1+1:0] tmp01_44_72;
	wire [WIDTH*2-1+1:0] tmp01_44_73;
	wire [WIDTH*2-1+1:0] tmp01_44_74;
	wire [WIDTH*2-1+1:0] tmp01_44_75;
	wire [WIDTH*2-1+1:0] tmp01_44_76;
	wire [WIDTH*2-1+1:0] tmp01_44_77;
	wire [WIDTH*2-1+1:0] tmp01_44_78;
	wire [WIDTH*2-1+1:0] tmp01_44_79;
	wire [WIDTH*2-1+1:0] tmp01_44_80;
	wire [WIDTH*2-1+1:0] tmp01_44_81;
	wire [WIDTH*2-1+1:0] tmp01_44_82;
	wire [WIDTH*2-1+1:0] tmp01_44_83;
	wire [WIDTH*2-1+1:0] tmp01_45_0;
	wire [WIDTH*2-1+1:0] tmp01_45_1;
	wire [WIDTH*2-1+1:0] tmp01_45_2;
	wire [WIDTH*2-1+1:0] tmp01_45_3;
	wire [WIDTH*2-1+1:0] tmp01_45_4;
	wire [WIDTH*2-1+1:0] tmp01_45_5;
	wire [WIDTH*2-1+1:0] tmp01_45_6;
	wire [WIDTH*2-1+1:0] tmp01_45_7;
	wire [WIDTH*2-1+1:0] tmp01_45_8;
	wire [WIDTH*2-1+1:0] tmp01_45_9;
	wire [WIDTH*2-1+1:0] tmp01_45_10;
	wire [WIDTH*2-1+1:0] tmp01_45_11;
	wire [WIDTH*2-1+1:0] tmp01_45_12;
	wire [WIDTH*2-1+1:0] tmp01_45_13;
	wire [WIDTH*2-1+1:0] tmp01_45_14;
	wire [WIDTH*2-1+1:0] tmp01_45_15;
	wire [WIDTH*2-1+1:0] tmp01_45_16;
	wire [WIDTH*2-1+1:0] tmp01_45_17;
	wire [WIDTH*2-1+1:0] tmp01_45_18;
	wire [WIDTH*2-1+1:0] tmp01_45_19;
	wire [WIDTH*2-1+1:0] tmp01_45_20;
	wire [WIDTH*2-1+1:0] tmp01_45_21;
	wire [WIDTH*2-1+1:0] tmp01_45_22;
	wire [WIDTH*2-1+1:0] tmp01_45_23;
	wire [WIDTH*2-1+1:0] tmp01_45_24;
	wire [WIDTH*2-1+1:0] tmp01_45_25;
	wire [WIDTH*2-1+1:0] tmp01_45_26;
	wire [WIDTH*2-1+1:0] tmp01_45_27;
	wire [WIDTH*2-1+1:0] tmp01_45_28;
	wire [WIDTH*2-1+1:0] tmp01_45_29;
	wire [WIDTH*2-1+1:0] tmp01_45_30;
	wire [WIDTH*2-1+1:0] tmp01_45_31;
	wire [WIDTH*2-1+1:0] tmp01_45_32;
	wire [WIDTH*2-1+1:0] tmp01_45_33;
	wire [WIDTH*2-1+1:0] tmp01_45_34;
	wire [WIDTH*2-1+1:0] tmp01_45_35;
	wire [WIDTH*2-1+1:0] tmp01_45_36;
	wire [WIDTH*2-1+1:0] tmp01_45_37;
	wire [WIDTH*2-1+1:0] tmp01_45_38;
	wire [WIDTH*2-1+1:0] tmp01_45_39;
	wire [WIDTH*2-1+1:0] tmp01_45_40;
	wire [WIDTH*2-1+1:0] tmp01_45_41;
	wire [WIDTH*2-1+1:0] tmp01_45_42;
	wire [WIDTH*2-1+1:0] tmp01_45_43;
	wire [WIDTH*2-1+1:0] tmp01_45_44;
	wire [WIDTH*2-1+1:0] tmp01_45_45;
	wire [WIDTH*2-1+1:0] tmp01_45_46;
	wire [WIDTH*2-1+1:0] tmp01_45_47;
	wire [WIDTH*2-1+1:0] tmp01_45_48;
	wire [WIDTH*2-1+1:0] tmp01_45_49;
	wire [WIDTH*2-1+1:0] tmp01_45_50;
	wire [WIDTH*2-1+1:0] tmp01_45_51;
	wire [WIDTH*2-1+1:0] tmp01_45_52;
	wire [WIDTH*2-1+1:0] tmp01_45_53;
	wire [WIDTH*2-1+1:0] tmp01_45_54;
	wire [WIDTH*2-1+1:0] tmp01_45_55;
	wire [WIDTH*2-1+1:0] tmp01_45_56;
	wire [WIDTH*2-1+1:0] tmp01_45_57;
	wire [WIDTH*2-1+1:0] tmp01_45_58;
	wire [WIDTH*2-1+1:0] tmp01_45_59;
	wire [WIDTH*2-1+1:0] tmp01_45_60;
	wire [WIDTH*2-1+1:0] tmp01_45_61;
	wire [WIDTH*2-1+1:0] tmp01_45_62;
	wire [WIDTH*2-1+1:0] tmp01_45_63;
	wire [WIDTH*2-1+1:0] tmp01_45_64;
	wire [WIDTH*2-1+1:0] tmp01_45_65;
	wire [WIDTH*2-1+1:0] tmp01_45_66;
	wire [WIDTH*2-1+1:0] tmp01_45_67;
	wire [WIDTH*2-1+1:0] tmp01_45_68;
	wire [WIDTH*2-1+1:0] tmp01_45_69;
	wire [WIDTH*2-1+1:0] tmp01_45_70;
	wire [WIDTH*2-1+1:0] tmp01_45_71;
	wire [WIDTH*2-1+1:0] tmp01_45_72;
	wire [WIDTH*2-1+1:0] tmp01_45_73;
	wire [WIDTH*2-1+1:0] tmp01_45_74;
	wire [WIDTH*2-1+1:0] tmp01_45_75;
	wire [WIDTH*2-1+1:0] tmp01_45_76;
	wire [WIDTH*2-1+1:0] tmp01_45_77;
	wire [WIDTH*2-1+1:0] tmp01_45_78;
	wire [WIDTH*2-1+1:0] tmp01_45_79;
	wire [WIDTH*2-1+1:0] tmp01_45_80;
	wire [WIDTH*2-1+1:0] tmp01_45_81;
	wire [WIDTH*2-1+1:0] tmp01_45_82;
	wire [WIDTH*2-1+1:0] tmp01_45_83;
	wire [WIDTH*2-1+1:0] tmp01_46_0;
	wire [WIDTH*2-1+1:0] tmp01_46_1;
	wire [WIDTH*2-1+1:0] tmp01_46_2;
	wire [WIDTH*2-1+1:0] tmp01_46_3;
	wire [WIDTH*2-1+1:0] tmp01_46_4;
	wire [WIDTH*2-1+1:0] tmp01_46_5;
	wire [WIDTH*2-1+1:0] tmp01_46_6;
	wire [WIDTH*2-1+1:0] tmp01_46_7;
	wire [WIDTH*2-1+1:0] tmp01_46_8;
	wire [WIDTH*2-1+1:0] tmp01_46_9;
	wire [WIDTH*2-1+1:0] tmp01_46_10;
	wire [WIDTH*2-1+1:0] tmp01_46_11;
	wire [WIDTH*2-1+1:0] tmp01_46_12;
	wire [WIDTH*2-1+1:0] tmp01_46_13;
	wire [WIDTH*2-1+1:0] tmp01_46_14;
	wire [WIDTH*2-1+1:0] tmp01_46_15;
	wire [WIDTH*2-1+1:0] tmp01_46_16;
	wire [WIDTH*2-1+1:0] tmp01_46_17;
	wire [WIDTH*2-1+1:0] tmp01_46_18;
	wire [WIDTH*2-1+1:0] tmp01_46_19;
	wire [WIDTH*2-1+1:0] tmp01_46_20;
	wire [WIDTH*2-1+1:0] tmp01_46_21;
	wire [WIDTH*2-1+1:0] tmp01_46_22;
	wire [WIDTH*2-1+1:0] tmp01_46_23;
	wire [WIDTH*2-1+1:0] tmp01_46_24;
	wire [WIDTH*2-1+1:0] tmp01_46_25;
	wire [WIDTH*2-1+1:0] tmp01_46_26;
	wire [WIDTH*2-1+1:0] tmp01_46_27;
	wire [WIDTH*2-1+1:0] tmp01_46_28;
	wire [WIDTH*2-1+1:0] tmp01_46_29;
	wire [WIDTH*2-1+1:0] tmp01_46_30;
	wire [WIDTH*2-1+1:0] tmp01_46_31;
	wire [WIDTH*2-1+1:0] tmp01_46_32;
	wire [WIDTH*2-1+1:0] tmp01_46_33;
	wire [WIDTH*2-1+1:0] tmp01_46_34;
	wire [WIDTH*2-1+1:0] tmp01_46_35;
	wire [WIDTH*2-1+1:0] tmp01_46_36;
	wire [WIDTH*2-1+1:0] tmp01_46_37;
	wire [WIDTH*2-1+1:0] tmp01_46_38;
	wire [WIDTH*2-1+1:0] tmp01_46_39;
	wire [WIDTH*2-1+1:0] tmp01_46_40;
	wire [WIDTH*2-1+1:0] tmp01_46_41;
	wire [WIDTH*2-1+1:0] tmp01_46_42;
	wire [WIDTH*2-1+1:0] tmp01_46_43;
	wire [WIDTH*2-1+1:0] tmp01_46_44;
	wire [WIDTH*2-1+1:0] tmp01_46_45;
	wire [WIDTH*2-1+1:0] tmp01_46_46;
	wire [WIDTH*2-1+1:0] tmp01_46_47;
	wire [WIDTH*2-1+1:0] tmp01_46_48;
	wire [WIDTH*2-1+1:0] tmp01_46_49;
	wire [WIDTH*2-1+1:0] tmp01_46_50;
	wire [WIDTH*2-1+1:0] tmp01_46_51;
	wire [WIDTH*2-1+1:0] tmp01_46_52;
	wire [WIDTH*2-1+1:0] tmp01_46_53;
	wire [WIDTH*2-1+1:0] tmp01_46_54;
	wire [WIDTH*2-1+1:0] tmp01_46_55;
	wire [WIDTH*2-1+1:0] tmp01_46_56;
	wire [WIDTH*2-1+1:0] tmp01_46_57;
	wire [WIDTH*2-1+1:0] tmp01_46_58;
	wire [WIDTH*2-1+1:0] tmp01_46_59;
	wire [WIDTH*2-1+1:0] tmp01_46_60;
	wire [WIDTH*2-1+1:0] tmp01_46_61;
	wire [WIDTH*2-1+1:0] tmp01_46_62;
	wire [WIDTH*2-1+1:0] tmp01_46_63;
	wire [WIDTH*2-1+1:0] tmp01_46_64;
	wire [WIDTH*2-1+1:0] tmp01_46_65;
	wire [WIDTH*2-1+1:0] tmp01_46_66;
	wire [WIDTH*2-1+1:0] tmp01_46_67;
	wire [WIDTH*2-1+1:0] tmp01_46_68;
	wire [WIDTH*2-1+1:0] tmp01_46_69;
	wire [WIDTH*2-1+1:0] tmp01_46_70;
	wire [WIDTH*2-1+1:0] tmp01_46_71;
	wire [WIDTH*2-1+1:0] tmp01_46_72;
	wire [WIDTH*2-1+1:0] tmp01_46_73;
	wire [WIDTH*2-1+1:0] tmp01_46_74;
	wire [WIDTH*2-1+1:0] tmp01_46_75;
	wire [WIDTH*2-1+1:0] tmp01_46_76;
	wire [WIDTH*2-1+1:0] tmp01_46_77;
	wire [WIDTH*2-1+1:0] tmp01_46_78;
	wire [WIDTH*2-1+1:0] tmp01_46_79;
	wire [WIDTH*2-1+1:0] tmp01_46_80;
	wire [WIDTH*2-1+1:0] tmp01_46_81;
	wire [WIDTH*2-1+1:0] tmp01_46_82;
	wire [WIDTH*2-1+1:0] tmp01_46_83;
	wire [WIDTH*2-1+1:0] tmp01_47_0;
	wire [WIDTH*2-1+1:0] tmp01_47_1;
	wire [WIDTH*2-1+1:0] tmp01_47_2;
	wire [WIDTH*2-1+1:0] tmp01_47_3;
	wire [WIDTH*2-1+1:0] tmp01_47_4;
	wire [WIDTH*2-1+1:0] tmp01_47_5;
	wire [WIDTH*2-1+1:0] tmp01_47_6;
	wire [WIDTH*2-1+1:0] tmp01_47_7;
	wire [WIDTH*2-1+1:0] tmp01_47_8;
	wire [WIDTH*2-1+1:0] tmp01_47_9;
	wire [WIDTH*2-1+1:0] tmp01_47_10;
	wire [WIDTH*2-1+1:0] tmp01_47_11;
	wire [WIDTH*2-1+1:0] tmp01_47_12;
	wire [WIDTH*2-1+1:0] tmp01_47_13;
	wire [WIDTH*2-1+1:0] tmp01_47_14;
	wire [WIDTH*2-1+1:0] tmp01_47_15;
	wire [WIDTH*2-1+1:0] tmp01_47_16;
	wire [WIDTH*2-1+1:0] tmp01_47_17;
	wire [WIDTH*2-1+1:0] tmp01_47_18;
	wire [WIDTH*2-1+1:0] tmp01_47_19;
	wire [WIDTH*2-1+1:0] tmp01_47_20;
	wire [WIDTH*2-1+1:0] tmp01_47_21;
	wire [WIDTH*2-1+1:0] tmp01_47_22;
	wire [WIDTH*2-1+1:0] tmp01_47_23;
	wire [WIDTH*2-1+1:0] tmp01_47_24;
	wire [WIDTH*2-1+1:0] tmp01_47_25;
	wire [WIDTH*2-1+1:0] tmp01_47_26;
	wire [WIDTH*2-1+1:0] tmp01_47_27;
	wire [WIDTH*2-1+1:0] tmp01_47_28;
	wire [WIDTH*2-1+1:0] tmp01_47_29;
	wire [WIDTH*2-1+1:0] tmp01_47_30;
	wire [WIDTH*2-1+1:0] tmp01_47_31;
	wire [WIDTH*2-1+1:0] tmp01_47_32;
	wire [WIDTH*2-1+1:0] tmp01_47_33;
	wire [WIDTH*2-1+1:0] tmp01_47_34;
	wire [WIDTH*2-1+1:0] tmp01_47_35;
	wire [WIDTH*2-1+1:0] tmp01_47_36;
	wire [WIDTH*2-1+1:0] tmp01_47_37;
	wire [WIDTH*2-1+1:0] tmp01_47_38;
	wire [WIDTH*2-1+1:0] tmp01_47_39;
	wire [WIDTH*2-1+1:0] tmp01_47_40;
	wire [WIDTH*2-1+1:0] tmp01_47_41;
	wire [WIDTH*2-1+1:0] tmp01_47_42;
	wire [WIDTH*2-1+1:0] tmp01_47_43;
	wire [WIDTH*2-1+1:0] tmp01_47_44;
	wire [WIDTH*2-1+1:0] tmp01_47_45;
	wire [WIDTH*2-1+1:0] tmp01_47_46;
	wire [WIDTH*2-1+1:0] tmp01_47_47;
	wire [WIDTH*2-1+1:0] tmp01_47_48;
	wire [WIDTH*2-1+1:0] tmp01_47_49;
	wire [WIDTH*2-1+1:0] tmp01_47_50;
	wire [WIDTH*2-1+1:0] tmp01_47_51;
	wire [WIDTH*2-1+1:0] tmp01_47_52;
	wire [WIDTH*2-1+1:0] tmp01_47_53;
	wire [WIDTH*2-1+1:0] tmp01_47_54;
	wire [WIDTH*2-1+1:0] tmp01_47_55;
	wire [WIDTH*2-1+1:0] tmp01_47_56;
	wire [WIDTH*2-1+1:0] tmp01_47_57;
	wire [WIDTH*2-1+1:0] tmp01_47_58;
	wire [WIDTH*2-1+1:0] tmp01_47_59;
	wire [WIDTH*2-1+1:0] tmp01_47_60;
	wire [WIDTH*2-1+1:0] tmp01_47_61;
	wire [WIDTH*2-1+1:0] tmp01_47_62;
	wire [WIDTH*2-1+1:0] tmp01_47_63;
	wire [WIDTH*2-1+1:0] tmp01_47_64;
	wire [WIDTH*2-1+1:0] tmp01_47_65;
	wire [WIDTH*2-1+1:0] tmp01_47_66;
	wire [WIDTH*2-1+1:0] tmp01_47_67;
	wire [WIDTH*2-1+1:0] tmp01_47_68;
	wire [WIDTH*2-1+1:0] tmp01_47_69;
	wire [WIDTH*2-1+1:0] tmp01_47_70;
	wire [WIDTH*2-1+1:0] tmp01_47_71;
	wire [WIDTH*2-1+1:0] tmp01_47_72;
	wire [WIDTH*2-1+1:0] tmp01_47_73;
	wire [WIDTH*2-1+1:0] tmp01_47_74;
	wire [WIDTH*2-1+1:0] tmp01_47_75;
	wire [WIDTH*2-1+1:0] tmp01_47_76;
	wire [WIDTH*2-1+1:0] tmp01_47_77;
	wire [WIDTH*2-1+1:0] tmp01_47_78;
	wire [WIDTH*2-1+1:0] tmp01_47_79;
	wire [WIDTH*2-1+1:0] tmp01_47_80;
	wire [WIDTH*2-1+1:0] tmp01_47_81;
	wire [WIDTH*2-1+1:0] tmp01_47_82;
	wire [WIDTH*2-1+1:0] tmp01_47_83;
	wire [WIDTH*2-1+1:0] tmp01_48_0;
	wire [WIDTH*2-1+1:0] tmp01_48_1;
	wire [WIDTH*2-1+1:0] tmp01_48_2;
	wire [WIDTH*2-1+1:0] tmp01_48_3;
	wire [WIDTH*2-1+1:0] tmp01_48_4;
	wire [WIDTH*2-1+1:0] tmp01_48_5;
	wire [WIDTH*2-1+1:0] tmp01_48_6;
	wire [WIDTH*2-1+1:0] tmp01_48_7;
	wire [WIDTH*2-1+1:0] tmp01_48_8;
	wire [WIDTH*2-1+1:0] tmp01_48_9;
	wire [WIDTH*2-1+1:0] tmp01_48_10;
	wire [WIDTH*2-1+1:0] tmp01_48_11;
	wire [WIDTH*2-1+1:0] tmp01_48_12;
	wire [WIDTH*2-1+1:0] tmp01_48_13;
	wire [WIDTH*2-1+1:0] tmp01_48_14;
	wire [WIDTH*2-1+1:0] tmp01_48_15;
	wire [WIDTH*2-1+1:0] tmp01_48_16;
	wire [WIDTH*2-1+1:0] tmp01_48_17;
	wire [WIDTH*2-1+1:0] tmp01_48_18;
	wire [WIDTH*2-1+1:0] tmp01_48_19;
	wire [WIDTH*2-1+1:0] tmp01_48_20;
	wire [WIDTH*2-1+1:0] tmp01_48_21;
	wire [WIDTH*2-1+1:0] tmp01_48_22;
	wire [WIDTH*2-1+1:0] tmp01_48_23;
	wire [WIDTH*2-1+1:0] tmp01_48_24;
	wire [WIDTH*2-1+1:0] tmp01_48_25;
	wire [WIDTH*2-1+1:0] tmp01_48_26;
	wire [WIDTH*2-1+1:0] tmp01_48_27;
	wire [WIDTH*2-1+1:0] tmp01_48_28;
	wire [WIDTH*2-1+1:0] tmp01_48_29;
	wire [WIDTH*2-1+1:0] tmp01_48_30;
	wire [WIDTH*2-1+1:0] tmp01_48_31;
	wire [WIDTH*2-1+1:0] tmp01_48_32;
	wire [WIDTH*2-1+1:0] tmp01_48_33;
	wire [WIDTH*2-1+1:0] tmp01_48_34;
	wire [WIDTH*2-1+1:0] tmp01_48_35;
	wire [WIDTH*2-1+1:0] tmp01_48_36;
	wire [WIDTH*2-1+1:0] tmp01_48_37;
	wire [WIDTH*2-1+1:0] tmp01_48_38;
	wire [WIDTH*2-1+1:0] tmp01_48_39;
	wire [WIDTH*2-1+1:0] tmp01_48_40;
	wire [WIDTH*2-1+1:0] tmp01_48_41;
	wire [WIDTH*2-1+1:0] tmp01_48_42;
	wire [WIDTH*2-1+1:0] tmp01_48_43;
	wire [WIDTH*2-1+1:0] tmp01_48_44;
	wire [WIDTH*2-1+1:0] tmp01_48_45;
	wire [WIDTH*2-1+1:0] tmp01_48_46;
	wire [WIDTH*2-1+1:0] tmp01_48_47;
	wire [WIDTH*2-1+1:0] tmp01_48_48;
	wire [WIDTH*2-1+1:0] tmp01_48_49;
	wire [WIDTH*2-1+1:0] tmp01_48_50;
	wire [WIDTH*2-1+1:0] tmp01_48_51;
	wire [WIDTH*2-1+1:0] tmp01_48_52;
	wire [WIDTH*2-1+1:0] tmp01_48_53;
	wire [WIDTH*2-1+1:0] tmp01_48_54;
	wire [WIDTH*2-1+1:0] tmp01_48_55;
	wire [WIDTH*2-1+1:0] tmp01_48_56;
	wire [WIDTH*2-1+1:0] tmp01_48_57;
	wire [WIDTH*2-1+1:0] tmp01_48_58;
	wire [WIDTH*2-1+1:0] tmp01_48_59;
	wire [WIDTH*2-1+1:0] tmp01_48_60;
	wire [WIDTH*2-1+1:0] tmp01_48_61;
	wire [WIDTH*2-1+1:0] tmp01_48_62;
	wire [WIDTH*2-1+1:0] tmp01_48_63;
	wire [WIDTH*2-1+1:0] tmp01_48_64;
	wire [WIDTH*2-1+1:0] tmp01_48_65;
	wire [WIDTH*2-1+1:0] tmp01_48_66;
	wire [WIDTH*2-1+1:0] tmp01_48_67;
	wire [WIDTH*2-1+1:0] tmp01_48_68;
	wire [WIDTH*2-1+1:0] tmp01_48_69;
	wire [WIDTH*2-1+1:0] tmp01_48_70;
	wire [WIDTH*2-1+1:0] tmp01_48_71;
	wire [WIDTH*2-1+1:0] tmp01_48_72;
	wire [WIDTH*2-1+1:0] tmp01_48_73;
	wire [WIDTH*2-1+1:0] tmp01_48_74;
	wire [WIDTH*2-1+1:0] tmp01_48_75;
	wire [WIDTH*2-1+1:0] tmp01_48_76;
	wire [WIDTH*2-1+1:0] tmp01_48_77;
	wire [WIDTH*2-1+1:0] tmp01_48_78;
	wire [WIDTH*2-1+1:0] tmp01_48_79;
	wire [WIDTH*2-1+1:0] tmp01_48_80;
	wire [WIDTH*2-1+1:0] tmp01_48_81;
	wire [WIDTH*2-1+1:0] tmp01_48_82;
	wire [WIDTH*2-1+1:0] tmp01_48_83;
	wire [WIDTH*2-1+1:0] tmp01_49_0;
	wire [WIDTH*2-1+1:0] tmp01_49_1;
	wire [WIDTH*2-1+1:0] tmp01_49_2;
	wire [WIDTH*2-1+1:0] tmp01_49_3;
	wire [WIDTH*2-1+1:0] tmp01_49_4;
	wire [WIDTH*2-1+1:0] tmp01_49_5;
	wire [WIDTH*2-1+1:0] tmp01_49_6;
	wire [WIDTH*2-1+1:0] tmp01_49_7;
	wire [WIDTH*2-1+1:0] tmp01_49_8;
	wire [WIDTH*2-1+1:0] tmp01_49_9;
	wire [WIDTH*2-1+1:0] tmp01_49_10;
	wire [WIDTH*2-1+1:0] tmp01_49_11;
	wire [WIDTH*2-1+1:0] tmp01_49_12;
	wire [WIDTH*2-1+1:0] tmp01_49_13;
	wire [WIDTH*2-1+1:0] tmp01_49_14;
	wire [WIDTH*2-1+1:0] tmp01_49_15;
	wire [WIDTH*2-1+1:0] tmp01_49_16;
	wire [WIDTH*2-1+1:0] tmp01_49_17;
	wire [WIDTH*2-1+1:0] tmp01_49_18;
	wire [WIDTH*2-1+1:0] tmp01_49_19;
	wire [WIDTH*2-1+1:0] tmp01_49_20;
	wire [WIDTH*2-1+1:0] tmp01_49_21;
	wire [WIDTH*2-1+1:0] tmp01_49_22;
	wire [WIDTH*2-1+1:0] tmp01_49_23;
	wire [WIDTH*2-1+1:0] tmp01_49_24;
	wire [WIDTH*2-1+1:0] tmp01_49_25;
	wire [WIDTH*2-1+1:0] tmp01_49_26;
	wire [WIDTH*2-1+1:0] tmp01_49_27;
	wire [WIDTH*2-1+1:0] tmp01_49_28;
	wire [WIDTH*2-1+1:0] tmp01_49_29;
	wire [WIDTH*2-1+1:0] tmp01_49_30;
	wire [WIDTH*2-1+1:0] tmp01_49_31;
	wire [WIDTH*2-1+1:0] tmp01_49_32;
	wire [WIDTH*2-1+1:0] tmp01_49_33;
	wire [WIDTH*2-1+1:0] tmp01_49_34;
	wire [WIDTH*2-1+1:0] tmp01_49_35;
	wire [WIDTH*2-1+1:0] tmp01_49_36;
	wire [WIDTH*2-1+1:0] tmp01_49_37;
	wire [WIDTH*2-1+1:0] tmp01_49_38;
	wire [WIDTH*2-1+1:0] tmp01_49_39;
	wire [WIDTH*2-1+1:0] tmp01_49_40;
	wire [WIDTH*2-1+1:0] tmp01_49_41;
	wire [WIDTH*2-1+1:0] tmp01_49_42;
	wire [WIDTH*2-1+1:0] tmp01_49_43;
	wire [WIDTH*2-1+1:0] tmp01_49_44;
	wire [WIDTH*2-1+1:0] tmp01_49_45;
	wire [WIDTH*2-1+1:0] tmp01_49_46;
	wire [WIDTH*2-1+1:0] tmp01_49_47;
	wire [WIDTH*2-1+1:0] tmp01_49_48;
	wire [WIDTH*2-1+1:0] tmp01_49_49;
	wire [WIDTH*2-1+1:0] tmp01_49_50;
	wire [WIDTH*2-1+1:0] tmp01_49_51;
	wire [WIDTH*2-1+1:0] tmp01_49_52;
	wire [WIDTH*2-1+1:0] tmp01_49_53;
	wire [WIDTH*2-1+1:0] tmp01_49_54;
	wire [WIDTH*2-1+1:0] tmp01_49_55;
	wire [WIDTH*2-1+1:0] tmp01_49_56;
	wire [WIDTH*2-1+1:0] tmp01_49_57;
	wire [WIDTH*2-1+1:0] tmp01_49_58;
	wire [WIDTH*2-1+1:0] tmp01_49_59;
	wire [WIDTH*2-1+1:0] tmp01_49_60;
	wire [WIDTH*2-1+1:0] tmp01_49_61;
	wire [WIDTH*2-1+1:0] tmp01_49_62;
	wire [WIDTH*2-1+1:0] tmp01_49_63;
	wire [WIDTH*2-1+1:0] tmp01_49_64;
	wire [WIDTH*2-1+1:0] tmp01_49_65;
	wire [WIDTH*2-1+1:0] tmp01_49_66;
	wire [WIDTH*2-1+1:0] tmp01_49_67;
	wire [WIDTH*2-1+1:0] tmp01_49_68;
	wire [WIDTH*2-1+1:0] tmp01_49_69;
	wire [WIDTH*2-1+1:0] tmp01_49_70;
	wire [WIDTH*2-1+1:0] tmp01_49_71;
	wire [WIDTH*2-1+1:0] tmp01_49_72;
	wire [WIDTH*2-1+1:0] tmp01_49_73;
	wire [WIDTH*2-1+1:0] tmp01_49_74;
	wire [WIDTH*2-1+1:0] tmp01_49_75;
	wire [WIDTH*2-1+1:0] tmp01_49_76;
	wire [WIDTH*2-1+1:0] tmp01_49_77;
	wire [WIDTH*2-1+1:0] tmp01_49_78;
	wire [WIDTH*2-1+1:0] tmp01_49_79;
	wire [WIDTH*2-1+1:0] tmp01_49_80;
	wire [WIDTH*2-1+1:0] tmp01_49_81;
	wire [WIDTH*2-1+1:0] tmp01_49_82;
	wire [WIDTH*2-1+1:0] tmp01_49_83;
	wire [WIDTH*2-1+1:0] tmp01_50_0;
	wire [WIDTH*2-1+1:0] tmp01_50_1;
	wire [WIDTH*2-1+1:0] tmp01_50_2;
	wire [WIDTH*2-1+1:0] tmp01_50_3;
	wire [WIDTH*2-1+1:0] tmp01_50_4;
	wire [WIDTH*2-1+1:0] tmp01_50_5;
	wire [WIDTH*2-1+1:0] tmp01_50_6;
	wire [WIDTH*2-1+1:0] tmp01_50_7;
	wire [WIDTH*2-1+1:0] tmp01_50_8;
	wire [WIDTH*2-1+1:0] tmp01_50_9;
	wire [WIDTH*2-1+1:0] tmp01_50_10;
	wire [WIDTH*2-1+1:0] tmp01_50_11;
	wire [WIDTH*2-1+1:0] tmp01_50_12;
	wire [WIDTH*2-1+1:0] tmp01_50_13;
	wire [WIDTH*2-1+1:0] tmp01_50_14;
	wire [WIDTH*2-1+1:0] tmp01_50_15;
	wire [WIDTH*2-1+1:0] tmp01_50_16;
	wire [WIDTH*2-1+1:0] tmp01_50_17;
	wire [WIDTH*2-1+1:0] tmp01_50_18;
	wire [WIDTH*2-1+1:0] tmp01_50_19;
	wire [WIDTH*2-1+1:0] tmp01_50_20;
	wire [WIDTH*2-1+1:0] tmp01_50_21;
	wire [WIDTH*2-1+1:0] tmp01_50_22;
	wire [WIDTH*2-1+1:0] tmp01_50_23;
	wire [WIDTH*2-1+1:0] tmp01_50_24;
	wire [WIDTH*2-1+1:0] tmp01_50_25;
	wire [WIDTH*2-1+1:0] tmp01_50_26;
	wire [WIDTH*2-1+1:0] tmp01_50_27;
	wire [WIDTH*2-1+1:0] tmp01_50_28;
	wire [WIDTH*2-1+1:0] tmp01_50_29;
	wire [WIDTH*2-1+1:0] tmp01_50_30;
	wire [WIDTH*2-1+1:0] tmp01_50_31;
	wire [WIDTH*2-1+1:0] tmp01_50_32;
	wire [WIDTH*2-1+1:0] tmp01_50_33;
	wire [WIDTH*2-1+1:0] tmp01_50_34;
	wire [WIDTH*2-1+1:0] tmp01_50_35;
	wire [WIDTH*2-1+1:0] tmp01_50_36;
	wire [WIDTH*2-1+1:0] tmp01_50_37;
	wire [WIDTH*2-1+1:0] tmp01_50_38;
	wire [WIDTH*2-1+1:0] tmp01_50_39;
	wire [WIDTH*2-1+1:0] tmp01_50_40;
	wire [WIDTH*2-1+1:0] tmp01_50_41;
	wire [WIDTH*2-1+1:0] tmp01_50_42;
	wire [WIDTH*2-1+1:0] tmp01_50_43;
	wire [WIDTH*2-1+1:0] tmp01_50_44;
	wire [WIDTH*2-1+1:0] tmp01_50_45;
	wire [WIDTH*2-1+1:0] tmp01_50_46;
	wire [WIDTH*2-1+1:0] tmp01_50_47;
	wire [WIDTH*2-1+1:0] tmp01_50_48;
	wire [WIDTH*2-1+1:0] tmp01_50_49;
	wire [WIDTH*2-1+1:0] tmp01_50_50;
	wire [WIDTH*2-1+1:0] tmp01_50_51;
	wire [WIDTH*2-1+1:0] tmp01_50_52;
	wire [WIDTH*2-1+1:0] tmp01_50_53;
	wire [WIDTH*2-1+1:0] tmp01_50_54;
	wire [WIDTH*2-1+1:0] tmp01_50_55;
	wire [WIDTH*2-1+1:0] tmp01_50_56;
	wire [WIDTH*2-1+1:0] tmp01_50_57;
	wire [WIDTH*2-1+1:0] tmp01_50_58;
	wire [WIDTH*2-1+1:0] tmp01_50_59;
	wire [WIDTH*2-1+1:0] tmp01_50_60;
	wire [WIDTH*2-1+1:0] tmp01_50_61;
	wire [WIDTH*2-1+1:0] tmp01_50_62;
	wire [WIDTH*2-1+1:0] tmp01_50_63;
	wire [WIDTH*2-1+1:0] tmp01_50_64;
	wire [WIDTH*2-1+1:0] tmp01_50_65;
	wire [WIDTH*2-1+1:0] tmp01_50_66;
	wire [WIDTH*2-1+1:0] tmp01_50_67;
	wire [WIDTH*2-1+1:0] tmp01_50_68;
	wire [WIDTH*2-1+1:0] tmp01_50_69;
	wire [WIDTH*2-1+1:0] tmp01_50_70;
	wire [WIDTH*2-1+1:0] tmp01_50_71;
	wire [WIDTH*2-1+1:0] tmp01_50_72;
	wire [WIDTH*2-1+1:0] tmp01_50_73;
	wire [WIDTH*2-1+1:0] tmp01_50_74;
	wire [WIDTH*2-1+1:0] tmp01_50_75;
	wire [WIDTH*2-1+1:0] tmp01_50_76;
	wire [WIDTH*2-1+1:0] tmp01_50_77;
	wire [WIDTH*2-1+1:0] tmp01_50_78;
	wire [WIDTH*2-1+1:0] tmp01_50_79;
	wire [WIDTH*2-1+1:0] tmp01_50_80;
	wire [WIDTH*2-1+1:0] tmp01_50_81;
	wire [WIDTH*2-1+1:0] tmp01_50_82;
	wire [WIDTH*2-1+1:0] tmp01_50_83;
	wire [WIDTH*2-1+1:0] tmp01_51_0;
	wire [WIDTH*2-1+1:0] tmp01_51_1;
	wire [WIDTH*2-1+1:0] tmp01_51_2;
	wire [WIDTH*2-1+1:0] tmp01_51_3;
	wire [WIDTH*2-1+1:0] tmp01_51_4;
	wire [WIDTH*2-1+1:0] tmp01_51_5;
	wire [WIDTH*2-1+1:0] tmp01_51_6;
	wire [WIDTH*2-1+1:0] tmp01_51_7;
	wire [WIDTH*2-1+1:0] tmp01_51_8;
	wire [WIDTH*2-1+1:0] tmp01_51_9;
	wire [WIDTH*2-1+1:0] tmp01_51_10;
	wire [WIDTH*2-1+1:0] tmp01_51_11;
	wire [WIDTH*2-1+1:0] tmp01_51_12;
	wire [WIDTH*2-1+1:0] tmp01_51_13;
	wire [WIDTH*2-1+1:0] tmp01_51_14;
	wire [WIDTH*2-1+1:0] tmp01_51_15;
	wire [WIDTH*2-1+1:0] tmp01_51_16;
	wire [WIDTH*2-1+1:0] tmp01_51_17;
	wire [WIDTH*2-1+1:0] tmp01_51_18;
	wire [WIDTH*2-1+1:0] tmp01_51_19;
	wire [WIDTH*2-1+1:0] tmp01_51_20;
	wire [WIDTH*2-1+1:0] tmp01_51_21;
	wire [WIDTH*2-1+1:0] tmp01_51_22;
	wire [WIDTH*2-1+1:0] tmp01_51_23;
	wire [WIDTH*2-1+1:0] tmp01_51_24;
	wire [WIDTH*2-1+1:0] tmp01_51_25;
	wire [WIDTH*2-1+1:0] tmp01_51_26;
	wire [WIDTH*2-1+1:0] tmp01_51_27;
	wire [WIDTH*2-1+1:0] tmp01_51_28;
	wire [WIDTH*2-1+1:0] tmp01_51_29;
	wire [WIDTH*2-1+1:0] tmp01_51_30;
	wire [WIDTH*2-1+1:0] tmp01_51_31;
	wire [WIDTH*2-1+1:0] tmp01_51_32;
	wire [WIDTH*2-1+1:0] tmp01_51_33;
	wire [WIDTH*2-1+1:0] tmp01_51_34;
	wire [WIDTH*2-1+1:0] tmp01_51_35;
	wire [WIDTH*2-1+1:0] tmp01_51_36;
	wire [WIDTH*2-1+1:0] tmp01_51_37;
	wire [WIDTH*2-1+1:0] tmp01_51_38;
	wire [WIDTH*2-1+1:0] tmp01_51_39;
	wire [WIDTH*2-1+1:0] tmp01_51_40;
	wire [WIDTH*2-1+1:0] tmp01_51_41;
	wire [WIDTH*2-1+1:0] tmp01_51_42;
	wire [WIDTH*2-1+1:0] tmp01_51_43;
	wire [WIDTH*2-1+1:0] tmp01_51_44;
	wire [WIDTH*2-1+1:0] tmp01_51_45;
	wire [WIDTH*2-1+1:0] tmp01_51_46;
	wire [WIDTH*2-1+1:0] tmp01_51_47;
	wire [WIDTH*2-1+1:0] tmp01_51_48;
	wire [WIDTH*2-1+1:0] tmp01_51_49;
	wire [WIDTH*2-1+1:0] tmp01_51_50;
	wire [WIDTH*2-1+1:0] tmp01_51_51;
	wire [WIDTH*2-1+1:0] tmp01_51_52;
	wire [WIDTH*2-1+1:0] tmp01_51_53;
	wire [WIDTH*2-1+1:0] tmp01_51_54;
	wire [WIDTH*2-1+1:0] tmp01_51_55;
	wire [WIDTH*2-1+1:0] tmp01_51_56;
	wire [WIDTH*2-1+1:0] tmp01_51_57;
	wire [WIDTH*2-1+1:0] tmp01_51_58;
	wire [WIDTH*2-1+1:0] tmp01_51_59;
	wire [WIDTH*2-1+1:0] tmp01_51_60;
	wire [WIDTH*2-1+1:0] tmp01_51_61;
	wire [WIDTH*2-1+1:0] tmp01_51_62;
	wire [WIDTH*2-1+1:0] tmp01_51_63;
	wire [WIDTH*2-1+1:0] tmp01_51_64;
	wire [WIDTH*2-1+1:0] tmp01_51_65;
	wire [WIDTH*2-1+1:0] tmp01_51_66;
	wire [WIDTH*2-1+1:0] tmp01_51_67;
	wire [WIDTH*2-1+1:0] tmp01_51_68;
	wire [WIDTH*2-1+1:0] tmp01_51_69;
	wire [WIDTH*2-1+1:0] tmp01_51_70;
	wire [WIDTH*2-1+1:0] tmp01_51_71;
	wire [WIDTH*2-1+1:0] tmp01_51_72;
	wire [WIDTH*2-1+1:0] tmp01_51_73;
	wire [WIDTH*2-1+1:0] tmp01_51_74;
	wire [WIDTH*2-1+1:0] tmp01_51_75;
	wire [WIDTH*2-1+1:0] tmp01_51_76;
	wire [WIDTH*2-1+1:0] tmp01_51_77;
	wire [WIDTH*2-1+1:0] tmp01_51_78;
	wire [WIDTH*2-1+1:0] tmp01_51_79;
	wire [WIDTH*2-1+1:0] tmp01_51_80;
	wire [WIDTH*2-1+1:0] tmp01_51_81;
	wire [WIDTH*2-1+1:0] tmp01_51_82;
	wire [WIDTH*2-1+1:0] tmp01_51_83;
	wire [WIDTH*2-1+1:0] tmp01_52_0;
	wire [WIDTH*2-1+1:0] tmp01_52_1;
	wire [WIDTH*2-1+1:0] tmp01_52_2;
	wire [WIDTH*2-1+1:0] tmp01_52_3;
	wire [WIDTH*2-1+1:0] tmp01_52_4;
	wire [WIDTH*2-1+1:0] tmp01_52_5;
	wire [WIDTH*2-1+1:0] tmp01_52_6;
	wire [WIDTH*2-1+1:0] tmp01_52_7;
	wire [WIDTH*2-1+1:0] tmp01_52_8;
	wire [WIDTH*2-1+1:0] tmp01_52_9;
	wire [WIDTH*2-1+1:0] tmp01_52_10;
	wire [WIDTH*2-1+1:0] tmp01_52_11;
	wire [WIDTH*2-1+1:0] tmp01_52_12;
	wire [WIDTH*2-1+1:0] tmp01_52_13;
	wire [WIDTH*2-1+1:0] tmp01_52_14;
	wire [WIDTH*2-1+1:0] tmp01_52_15;
	wire [WIDTH*2-1+1:0] tmp01_52_16;
	wire [WIDTH*2-1+1:0] tmp01_52_17;
	wire [WIDTH*2-1+1:0] tmp01_52_18;
	wire [WIDTH*2-1+1:0] tmp01_52_19;
	wire [WIDTH*2-1+1:0] tmp01_52_20;
	wire [WIDTH*2-1+1:0] tmp01_52_21;
	wire [WIDTH*2-1+1:0] tmp01_52_22;
	wire [WIDTH*2-1+1:0] tmp01_52_23;
	wire [WIDTH*2-1+1:0] tmp01_52_24;
	wire [WIDTH*2-1+1:0] tmp01_52_25;
	wire [WIDTH*2-1+1:0] tmp01_52_26;
	wire [WIDTH*2-1+1:0] tmp01_52_27;
	wire [WIDTH*2-1+1:0] tmp01_52_28;
	wire [WIDTH*2-1+1:0] tmp01_52_29;
	wire [WIDTH*2-1+1:0] tmp01_52_30;
	wire [WIDTH*2-1+1:0] tmp01_52_31;
	wire [WIDTH*2-1+1:0] tmp01_52_32;
	wire [WIDTH*2-1+1:0] tmp01_52_33;
	wire [WIDTH*2-1+1:0] tmp01_52_34;
	wire [WIDTH*2-1+1:0] tmp01_52_35;
	wire [WIDTH*2-1+1:0] tmp01_52_36;
	wire [WIDTH*2-1+1:0] tmp01_52_37;
	wire [WIDTH*2-1+1:0] tmp01_52_38;
	wire [WIDTH*2-1+1:0] tmp01_52_39;
	wire [WIDTH*2-1+1:0] tmp01_52_40;
	wire [WIDTH*2-1+1:0] tmp01_52_41;
	wire [WIDTH*2-1+1:0] tmp01_52_42;
	wire [WIDTH*2-1+1:0] tmp01_52_43;
	wire [WIDTH*2-1+1:0] tmp01_52_44;
	wire [WIDTH*2-1+1:0] tmp01_52_45;
	wire [WIDTH*2-1+1:0] tmp01_52_46;
	wire [WIDTH*2-1+1:0] tmp01_52_47;
	wire [WIDTH*2-1+1:0] tmp01_52_48;
	wire [WIDTH*2-1+1:0] tmp01_52_49;
	wire [WIDTH*2-1+1:0] tmp01_52_50;
	wire [WIDTH*2-1+1:0] tmp01_52_51;
	wire [WIDTH*2-1+1:0] tmp01_52_52;
	wire [WIDTH*2-1+1:0] tmp01_52_53;
	wire [WIDTH*2-1+1:0] tmp01_52_54;
	wire [WIDTH*2-1+1:0] tmp01_52_55;
	wire [WIDTH*2-1+1:0] tmp01_52_56;
	wire [WIDTH*2-1+1:0] tmp01_52_57;
	wire [WIDTH*2-1+1:0] tmp01_52_58;
	wire [WIDTH*2-1+1:0] tmp01_52_59;
	wire [WIDTH*2-1+1:0] tmp01_52_60;
	wire [WIDTH*2-1+1:0] tmp01_52_61;
	wire [WIDTH*2-1+1:0] tmp01_52_62;
	wire [WIDTH*2-1+1:0] tmp01_52_63;
	wire [WIDTH*2-1+1:0] tmp01_52_64;
	wire [WIDTH*2-1+1:0] tmp01_52_65;
	wire [WIDTH*2-1+1:0] tmp01_52_66;
	wire [WIDTH*2-1+1:0] tmp01_52_67;
	wire [WIDTH*2-1+1:0] tmp01_52_68;
	wire [WIDTH*2-1+1:0] tmp01_52_69;
	wire [WIDTH*2-1+1:0] tmp01_52_70;
	wire [WIDTH*2-1+1:0] tmp01_52_71;
	wire [WIDTH*2-1+1:0] tmp01_52_72;
	wire [WIDTH*2-1+1:0] tmp01_52_73;
	wire [WIDTH*2-1+1:0] tmp01_52_74;
	wire [WIDTH*2-1+1:0] tmp01_52_75;
	wire [WIDTH*2-1+1:0] tmp01_52_76;
	wire [WIDTH*2-1+1:0] tmp01_52_77;
	wire [WIDTH*2-1+1:0] tmp01_52_78;
	wire [WIDTH*2-1+1:0] tmp01_52_79;
	wire [WIDTH*2-1+1:0] tmp01_52_80;
	wire [WIDTH*2-1+1:0] tmp01_52_81;
	wire [WIDTH*2-1+1:0] tmp01_52_82;
	wire [WIDTH*2-1+1:0] tmp01_52_83;
	wire [WIDTH*2-1+1:0] tmp01_53_0;
	wire [WIDTH*2-1+1:0] tmp01_53_1;
	wire [WIDTH*2-1+1:0] tmp01_53_2;
	wire [WIDTH*2-1+1:0] tmp01_53_3;
	wire [WIDTH*2-1+1:0] tmp01_53_4;
	wire [WIDTH*2-1+1:0] tmp01_53_5;
	wire [WIDTH*2-1+1:0] tmp01_53_6;
	wire [WIDTH*2-1+1:0] tmp01_53_7;
	wire [WIDTH*2-1+1:0] tmp01_53_8;
	wire [WIDTH*2-1+1:0] tmp01_53_9;
	wire [WIDTH*2-1+1:0] tmp01_53_10;
	wire [WIDTH*2-1+1:0] tmp01_53_11;
	wire [WIDTH*2-1+1:0] tmp01_53_12;
	wire [WIDTH*2-1+1:0] tmp01_53_13;
	wire [WIDTH*2-1+1:0] tmp01_53_14;
	wire [WIDTH*2-1+1:0] tmp01_53_15;
	wire [WIDTH*2-1+1:0] tmp01_53_16;
	wire [WIDTH*2-1+1:0] tmp01_53_17;
	wire [WIDTH*2-1+1:0] tmp01_53_18;
	wire [WIDTH*2-1+1:0] tmp01_53_19;
	wire [WIDTH*2-1+1:0] tmp01_53_20;
	wire [WIDTH*2-1+1:0] tmp01_53_21;
	wire [WIDTH*2-1+1:0] tmp01_53_22;
	wire [WIDTH*2-1+1:0] tmp01_53_23;
	wire [WIDTH*2-1+1:0] tmp01_53_24;
	wire [WIDTH*2-1+1:0] tmp01_53_25;
	wire [WIDTH*2-1+1:0] tmp01_53_26;
	wire [WIDTH*2-1+1:0] tmp01_53_27;
	wire [WIDTH*2-1+1:0] tmp01_53_28;
	wire [WIDTH*2-1+1:0] tmp01_53_29;
	wire [WIDTH*2-1+1:0] tmp01_53_30;
	wire [WIDTH*2-1+1:0] tmp01_53_31;
	wire [WIDTH*2-1+1:0] tmp01_53_32;
	wire [WIDTH*2-1+1:0] tmp01_53_33;
	wire [WIDTH*2-1+1:0] tmp01_53_34;
	wire [WIDTH*2-1+1:0] tmp01_53_35;
	wire [WIDTH*2-1+1:0] tmp01_53_36;
	wire [WIDTH*2-1+1:0] tmp01_53_37;
	wire [WIDTH*2-1+1:0] tmp01_53_38;
	wire [WIDTH*2-1+1:0] tmp01_53_39;
	wire [WIDTH*2-1+1:0] tmp01_53_40;
	wire [WIDTH*2-1+1:0] tmp01_53_41;
	wire [WIDTH*2-1+1:0] tmp01_53_42;
	wire [WIDTH*2-1+1:0] tmp01_53_43;
	wire [WIDTH*2-1+1:0] tmp01_53_44;
	wire [WIDTH*2-1+1:0] tmp01_53_45;
	wire [WIDTH*2-1+1:0] tmp01_53_46;
	wire [WIDTH*2-1+1:0] tmp01_53_47;
	wire [WIDTH*2-1+1:0] tmp01_53_48;
	wire [WIDTH*2-1+1:0] tmp01_53_49;
	wire [WIDTH*2-1+1:0] tmp01_53_50;
	wire [WIDTH*2-1+1:0] tmp01_53_51;
	wire [WIDTH*2-1+1:0] tmp01_53_52;
	wire [WIDTH*2-1+1:0] tmp01_53_53;
	wire [WIDTH*2-1+1:0] tmp01_53_54;
	wire [WIDTH*2-1+1:0] tmp01_53_55;
	wire [WIDTH*2-1+1:0] tmp01_53_56;
	wire [WIDTH*2-1+1:0] tmp01_53_57;
	wire [WIDTH*2-1+1:0] tmp01_53_58;
	wire [WIDTH*2-1+1:0] tmp01_53_59;
	wire [WIDTH*2-1+1:0] tmp01_53_60;
	wire [WIDTH*2-1+1:0] tmp01_53_61;
	wire [WIDTH*2-1+1:0] tmp01_53_62;
	wire [WIDTH*2-1+1:0] tmp01_53_63;
	wire [WIDTH*2-1+1:0] tmp01_53_64;
	wire [WIDTH*2-1+1:0] tmp01_53_65;
	wire [WIDTH*2-1+1:0] tmp01_53_66;
	wire [WIDTH*2-1+1:0] tmp01_53_67;
	wire [WIDTH*2-1+1:0] tmp01_53_68;
	wire [WIDTH*2-1+1:0] tmp01_53_69;
	wire [WIDTH*2-1+1:0] tmp01_53_70;
	wire [WIDTH*2-1+1:0] tmp01_53_71;
	wire [WIDTH*2-1+1:0] tmp01_53_72;
	wire [WIDTH*2-1+1:0] tmp01_53_73;
	wire [WIDTH*2-1+1:0] tmp01_53_74;
	wire [WIDTH*2-1+1:0] tmp01_53_75;
	wire [WIDTH*2-1+1:0] tmp01_53_76;
	wire [WIDTH*2-1+1:0] tmp01_53_77;
	wire [WIDTH*2-1+1:0] tmp01_53_78;
	wire [WIDTH*2-1+1:0] tmp01_53_79;
	wire [WIDTH*2-1+1:0] tmp01_53_80;
	wire [WIDTH*2-1+1:0] tmp01_53_81;
	wire [WIDTH*2-1+1:0] tmp01_53_82;
	wire [WIDTH*2-1+1:0] tmp01_53_83;
	wire [WIDTH*2-1+1:0] tmp01_54_0;
	wire [WIDTH*2-1+1:0] tmp01_54_1;
	wire [WIDTH*2-1+1:0] tmp01_54_2;
	wire [WIDTH*2-1+1:0] tmp01_54_3;
	wire [WIDTH*2-1+1:0] tmp01_54_4;
	wire [WIDTH*2-1+1:0] tmp01_54_5;
	wire [WIDTH*2-1+1:0] tmp01_54_6;
	wire [WIDTH*2-1+1:0] tmp01_54_7;
	wire [WIDTH*2-1+1:0] tmp01_54_8;
	wire [WIDTH*2-1+1:0] tmp01_54_9;
	wire [WIDTH*2-1+1:0] tmp01_54_10;
	wire [WIDTH*2-1+1:0] tmp01_54_11;
	wire [WIDTH*2-1+1:0] tmp01_54_12;
	wire [WIDTH*2-1+1:0] tmp01_54_13;
	wire [WIDTH*2-1+1:0] tmp01_54_14;
	wire [WIDTH*2-1+1:0] tmp01_54_15;
	wire [WIDTH*2-1+1:0] tmp01_54_16;
	wire [WIDTH*2-1+1:0] tmp01_54_17;
	wire [WIDTH*2-1+1:0] tmp01_54_18;
	wire [WIDTH*2-1+1:0] tmp01_54_19;
	wire [WIDTH*2-1+1:0] tmp01_54_20;
	wire [WIDTH*2-1+1:0] tmp01_54_21;
	wire [WIDTH*2-1+1:0] tmp01_54_22;
	wire [WIDTH*2-1+1:0] tmp01_54_23;
	wire [WIDTH*2-1+1:0] tmp01_54_24;
	wire [WIDTH*2-1+1:0] tmp01_54_25;
	wire [WIDTH*2-1+1:0] tmp01_54_26;
	wire [WIDTH*2-1+1:0] tmp01_54_27;
	wire [WIDTH*2-1+1:0] tmp01_54_28;
	wire [WIDTH*2-1+1:0] tmp01_54_29;
	wire [WIDTH*2-1+1:0] tmp01_54_30;
	wire [WIDTH*2-1+1:0] tmp01_54_31;
	wire [WIDTH*2-1+1:0] tmp01_54_32;
	wire [WIDTH*2-1+1:0] tmp01_54_33;
	wire [WIDTH*2-1+1:0] tmp01_54_34;
	wire [WIDTH*2-1+1:0] tmp01_54_35;
	wire [WIDTH*2-1+1:0] tmp01_54_36;
	wire [WIDTH*2-1+1:0] tmp01_54_37;
	wire [WIDTH*2-1+1:0] tmp01_54_38;
	wire [WIDTH*2-1+1:0] tmp01_54_39;
	wire [WIDTH*2-1+1:0] tmp01_54_40;
	wire [WIDTH*2-1+1:0] tmp01_54_41;
	wire [WIDTH*2-1+1:0] tmp01_54_42;
	wire [WIDTH*2-1+1:0] tmp01_54_43;
	wire [WIDTH*2-1+1:0] tmp01_54_44;
	wire [WIDTH*2-1+1:0] tmp01_54_45;
	wire [WIDTH*2-1+1:0] tmp01_54_46;
	wire [WIDTH*2-1+1:0] tmp01_54_47;
	wire [WIDTH*2-1+1:0] tmp01_54_48;
	wire [WIDTH*2-1+1:0] tmp01_54_49;
	wire [WIDTH*2-1+1:0] tmp01_54_50;
	wire [WIDTH*2-1+1:0] tmp01_54_51;
	wire [WIDTH*2-1+1:0] tmp01_54_52;
	wire [WIDTH*2-1+1:0] tmp01_54_53;
	wire [WIDTH*2-1+1:0] tmp01_54_54;
	wire [WIDTH*2-1+1:0] tmp01_54_55;
	wire [WIDTH*2-1+1:0] tmp01_54_56;
	wire [WIDTH*2-1+1:0] tmp01_54_57;
	wire [WIDTH*2-1+1:0] tmp01_54_58;
	wire [WIDTH*2-1+1:0] tmp01_54_59;
	wire [WIDTH*2-1+1:0] tmp01_54_60;
	wire [WIDTH*2-1+1:0] tmp01_54_61;
	wire [WIDTH*2-1+1:0] tmp01_54_62;
	wire [WIDTH*2-1+1:0] tmp01_54_63;
	wire [WIDTH*2-1+1:0] tmp01_54_64;
	wire [WIDTH*2-1+1:0] tmp01_54_65;
	wire [WIDTH*2-1+1:0] tmp01_54_66;
	wire [WIDTH*2-1+1:0] tmp01_54_67;
	wire [WIDTH*2-1+1:0] tmp01_54_68;
	wire [WIDTH*2-1+1:0] tmp01_54_69;
	wire [WIDTH*2-1+1:0] tmp01_54_70;
	wire [WIDTH*2-1+1:0] tmp01_54_71;
	wire [WIDTH*2-1+1:0] tmp01_54_72;
	wire [WIDTH*2-1+1:0] tmp01_54_73;
	wire [WIDTH*2-1+1:0] tmp01_54_74;
	wire [WIDTH*2-1+1:0] tmp01_54_75;
	wire [WIDTH*2-1+1:0] tmp01_54_76;
	wire [WIDTH*2-1+1:0] tmp01_54_77;
	wire [WIDTH*2-1+1:0] tmp01_54_78;
	wire [WIDTH*2-1+1:0] tmp01_54_79;
	wire [WIDTH*2-1+1:0] tmp01_54_80;
	wire [WIDTH*2-1+1:0] tmp01_54_81;
	wire [WIDTH*2-1+1:0] tmp01_54_82;
	wire [WIDTH*2-1+1:0] tmp01_54_83;
	wire [WIDTH*2-1+1:0] tmp01_55_0;
	wire [WIDTH*2-1+1:0] tmp01_55_1;
	wire [WIDTH*2-1+1:0] tmp01_55_2;
	wire [WIDTH*2-1+1:0] tmp01_55_3;
	wire [WIDTH*2-1+1:0] tmp01_55_4;
	wire [WIDTH*2-1+1:0] tmp01_55_5;
	wire [WIDTH*2-1+1:0] tmp01_55_6;
	wire [WIDTH*2-1+1:0] tmp01_55_7;
	wire [WIDTH*2-1+1:0] tmp01_55_8;
	wire [WIDTH*2-1+1:0] tmp01_55_9;
	wire [WIDTH*2-1+1:0] tmp01_55_10;
	wire [WIDTH*2-1+1:0] tmp01_55_11;
	wire [WIDTH*2-1+1:0] tmp01_55_12;
	wire [WIDTH*2-1+1:0] tmp01_55_13;
	wire [WIDTH*2-1+1:0] tmp01_55_14;
	wire [WIDTH*2-1+1:0] tmp01_55_15;
	wire [WIDTH*2-1+1:0] tmp01_55_16;
	wire [WIDTH*2-1+1:0] tmp01_55_17;
	wire [WIDTH*2-1+1:0] tmp01_55_18;
	wire [WIDTH*2-1+1:0] tmp01_55_19;
	wire [WIDTH*2-1+1:0] tmp01_55_20;
	wire [WIDTH*2-1+1:0] tmp01_55_21;
	wire [WIDTH*2-1+1:0] tmp01_55_22;
	wire [WIDTH*2-1+1:0] tmp01_55_23;
	wire [WIDTH*2-1+1:0] tmp01_55_24;
	wire [WIDTH*2-1+1:0] tmp01_55_25;
	wire [WIDTH*2-1+1:0] tmp01_55_26;
	wire [WIDTH*2-1+1:0] tmp01_55_27;
	wire [WIDTH*2-1+1:0] tmp01_55_28;
	wire [WIDTH*2-1+1:0] tmp01_55_29;
	wire [WIDTH*2-1+1:0] tmp01_55_30;
	wire [WIDTH*2-1+1:0] tmp01_55_31;
	wire [WIDTH*2-1+1:0] tmp01_55_32;
	wire [WIDTH*2-1+1:0] tmp01_55_33;
	wire [WIDTH*2-1+1:0] tmp01_55_34;
	wire [WIDTH*2-1+1:0] tmp01_55_35;
	wire [WIDTH*2-1+1:0] tmp01_55_36;
	wire [WIDTH*2-1+1:0] tmp01_55_37;
	wire [WIDTH*2-1+1:0] tmp01_55_38;
	wire [WIDTH*2-1+1:0] tmp01_55_39;
	wire [WIDTH*2-1+1:0] tmp01_55_40;
	wire [WIDTH*2-1+1:0] tmp01_55_41;
	wire [WIDTH*2-1+1:0] tmp01_55_42;
	wire [WIDTH*2-1+1:0] tmp01_55_43;
	wire [WIDTH*2-1+1:0] tmp01_55_44;
	wire [WIDTH*2-1+1:0] tmp01_55_45;
	wire [WIDTH*2-1+1:0] tmp01_55_46;
	wire [WIDTH*2-1+1:0] tmp01_55_47;
	wire [WIDTH*2-1+1:0] tmp01_55_48;
	wire [WIDTH*2-1+1:0] tmp01_55_49;
	wire [WIDTH*2-1+1:0] tmp01_55_50;
	wire [WIDTH*2-1+1:0] tmp01_55_51;
	wire [WIDTH*2-1+1:0] tmp01_55_52;
	wire [WIDTH*2-1+1:0] tmp01_55_53;
	wire [WIDTH*2-1+1:0] tmp01_55_54;
	wire [WIDTH*2-1+1:0] tmp01_55_55;
	wire [WIDTH*2-1+1:0] tmp01_55_56;
	wire [WIDTH*2-1+1:0] tmp01_55_57;
	wire [WIDTH*2-1+1:0] tmp01_55_58;
	wire [WIDTH*2-1+1:0] tmp01_55_59;
	wire [WIDTH*2-1+1:0] tmp01_55_60;
	wire [WIDTH*2-1+1:0] tmp01_55_61;
	wire [WIDTH*2-1+1:0] tmp01_55_62;
	wire [WIDTH*2-1+1:0] tmp01_55_63;
	wire [WIDTH*2-1+1:0] tmp01_55_64;
	wire [WIDTH*2-1+1:0] tmp01_55_65;
	wire [WIDTH*2-1+1:0] tmp01_55_66;
	wire [WIDTH*2-1+1:0] tmp01_55_67;
	wire [WIDTH*2-1+1:0] tmp01_55_68;
	wire [WIDTH*2-1+1:0] tmp01_55_69;
	wire [WIDTH*2-1+1:0] tmp01_55_70;
	wire [WIDTH*2-1+1:0] tmp01_55_71;
	wire [WIDTH*2-1+1:0] tmp01_55_72;
	wire [WIDTH*2-1+1:0] tmp01_55_73;
	wire [WIDTH*2-1+1:0] tmp01_55_74;
	wire [WIDTH*2-1+1:0] tmp01_55_75;
	wire [WIDTH*2-1+1:0] tmp01_55_76;
	wire [WIDTH*2-1+1:0] tmp01_55_77;
	wire [WIDTH*2-1+1:0] tmp01_55_78;
	wire [WIDTH*2-1+1:0] tmp01_55_79;
	wire [WIDTH*2-1+1:0] tmp01_55_80;
	wire [WIDTH*2-1+1:0] tmp01_55_81;
	wire [WIDTH*2-1+1:0] tmp01_55_82;
	wire [WIDTH*2-1+1:0] tmp01_55_83;
	wire [WIDTH*2-1+1:0] tmp01_56_0;
	wire [WIDTH*2-1+1:0] tmp01_56_1;
	wire [WIDTH*2-1+1:0] tmp01_56_2;
	wire [WIDTH*2-1+1:0] tmp01_56_3;
	wire [WIDTH*2-1+1:0] tmp01_56_4;
	wire [WIDTH*2-1+1:0] tmp01_56_5;
	wire [WIDTH*2-1+1:0] tmp01_56_6;
	wire [WIDTH*2-1+1:0] tmp01_56_7;
	wire [WIDTH*2-1+1:0] tmp01_56_8;
	wire [WIDTH*2-1+1:0] tmp01_56_9;
	wire [WIDTH*2-1+1:0] tmp01_56_10;
	wire [WIDTH*2-1+1:0] tmp01_56_11;
	wire [WIDTH*2-1+1:0] tmp01_56_12;
	wire [WIDTH*2-1+1:0] tmp01_56_13;
	wire [WIDTH*2-1+1:0] tmp01_56_14;
	wire [WIDTH*2-1+1:0] tmp01_56_15;
	wire [WIDTH*2-1+1:0] tmp01_56_16;
	wire [WIDTH*2-1+1:0] tmp01_56_17;
	wire [WIDTH*2-1+1:0] tmp01_56_18;
	wire [WIDTH*2-1+1:0] tmp01_56_19;
	wire [WIDTH*2-1+1:0] tmp01_56_20;
	wire [WIDTH*2-1+1:0] tmp01_56_21;
	wire [WIDTH*2-1+1:0] tmp01_56_22;
	wire [WIDTH*2-1+1:0] tmp01_56_23;
	wire [WIDTH*2-1+1:0] tmp01_56_24;
	wire [WIDTH*2-1+1:0] tmp01_56_25;
	wire [WIDTH*2-1+1:0] tmp01_56_26;
	wire [WIDTH*2-1+1:0] tmp01_56_27;
	wire [WIDTH*2-1+1:0] tmp01_56_28;
	wire [WIDTH*2-1+1:0] tmp01_56_29;
	wire [WIDTH*2-1+1:0] tmp01_56_30;
	wire [WIDTH*2-1+1:0] tmp01_56_31;
	wire [WIDTH*2-1+1:0] tmp01_56_32;
	wire [WIDTH*2-1+1:0] tmp01_56_33;
	wire [WIDTH*2-1+1:0] tmp01_56_34;
	wire [WIDTH*2-1+1:0] tmp01_56_35;
	wire [WIDTH*2-1+1:0] tmp01_56_36;
	wire [WIDTH*2-1+1:0] tmp01_56_37;
	wire [WIDTH*2-1+1:0] tmp01_56_38;
	wire [WIDTH*2-1+1:0] tmp01_56_39;
	wire [WIDTH*2-1+1:0] tmp01_56_40;
	wire [WIDTH*2-1+1:0] tmp01_56_41;
	wire [WIDTH*2-1+1:0] tmp01_56_42;
	wire [WIDTH*2-1+1:0] tmp01_56_43;
	wire [WIDTH*2-1+1:0] tmp01_56_44;
	wire [WIDTH*2-1+1:0] tmp01_56_45;
	wire [WIDTH*2-1+1:0] tmp01_56_46;
	wire [WIDTH*2-1+1:0] tmp01_56_47;
	wire [WIDTH*2-1+1:0] tmp01_56_48;
	wire [WIDTH*2-1+1:0] tmp01_56_49;
	wire [WIDTH*2-1+1:0] tmp01_56_50;
	wire [WIDTH*2-1+1:0] tmp01_56_51;
	wire [WIDTH*2-1+1:0] tmp01_56_52;
	wire [WIDTH*2-1+1:0] tmp01_56_53;
	wire [WIDTH*2-1+1:0] tmp01_56_54;
	wire [WIDTH*2-1+1:0] tmp01_56_55;
	wire [WIDTH*2-1+1:0] tmp01_56_56;
	wire [WIDTH*2-1+1:0] tmp01_56_57;
	wire [WIDTH*2-1+1:0] tmp01_56_58;
	wire [WIDTH*2-1+1:0] tmp01_56_59;
	wire [WIDTH*2-1+1:0] tmp01_56_60;
	wire [WIDTH*2-1+1:0] tmp01_56_61;
	wire [WIDTH*2-1+1:0] tmp01_56_62;
	wire [WIDTH*2-1+1:0] tmp01_56_63;
	wire [WIDTH*2-1+1:0] tmp01_56_64;
	wire [WIDTH*2-1+1:0] tmp01_56_65;
	wire [WIDTH*2-1+1:0] tmp01_56_66;
	wire [WIDTH*2-1+1:0] tmp01_56_67;
	wire [WIDTH*2-1+1:0] tmp01_56_68;
	wire [WIDTH*2-1+1:0] tmp01_56_69;
	wire [WIDTH*2-1+1:0] tmp01_56_70;
	wire [WIDTH*2-1+1:0] tmp01_56_71;
	wire [WIDTH*2-1+1:0] tmp01_56_72;
	wire [WIDTH*2-1+1:0] tmp01_56_73;
	wire [WIDTH*2-1+1:0] tmp01_56_74;
	wire [WIDTH*2-1+1:0] tmp01_56_75;
	wire [WIDTH*2-1+1:0] tmp01_56_76;
	wire [WIDTH*2-1+1:0] tmp01_56_77;
	wire [WIDTH*2-1+1:0] tmp01_56_78;
	wire [WIDTH*2-1+1:0] tmp01_56_79;
	wire [WIDTH*2-1+1:0] tmp01_56_80;
	wire [WIDTH*2-1+1:0] tmp01_56_81;
	wire [WIDTH*2-1+1:0] tmp01_56_82;
	wire [WIDTH*2-1+1:0] tmp01_56_83;
	wire [WIDTH*2-1+1:0] tmp01_57_0;
	wire [WIDTH*2-1+1:0] tmp01_57_1;
	wire [WIDTH*2-1+1:0] tmp01_57_2;
	wire [WIDTH*2-1+1:0] tmp01_57_3;
	wire [WIDTH*2-1+1:0] tmp01_57_4;
	wire [WIDTH*2-1+1:0] tmp01_57_5;
	wire [WIDTH*2-1+1:0] tmp01_57_6;
	wire [WIDTH*2-1+1:0] tmp01_57_7;
	wire [WIDTH*2-1+1:0] tmp01_57_8;
	wire [WIDTH*2-1+1:0] tmp01_57_9;
	wire [WIDTH*2-1+1:0] tmp01_57_10;
	wire [WIDTH*2-1+1:0] tmp01_57_11;
	wire [WIDTH*2-1+1:0] tmp01_57_12;
	wire [WIDTH*2-1+1:0] tmp01_57_13;
	wire [WIDTH*2-1+1:0] tmp01_57_14;
	wire [WIDTH*2-1+1:0] tmp01_57_15;
	wire [WIDTH*2-1+1:0] tmp01_57_16;
	wire [WIDTH*2-1+1:0] tmp01_57_17;
	wire [WIDTH*2-1+1:0] tmp01_57_18;
	wire [WIDTH*2-1+1:0] tmp01_57_19;
	wire [WIDTH*2-1+1:0] tmp01_57_20;
	wire [WIDTH*2-1+1:0] tmp01_57_21;
	wire [WIDTH*2-1+1:0] tmp01_57_22;
	wire [WIDTH*2-1+1:0] tmp01_57_23;
	wire [WIDTH*2-1+1:0] tmp01_57_24;
	wire [WIDTH*2-1+1:0] tmp01_57_25;
	wire [WIDTH*2-1+1:0] tmp01_57_26;
	wire [WIDTH*2-1+1:0] tmp01_57_27;
	wire [WIDTH*2-1+1:0] tmp01_57_28;
	wire [WIDTH*2-1+1:0] tmp01_57_29;
	wire [WIDTH*2-1+1:0] tmp01_57_30;
	wire [WIDTH*2-1+1:0] tmp01_57_31;
	wire [WIDTH*2-1+1:0] tmp01_57_32;
	wire [WIDTH*2-1+1:0] tmp01_57_33;
	wire [WIDTH*2-1+1:0] tmp01_57_34;
	wire [WIDTH*2-1+1:0] tmp01_57_35;
	wire [WIDTH*2-1+1:0] tmp01_57_36;
	wire [WIDTH*2-1+1:0] tmp01_57_37;
	wire [WIDTH*2-1+1:0] tmp01_57_38;
	wire [WIDTH*2-1+1:0] tmp01_57_39;
	wire [WIDTH*2-1+1:0] tmp01_57_40;
	wire [WIDTH*2-1+1:0] tmp01_57_41;
	wire [WIDTH*2-1+1:0] tmp01_57_42;
	wire [WIDTH*2-1+1:0] tmp01_57_43;
	wire [WIDTH*2-1+1:0] tmp01_57_44;
	wire [WIDTH*2-1+1:0] tmp01_57_45;
	wire [WIDTH*2-1+1:0] tmp01_57_46;
	wire [WIDTH*2-1+1:0] tmp01_57_47;
	wire [WIDTH*2-1+1:0] tmp01_57_48;
	wire [WIDTH*2-1+1:0] tmp01_57_49;
	wire [WIDTH*2-1+1:0] tmp01_57_50;
	wire [WIDTH*2-1+1:0] tmp01_57_51;
	wire [WIDTH*2-1+1:0] tmp01_57_52;
	wire [WIDTH*2-1+1:0] tmp01_57_53;
	wire [WIDTH*2-1+1:0] tmp01_57_54;
	wire [WIDTH*2-1+1:0] tmp01_57_55;
	wire [WIDTH*2-1+1:0] tmp01_57_56;
	wire [WIDTH*2-1+1:0] tmp01_57_57;
	wire [WIDTH*2-1+1:0] tmp01_57_58;
	wire [WIDTH*2-1+1:0] tmp01_57_59;
	wire [WIDTH*2-1+1:0] tmp01_57_60;
	wire [WIDTH*2-1+1:0] tmp01_57_61;
	wire [WIDTH*2-1+1:0] tmp01_57_62;
	wire [WIDTH*2-1+1:0] tmp01_57_63;
	wire [WIDTH*2-1+1:0] tmp01_57_64;
	wire [WIDTH*2-1+1:0] tmp01_57_65;
	wire [WIDTH*2-1+1:0] tmp01_57_66;
	wire [WIDTH*2-1+1:0] tmp01_57_67;
	wire [WIDTH*2-1+1:0] tmp01_57_68;
	wire [WIDTH*2-1+1:0] tmp01_57_69;
	wire [WIDTH*2-1+1:0] tmp01_57_70;
	wire [WIDTH*2-1+1:0] tmp01_57_71;
	wire [WIDTH*2-1+1:0] tmp01_57_72;
	wire [WIDTH*2-1+1:0] tmp01_57_73;
	wire [WIDTH*2-1+1:0] tmp01_57_74;
	wire [WIDTH*2-1+1:0] tmp01_57_75;
	wire [WIDTH*2-1+1:0] tmp01_57_76;
	wire [WIDTH*2-1+1:0] tmp01_57_77;
	wire [WIDTH*2-1+1:0] tmp01_57_78;
	wire [WIDTH*2-1+1:0] tmp01_57_79;
	wire [WIDTH*2-1+1:0] tmp01_57_80;
	wire [WIDTH*2-1+1:0] tmp01_57_81;
	wire [WIDTH*2-1+1:0] tmp01_57_82;
	wire [WIDTH*2-1+1:0] tmp01_57_83;
	wire [WIDTH*2-1+1:0] tmp01_58_0;
	wire [WIDTH*2-1+1:0] tmp01_58_1;
	wire [WIDTH*2-1+1:0] tmp01_58_2;
	wire [WIDTH*2-1+1:0] tmp01_58_3;
	wire [WIDTH*2-1+1:0] tmp01_58_4;
	wire [WIDTH*2-1+1:0] tmp01_58_5;
	wire [WIDTH*2-1+1:0] tmp01_58_6;
	wire [WIDTH*2-1+1:0] tmp01_58_7;
	wire [WIDTH*2-1+1:0] tmp01_58_8;
	wire [WIDTH*2-1+1:0] tmp01_58_9;
	wire [WIDTH*2-1+1:0] tmp01_58_10;
	wire [WIDTH*2-1+1:0] tmp01_58_11;
	wire [WIDTH*2-1+1:0] tmp01_58_12;
	wire [WIDTH*2-1+1:0] tmp01_58_13;
	wire [WIDTH*2-1+1:0] tmp01_58_14;
	wire [WIDTH*2-1+1:0] tmp01_58_15;
	wire [WIDTH*2-1+1:0] tmp01_58_16;
	wire [WIDTH*2-1+1:0] tmp01_58_17;
	wire [WIDTH*2-1+1:0] tmp01_58_18;
	wire [WIDTH*2-1+1:0] tmp01_58_19;
	wire [WIDTH*2-1+1:0] tmp01_58_20;
	wire [WIDTH*2-1+1:0] tmp01_58_21;
	wire [WIDTH*2-1+1:0] tmp01_58_22;
	wire [WIDTH*2-1+1:0] tmp01_58_23;
	wire [WIDTH*2-1+1:0] tmp01_58_24;
	wire [WIDTH*2-1+1:0] tmp01_58_25;
	wire [WIDTH*2-1+1:0] tmp01_58_26;
	wire [WIDTH*2-1+1:0] tmp01_58_27;
	wire [WIDTH*2-1+1:0] tmp01_58_28;
	wire [WIDTH*2-1+1:0] tmp01_58_29;
	wire [WIDTH*2-1+1:0] tmp01_58_30;
	wire [WIDTH*2-1+1:0] tmp01_58_31;
	wire [WIDTH*2-1+1:0] tmp01_58_32;
	wire [WIDTH*2-1+1:0] tmp01_58_33;
	wire [WIDTH*2-1+1:0] tmp01_58_34;
	wire [WIDTH*2-1+1:0] tmp01_58_35;
	wire [WIDTH*2-1+1:0] tmp01_58_36;
	wire [WIDTH*2-1+1:0] tmp01_58_37;
	wire [WIDTH*2-1+1:0] tmp01_58_38;
	wire [WIDTH*2-1+1:0] tmp01_58_39;
	wire [WIDTH*2-1+1:0] tmp01_58_40;
	wire [WIDTH*2-1+1:0] tmp01_58_41;
	wire [WIDTH*2-1+1:0] tmp01_58_42;
	wire [WIDTH*2-1+1:0] tmp01_58_43;
	wire [WIDTH*2-1+1:0] tmp01_58_44;
	wire [WIDTH*2-1+1:0] tmp01_58_45;
	wire [WIDTH*2-1+1:0] tmp01_58_46;
	wire [WIDTH*2-1+1:0] tmp01_58_47;
	wire [WIDTH*2-1+1:0] tmp01_58_48;
	wire [WIDTH*2-1+1:0] tmp01_58_49;
	wire [WIDTH*2-1+1:0] tmp01_58_50;
	wire [WIDTH*2-1+1:0] tmp01_58_51;
	wire [WIDTH*2-1+1:0] tmp01_58_52;
	wire [WIDTH*2-1+1:0] tmp01_58_53;
	wire [WIDTH*2-1+1:0] tmp01_58_54;
	wire [WIDTH*2-1+1:0] tmp01_58_55;
	wire [WIDTH*2-1+1:0] tmp01_58_56;
	wire [WIDTH*2-1+1:0] tmp01_58_57;
	wire [WIDTH*2-1+1:0] tmp01_58_58;
	wire [WIDTH*2-1+1:0] tmp01_58_59;
	wire [WIDTH*2-1+1:0] tmp01_58_60;
	wire [WIDTH*2-1+1:0] tmp01_58_61;
	wire [WIDTH*2-1+1:0] tmp01_58_62;
	wire [WIDTH*2-1+1:0] tmp01_58_63;
	wire [WIDTH*2-1+1:0] tmp01_58_64;
	wire [WIDTH*2-1+1:0] tmp01_58_65;
	wire [WIDTH*2-1+1:0] tmp01_58_66;
	wire [WIDTH*2-1+1:0] tmp01_58_67;
	wire [WIDTH*2-1+1:0] tmp01_58_68;
	wire [WIDTH*2-1+1:0] tmp01_58_69;
	wire [WIDTH*2-1+1:0] tmp01_58_70;
	wire [WIDTH*2-1+1:0] tmp01_58_71;
	wire [WIDTH*2-1+1:0] tmp01_58_72;
	wire [WIDTH*2-1+1:0] tmp01_58_73;
	wire [WIDTH*2-1+1:0] tmp01_58_74;
	wire [WIDTH*2-1+1:0] tmp01_58_75;
	wire [WIDTH*2-1+1:0] tmp01_58_76;
	wire [WIDTH*2-1+1:0] tmp01_58_77;
	wire [WIDTH*2-1+1:0] tmp01_58_78;
	wire [WIDTH*2-1+1:0] tmp01_58_79;
	wire [WIDTH*2-1+1:0] tmp01_58_80;
	wire [WIDTH*2-1+1:0] tmp01_58_81;
	wire [WIDTH*2-1+1:0] tmp01_58_82;
	wire [WIDTH*2-1+1:0] tmp01_58_83;
	wire [WIDTH*2-1+1:0] tmp01_59_0;
	wire [WIDTH*2-1+1:0] tmp01_59_1;
	wire [WIDTH*2-1+1:0] tmp01_59_2;
	wire [WIDTH*2-1+1:0] tmp01_59_3;
	wire [WIDTH*2-1+1:0] tmp01_59_4;
	wire [WIDTH*2-1+1:0] tmp01_59_5;
	wire [WIDTH*2-1+1:0] tmp01_59_6;
	wire [WIDTH*2-1+1:0] tmp01_59_7;
	wire [WIDTH*2-1+1:0] tmp01_59_8;
	wire [WIDTH*2-1+1:0] tmp01_59_9;
	wire [WIDTH*2-1+1:0] tmp01_59_10;
	wire [WIDTH*2-1+1:0] tmp01_59_11;
	wire [WIDTH*2-1+1:0] tmp01_59_12;
	wire [WIDTH*2-1+1:0] tmp01_59_13;
	wire [WIDTH*2-1+1:0] tmp01_59_14;
	wire [WIDTH*2-1+1:0] tmp01_59_15;
	wire [WIDTH*2-1+1:0] tmp01_59_16;
	wire [WIDTH*2-1+1:0] tmp01_59_17;
	wire [WIDTH*2-1+1:0] tmp01_59_18;
	wire [WIDTH*2-1+1:0] tmp01_59_19;
	wire [WIDTH*2-1+1:0] tmp01_59_20;
	wire [WIDTH*2-1+1:0] tmp01_59_21;
	wire [WIDTH*2-1+1:0] tmp01_59_22;
	wire [WIDTH*2-1+1:0] tmp01_59_23;
	wire [WIDTH*2-1+1:0] tmp01_59_24;
	wire [WIDTH*2-1+1:0] tmp01_59_25;
	wire [WIDTH*2-1+1:0] tmp01_59_26;
	wire [WIDTH*2-1+1:0] tmp01_59_27;
	wire [WIDTH*2-1+1:0] tmp01_59_28;
	wire [WIDTH*2-1+1:0] tmp01_59_29;
	wire [WIDTH*2-1+1:0] tmp01_59_30;
	wire [WIDTH*2-1+1:0] tmp01_59_31;
	wire [WIDTH*2-1+1:0] tmp01_59_32;
	wire [WIDTH*2-1+1:0] tmp01_59_33;
	wire [WIDTH*2-1+1:0] tmp01_59_34;
	wire [WIDTH*2-1+1:0] tmp01_59_35;
	wire [WIDTH*2-1+1:0] tmp01_59_36;
	wire [WIDTH*2-1+1:0] tmp01_59_37;
	wire [WIDTH*2-1+1:0] tmp01_59_38;
	wire [WIDTH*2-1+1:0] tmp01_59_39;
	wire [WIDTH*2-1+1:0] tmp01_59_40;
	wire [WIDTH*2-1+1:0] tmp01_59_41;
	wire [WIDTH*2-1+1:0] tmp01_59_42;
	wire [WIDTH*2-1+1:0] tmp01_59_43;
	wire [WIDTH*2-1+1:0] tmp01_59_44;
	wire [WIDTH*2-1+1:0] tmp01_59_45;
	wire [WIDTH*2-1+1:0] tmp01_59_46;
	wire [WIDTH*2-1+1:0] tmp01_59_47;
	wire [WIDTH*2-1+1:0] tmp01_59_48;
	wire [WIDTH*2-1+1:0] tmp01_59_49;
	wire [WIDTH*2-1+1:0] tmp01_59_50;
	wire [WIDTH*2-1+1:0] tmp01_59_51;
	wire [WIDTH*2-1+1:0] tmp01_59_52;
	wire [WIDTH*2-1+1:0] tmp01_59_53;
	wire [WIDTH*2-1+1:0] tmp01_59_54;
	wire [WIDTH*2-1+1:0] tmp01_59_55;
	wire [WIDTH*2-1+1:0] tmp01_59_56;
	wire [WIDTH*2-1+1:0] tmp01_59_57;
	wire [WIDTH*2-1+1:0] tmp01_59_58;
	wire [WIDTH*2-1+1:0] tmp01_59_59;
	wire [WIDTH*2-1+1:0] tmp01_59_60;
	wire [WIDTH*2-1+1:0] tmp01_59_61;
	wire [WIDTH*2-1+1:0] tmp01_59_62;
	wire [WIDTH*2-1+1:0] tmp01_59_63;
	wire [WIDTH*2-1+1:0] tmp01_59_64;
	wire [WIDTH*2-1+1:0] tmp01_59_65;
	wire [WIDTH*2-1+1:0] tmp01_59_66;
	wire [WIDTH*2-1+1:0] tmp01_59_67;
	wire [WIDTH*2-1+1:0] tmp01_59_68;
	wire [WIDTH*2-1+1:0] tmp01_59_69;
	wire [WIDTH*2-1+1:0] tmp01_59_70;
	wire [WIDTH*2-1+1:0] tmp01_59_71;
	wire [WIDTH*2-1+1:0] tmp01_59_72;
	wire [WIDTH*2-1+1:0] tmp01_59_73;
	wire [WIDTH*2-1+1:0] tmp01_59_74;
	wire [WIDTH*2-1+1:0] tmp01_59_75;
	wire [WIDTH*2-1+1:0] tmp01_59_76;
	wire [WIDTH*2-1+1:0] tmp01_59_77;
	wire [WIDTH*2-1+1:0] tmp01_59_78;
	wire [WIDTH*2-1+1:0] tmp01_59_79;
	wire [WIDTH*2-1+1:0] tmp01_59_80;
	wire [WIDTH*2-1+1:0] tmp01_59_81;
	wire [WIDTH*2-1+1:0] tmp01_59_82;
	wire [WIDTH*2-1+1:0] tmp01_59_83;
	wire [WIDTH*2-1+1:0] tmp01_60_0;
	wire [WIDTH*2-1+1:0] tmp01_60_1;
	wire [WIDTH*2-1+1:0] tmp01_60_2;
	wire [WIDTH*2-1+1:0] tmp01_60_3;
	wire [WIDTH*2-1+1:0] tmp01_60_4;
	wire [WIDTH*2-1+1:0] tmp01_60_5;
	wire [WIDTH*2-1+1:0] tmp01_60_6;
	wire [WIDTH*2-1+1:0] tmp01_60_7;
	wire [WIDTH*2-1+1:0] tmp01_60_8;
	wire [WIDTH*2-1+1:0] tmp01_60_9;
	wire [WIDTH*2-1+1:0] tmp01_60_10;
	wire [WIDTH*2-1+1:0] tmp01_60_11;
	wire [WIDTH*2-1+1:0] tmp01_60_12;
	wire [WIDTH*2-1+1:0] tmp01_60_13;
	wire [WIDTH*2-1+1:0] tmp01_60_14;
	wire [WIDTH*2-1+1:0] tmp01_60_15;
	wire [WIDTH*2-1+1:0] tmp01_60_16;
	wire [WIDTH*2-1+1:0] tmp01_60_17;
	wire [WIDTH*2-1+1:0] tmp01_60_18;
	wire [WIDTH*2-1+1:0] tmp01_60_19;
	wire [WIDTH*2-1+1:0] tmp01_60_20;
	wire [WIDTH*2-1+1:0] tmp01_60_21;
	wire [WIDTH*2-1+1:0] tmp01_60_22;
	wire [WIDTH*2-1+1:0] tmp01_60_23;
	wire [WIDTH*2-1+1:0] tmp01_60_24;
	wire [WIDTH*2-1+1:0] tmp01_60_25;
	wire [WIDTH*2-1+1:0] tmp01_60_26;
	wire [WIDTH*2-1+1:0] tmp01_60_27;
	wire [WIDTH*2-1+1:0] tmp01_60_28;
	wire [WIDTH*2-1+1:0] tmp01_60_29;
	wire [WIDTH*2-1+1:0] tmp01_60_30;
	wire [WIDTH*2-1+1:0] tmp01_60_31;
	wire [WIDTH*2-1+1:0] tmp01_60_32;
	wire [WIDTH*2-1+1:0] tmp01_60_33;
	wire [WIDTH*2-1+1:0] tmp01_60_34;
	wire [WIDTH*2-1+1:0] tmp01_60_35;
	wire [WIDTH*2-1+1:0] tmp01_60_36;
	wire [WIDTH*2-1+1:0] tmp01_60_37;
	wire [WIDTH*2-1+1:0] tmp01_60_38;
	wire [WIDTH*2-1+1:0] tmp01_60_39;
	wire [WIDTH*2-1+1:0] tmp01_60_40;
	wire [WIDTH*2-1+1:0] tmp01_60_41;
	wire [WIDTH*2-1+1:0] tmp01_60_42;
	wire [WIDTH*2-1+1:0] tmp01_60_43;
	wire [WIDTH*2-1+1:0] tmp01_60_44;
	wire [WIDTH*2-1+1:0] tmp01_60_45;
	wire [WIDTH*2-1+1:0] tmp01_60_46;
	wire [WIDTH*2-1+1:0] tmp01_60_47;
	wire [WIDTH*2-1+1:0] tmp01_60_48;
	wire [WIDTH*2-1+1:0] tmp01_60_49;
	wire [WIDTH*2-1+1:0] tmp01_60_50;
	wire [WIDTH*2-1+1:0] tmp01_60_51;
	wire [WIDTH*2-1+1:0] tmp01_60_52;
	wire [WIDTH*2-1+1:0] tmp01_60_53;
	wire [WIDTH*2-1+1:0] tmp01_60_54;
	wire [WIDTH*2-1+1:0] tmp01_60_55;
	wire [WIDTH*2-1+1:0] tmp01_60_56;
	wire [WIDTH*2-1+1:0] tmp01_60_57;
	wire [WIDTH*2-1+1:0] tmp01_60_58;
	wire [WIDTH*2-1+1:0] tmp01_60_59;
	wire [WIDTH*2-1+1:0] tmp01_60_60;
	wire [WIDTH*2-1+1:0] tmp01_60_61;
	wire [WIDTH*2-1+1:0] tmp01_60_62;
	wire [WIDTH*2-1+1:0] tmp01_60_63;
	wire [WIDTH*2-1+1:0] tmp01_60_64;
	wire [WIDTH*2-1+1:0] tmp01_60_65;
	wire [WIDTH*2-1+1:0] tmp01_60_66;
	wire [WIDTH*2-1+1:0] tmp01_60_67;
	wire [WIDTH*2-1+1:0] tmp01_60_68;
	wire [WIDTH*2-1+1:0] tmp01_60_69;
	wire [WIDTH*2-1+1:0] tmp01_60_70;
	wire [WIDTH*2-1+1:0] tmp01_60_71;
	wire [WIDTH*2-1+1:0] tmp01_60_72;
	wire [WIDTH*2-1+1:0] tmp01_60_73;
	wire [WIDTH*2-1+1:0] tmp01_60_74;
	wire [WIDTH*2-1+1:0] tmp01_60_75;
	wire [WIDTH*2-1+1:0] tmp01_60_76;
	wire [WIDTH*2-1+1:0] tmp01_60_77;
	wire [WIDTH*2-1+1:0] tmp01_60_78;
	wire [WIDTH*2-1+1:0] tmp01_60_79;
	wire [WIDTH*2-1+1:0] tmp01_60_80;
	wire [WIDTH*2-1+1:0] tmp01_60_81;
	wire [WIDTH*2-1+1:0] tmp01_60_82;
	wire [WIDTH*2-1+1:0] tmp01_60_83;
	wire [WIDTH*2-1+1:0] tmp01_61_0;
	wire [WIDTH*2-1+1:0] tmp01_61_1;
	wire [WIDTH*2-1+1:0] tmp01_61_2;
	wire [WIDTH*2-1+1:0] tmp01_61_3;
	wire [WIDTH*2-1+1:0] tmp01_61_4;
	wire [WIDTH*2-1+1:0] tmp01_61_5;
	wire [WIDTH*2-1+1:0] tmp01_61_6;
	wire [WIDTH*2-1+1:0] tmp01_61_7;
	wire [WIDTH*2-1+1:0] tmp01_61_8;
	wire [WIDTH*2-1+1:0] tmp01_61_9;
	wire [WIDTH*2-1+1:0] tmp01_61_10;
	wire [WIDTH*2-1+1:0] tmp01_61_11;
	wire [WIDTH*2-1+1:0] tmp01_61_12;
	wire [WIDTH*2-1+1:0] tmp01_61_13;
	wire [WIDTH*2-1+1:0] tmp01_61_14;
	wire [WIDTH*2-1+1:0] tmp01_61_15;
	wire [WIDTH*2-1+1:0] tmp01_61_16;
	wire [WIDTH*2-1+1:0] tmp01_61_17;
	wire [WIDTH*2-1+1:0] tmp01_61_18;
	wire [WIDTH*2-1+1:0] tmp01_61_19;
	wire [WIDTH*2-1+1:0] tmp01_61_20;
	wire [WIDTH*2-1+1:0] tmp01_61_21;
	wire [WIDTH*2-1+1:0] tmp01_61_22;
	wire [WIDTH*2-1+1:0] tmp01_61_23;
	wire [WIDTH*2-1+1:0] tmp01_61_24;
	wire [WIDTH*2-1+1:0] tmp01_61_25;
	wire [WIDTH*2-1+1:0] tmp01_61_26;
	wire [WIDTH*2-1+1:0] tmp01_61_27;
	wire [WIDTH*2-1+1:0] tmp01_61_28;
	wire [WIDTH*2-1+1:0] tmp01_61_29;
	wire [WIDTH*2-1+1:0] tmp01_61_30;
	wire [WIDTH*2-1+1:0] tmp01_61_31;
	wire [WIDTH*2-1+1:0] tmp01_61_32;
	wire [WIDTH*2-1+1:0] tmp01_61_33;
	wire [WIDTH*2-1+1:0] tmp01_61_34;
	wire [WIDTH*2-1+1:0] tmp01_61_35;
	wire [WIDTH*2-1+1:0] tmp01_61_36;
	wire [WIDTH*2-1+1:0] tmp01_61_37;
	wire [WIDTH*2-1+1:0] tmp01_61_38;
	wire [WIDTH*2-1+1:0] tmp01_61_39;
	wire [WIDTH*2-1+1:0] tmp01_61_40;
	wire [WIDTH*2-1+1:0] tmp01_61_41;
	wire [WIDTH*2-1+1:0] tmp01_61_42;
	wire [WIDTH*2-1+1:0] tmp01_61_43;
	wire [WIDTH*2-1+1:0] tmp01_61_44;
	wire [WIDTH*2-1+1:0] tmp01_61_45;
	wire [WIDTH*2-1+1:0] tmp01_61_46;
	wire [WIDTH*2-1+1:0] tmp01_61_47;
	wire [WIDTH*2-1+1:0] tmp01_61_48;
	wire [WIDTH*2-1+1:0] tmp01_61_49;
	wire [WIDTH*2-1+1:0] tmp01_61_50;
	wire [WIDTH*2-1+1:0] tmp01_61_51;
	wire [WIDTH*2-1+1:0] tmp01_61_52;
	wire [WIDTH*2-1+1:0] tmp01_61_53;
	wire [WIDTH*2-1+1:0] tmp01_61_54;
	wire [WIDTH*2-1+1:0] tmp01_61_55;
	wire [WIDTH*2-1+1:0] tmp01_61_56;
	wire [WIDTH*2-1+1:0] tmp01_61_57;
	wire [WIDTH*2-1+1:0] tmp01_61_58;
	wire [WIDTH*2-1+1:0] tmp01_61_59;
	wire [WIDTH*2-1+1:0] tmp01_61_60;
	wire [WIDTH*2-1+1:0] tmp01_61_61;
	wire [WIDTH*2-1+1:0] tmp01_61_62;
	wire [WIDTH*2-1+1:0] tmp01_61_63;
	wire [WIDTH*2-1+1:0] tmp01_61_64;
	wire [WIDTH*2-1+1:0] tmp01_61_65;
	wire [WIDTH*2-1+1:0] tmp01_61_66;
	wire [WIDTH*2-1+1:0] tmp01_61_67;
	wire [WIDTH*2-1+1:0] tmp01_61_68;
	wire [WIDTH*2-1+1:0] tmp01_61_69;
	wire [WIDTH*2-1+1:0] tmp01_61_70;
	wire [WIDTH*2-1+1:0] tmp01_61_71;
	wire [WIDTH*2-1+1:0] tmp01_61_72;
	wire [WIDTH*2-1+1:0] tmp01_61_73;
	wire [WIDTH*2-1+1:0] tmp01_61_74;
	wire [WIDTH*2-1+1:0] tmp01_61_75;
	wire [WIDTH*2-1+1:0] tmp01_61_76;
	wire [WIDTH*2-1+1:0] tmp01_61_77;
	wire [WIDTH*2-1+1:0] tmp01_61_78;
	wire [WIDTH*2-1+1:0] tmp01_61_79;
	wire [WIDTH*2-1+1:0] tmp01_61_80;
	wire [WIDTH*2-1+1:0] tmp01_61_81;
	wire [WIDTH*2-1+1:0] tmp01_61_82;
	wire [WIDTH*2-1+1:0] tmp01_61_83;
	wire [WIDTH*2-1+1:0] tmp01_62_0;
	wire [WIDTH*2-1+1:0] tmp01_62_1;
	wire [WIDTH*2-1+1:0] tmp01_62_2;
	wire [WIDTH*2-1+1:0] tmp01_62_3;
	wire [WIDTH*2-1+1:0] tmp01_62_4;
	wire [WIDTH*2-1+1:0] tmp01_62_5;
	wire [WIDTH*2-1+1:0] tmp01_62_6;
	wire [WIDTH*2-1+1:0] tmp01_62_7;
	wire [WIDTH*2-1+1:0] tmp01_62_8;
	wire [WIDTH*2-1+1:0] tmp01_62_9;
	wire [WIDTH*2-1+1:0] tmp01_62_10;
	wire [WIDTH*2-1+1:0] tmp01_62_11;
	wire [WIDTH*2-1+1:0] tmp01_62_12;
	wire [WIDTH*2-1+1:0] tmp01_62_13;
	wire [WIDTH*2-1+1:0] tmp01_62_14;
	wire [WIDTH*2-1+1:0] tmp01_62_15;
	wire [WIDTH*2-1+1:0] tmp01_62_16;
	wire [WIDTH*2-1+1:0] tmp01_62_17;
	wire [WIDTH*2-1+1:0] tmp01_62_18;
	wire [WIDTH*2-1+1:0] tmp01_62_19;
	wire [WIDTH*2-1+1:0] tmp01_62_20;
	wire [WIDTH*2-1+1:0] tmp01_62_21;
	wire [WIDTH*2-1+1:0] tmp01_62_22;
	wire [WIDTH*2-1+1:0] tmp01_62_23;
	wire [WIDTH*2-1+1:0] tmp01_62_24;
	wire [WIDTH*2-1+1:0] tmp01_62_25;
	wire [WIDTH*2-1+1:0] tmp01_62_26;
	wire [WIDTH*2-1+1:0] tmp01_62_27;
	wire [WIDTH*2-1+1:0] tmp01_62_28;
	wire [WIDTH*2-1+1:0] tmp01_62_29;
	wire [WIDTH*2-1+1:0] tmp01_62_30;
	wire [WIDTH*2-1+1:0] tmp01_62_31;
	wire [WIDTH*2-1+1:0] tmp01_62_32;
	wire [WIDTH*2-1+1:0] tmp01_62_33;
	wire [WIDTH*2-1+1:0] tmp01_62_34;
	wire [WIDTH*2-1+1:0] tmp01_62_35;
	wire [WIDTH*2-1+1:0] tmp01_62_36;
	wire [WIDTH*2-1+1:0] tmp01_62_37;
	wire [WIDTH*2-1+1:0] tmp01_62_38;
	wire [WIDTH*2-1+1:0] tmp01_62_39;
	wire [WIDTH*2-1+1:0] tmp01_62_40;
	wire [WIDTH*2-1+1:0] tmp01_62_41;
	wire [WIDTH*2-1+1:0] tmp01_62_42;
	wire [WIDTH*2-1+1:0] tmp01_62_43;
	wire [WIDTH*2-1+1:0] tmp01_62_44;
	wire [WIDTH*2-1+1:0] tmp01_62_45;
	wire [WIDTH*2-1+1:0] tmp01_62_46;
	wire [WIDTH*2-1+1:0] tmp01_62_47;
	wire [WIDTH*2-1+1:0] tmp01_62_48;
	wire [WIDTH*2-1+1:0] tmp01_62_49;
	wire [WIDTH*2-1+1:0] tmp01_62_50;
	wire [WIDTH*2-1+1:0] tmp01_62_51;
	wire [WIDTH*2-1+1:0] tmp01_62_52;
	wire [WIDTH*2-1+1:0] tmp01_62_53;
	wire [WIDTH*2-1+1:0] tmp01_62_54;
	wire [WIDTH*2-1+1:0] tmp01_62_55;
	wire [WIDTH*2-1+1:0] tmp01_62_56;
	wire [WIDTH*2-1+1:0] tmp01_62_57;
	wire [WIDTH*2-1+1:0] tmp01_62_58;
	wire [WIDTH*2-1+1:0] tmp01_62_59;
	wire [WIDTH*2-1+1:0] tmp01_62_60;
	wire [WIDTH*2-1+1:0] tmp01_62_61;
	wire [WIDTH*2-1+1:0] tmp01_62_62;
	wire [WIDTH*2-1+1:0] tmp01_62_63;
	wire [WIDTH*2-1+1:0] tmp01_62_64;
	wire [WIDTH*2-1+1:0] tmp01_62_65;
	wire [WIDTH*2-1+1:0] tmp01_62_66;
	wire [WIDTH*2-1+1:0] tmp01_62_67;
	wire [WIDTH*2-1+1:0] tmp01_62_68;
	wire [WIDTH*2-1+1:0] tmp01_62_69;
	wire [WIDTH*2-1+1:0] tmp01_62_70;
	wire [WIDTH*2-1+1:0] tmp01_62_71;
	wire [WIDTH*2-1+1:0] tmp01_62_72;
	wire [WIDTH*2-1+1:0] tmp01_62_73;
	wire [WIDTH*2-1+1:0] tmp01_62_74;
	wire [WIDTH*2-1+1:0] tmp01_62_75;
	wire [WIDTH*2-1+1:0] tmp01_62_76;
	wire [WIDTH*2-1+1:0] tmp01_62_77;
	wire [WIDTH*2-1+1:0] tmp01_62_78;
	wire [WIDTH*2-1+1:0] tmp01_62_79;
	wire [WIDTH*2-1+1:0] tmp01_62_80;
	wire [WIDTH*2-1+1:0] tmp01_62_81;
	wire [WIDTH*2-1+1:0] tmp01_62_82;
	wire [WIDTH*2-1+1:0] tmp01_62_83;
	wire [WIDTH*2-1+1:0] tmp01_63_0;
	wire [WIDTH*2-1+1:0] tmp01_63_1;
	wire [WIDTH*2-1+1:0] tmp01_63_2;
	wire [WIDTH*2-1+1:0] tmp01_63_3;
	wire [WIDTH*2-1+1:0] tmp01_63_4;
	wire [WIDTH*2-1+1:0] tmp01_63_5;
	wire [WIDTH*2-1+1:0] tmp01_63_6;
	wire [WIDTH*2-1+1:0] tmp01_63_7;
	wire [WIDTH*2-1+1:0] tmp01_63_8;
	wire [WIDTH*2-1+1:0] tmp01_63_9;
	wire [WIDTH*2-1+1:0] tmp01_63_10;
	wire [WIDTH*2-1+1:0] tmp01_63_11;
	wire [WIDTH*2-1+1:0] tmp01_63_12;
	wire [WIDTH*2-1+1:0] tmp01_63_13;
	wire [WIDTH*2-1+1:0] tmp01_63_14;
	wire [WIDTH*2-1+1:0] tmp01_63_15;
	wire [WIDTH*2-1+1:0] tmp01_63_16;
	wire [WIDTH*2-1+1:0] tmp01_63_17;
	wire [WIDTH*2-1+1:0] tmp01_63_18;
	wire [WIDTH*2-1+1:0] tmp01_63_19;
	wire [WIDTH*2-1+1:0] tmp01_63_20;
	wire [WIDTH*2-1+1:0] tmp01_63_21;
	wire [WIDTH*2-1+1:0] tmp01_63_22;
	wire [WIDTH*2-1+1:0] tmp01_63_23;
	wire [WIDTH*2-1+1:0] tmp01_63_24;
	wire [WIDTH*2-1+1:0] tmp01_63_25;
	wire [WIDTH*2-1+1:0] tmp01_63_26;
	wire [WIDTH*2-1+1:0] tmp01_63_27;
	wire [WIDTH*2-1+1:0] tmp01_63_28;
	wire [WIDTH*2-1+1:0] tmp01_63_29;
	wire [WIDTH*2-1+1:0] tmp01_63_30;
	wire [WIDTH*2-1+1:0] tmp01_63_31;
	wire [WIDTH*2-1+1:0] tmp01_63_32;
	wire [WIDTH*2-1+1:0] tmp01_63_33;
	wire [WIDTH*2-1+1:0] tmp01_63_34;
	wire [WIDTH*2-1+1:0] tmp01_63_35;
	wire [WIDTH*2-1+1:0] tmp01_63_36;
	wire [WIDTH*2-1+1:0] tmp01_63_37;
	wire [WIDTH*2-1+1:0] tmp01_63_38;
	wire [WIDTH*2-1+1:0] tmp01_63_39;
	wire [WIDTH*2-1+1:0] tmp01_63_40;
	wire [WIDTH*2-1+1:0] tmp01_63_41;
	wire [WIDTH*2-1+1:0] tmp01_63_42;
	wire [WIDTH*2-1+1:0] tmp01_63_43;
	wire [WIDTH*2-1+1:0] tmp01_63_44;
	wire [WIDTH*2-1+1:0] tmp01_63_45;
	wire [WIDTH*2-1+1:0] tmp01_63_46;
	wire [WIDTH*2-1+1:0] tmp01_63_47;
	wire [WIDTH*2-1+1:0] tmp01_63_48;
	wire [WIDTH*2-1+1:0] tmp01_63_49;
	wire [WIDTH*2-1+1:0] tmp01_63_50;
	wire [WIDTH*2-1+1:0] tmp01_63_51;
	wire [WIDTH*2-1+1:0] tmp01_63_52;
	wire [WIDTH*2-1+1:0] tmp01_63_53;
	wire [WIDTH*2-1+1:0] tmp01_63_54;
	wire [WIDTH*2-1+1:0] tmp01_63_55;
	wire [WIDTH*2-1+1:0] tmp01_63_56;
	wire [WIDTH*2-1+1:0] tmp01_63_57;
	wire [WIDTH*2-1+1:0] tmp01_63_58;
	wire [WIDTH*2-1+1:0] tmp01_63_59;
	wire [WIDTH*2-1+1:0] tmp01_63_60;
	wire [WIDTH*2-1+1:0] tmp01_63_61;
	wire [WIDTH*2-1+1:0] tmp01_63_62;
	wire [WIDTH*2-1+1:0] tmp01_63_63;
	wire [WIDTH*2-1+1:0] tmp01_63_64;
	wire [WIDTH*2-1+1:0] tmp01_63_65;
	wire [WIDTH*2-1+1:0] tmp01_63_66;
	wire [WIDTH*2-1+1:0] tmp01_63_67;
	wire [WIDTH*2-1+1:0] tmp01_63_68;
	wire [WIDTH*2-1+1:0] tmp01_63_69;
	wire [WIDTH*2-1+1:0] tmp01_63_70;
	wire [WIDTH*2-1+1:0] tmp01_63_71;
	wire [WIDTH*2-1+1:0] tmp01_63_72;
	wire [WIDTH*2-1+1:0] tmp01_63_73;
	wire [WIDTH*2-1+1:0] tmp01_63_74;
	wire [WIDTH*2-1+1:0] tmp01_63_75;
	wire [WIDTH*2-1+1:0] tmp01_63_76;
	wire [WIDTH*2-1+1:0] tmp01_63_77;
	wire [WIDTH*2-1+1:0] tmp01_63_78;
	wire [WIDTH*2-1+1:0] tmp01_63_79;
	wire [WIDTH*2-1+1:0] tmp01_63_80;
	wire [WIDTH*2-1+1:0] tmp01_63_81;
	wire [WIDTH*2-1+1:0] tmp01_63_82;
	wire [WIDTH*2-1+1:0] tmp01_63_83;
	wire [WIDTH*2-1+2:0] tmp02_0_0;
	wire [WIDTH*2-1+2:0] tmp02_0_1;
	wire [WIDTH*2-1+2:0] tmp02_0_2;
	wire [WIDTH*2-1+2:0] tmp02_0_3;
	wire [WIDTH*2-1+2:0] tmp02_0_4;
	wire [WIDTH*2-1+2:0] tmp02_0_5;
	wire [WIDTH*2-1+2:0] tmp02_0_6;
	wire [WIDTH*2-1+2:0] tmp02_0_7;
	wire [WIDTH*2-1+2:0] tmp02_0_8;
	wire [WIDTH*2-1+2:0] tmp02_0_9;
	wire [WIDTH*2-1+2:0] tmp02_0_10;
	wire [WIDTH*2-1+2:0] tmp02_0_11;
	wire [WIDTH*2-1+2:0] tmp02_0_12;
	wire [WIDTH*2-1+2:0] tmp02_0_13;
	wire [WIDTH*2-1+2:0] tmp02_0_14;
	wire [WIDTH*2-1+2:0] tmp02_0_15;
	wire [WIDTH*2-1+2:0] tmp02_0_16;
	wire [WIDTH*2-1+2:0] tmp02_0_17;
	wire [WIDTH*2-1+2:0] tmp02_0_18;
	wire [WIDTH*2-1+2:0] tmp02_0_19;
	wire [WIDTH*2-1+2:0] tmp02_0_20;
	wire [WIDTH*2-1+2:0] tmp02_0_21;
	wire [WIDTH*2-1+2:0] tmp02_0_22;
	wire [WIDTH*2-1+2:0] tmp02_0_23;
	wire [WIDTH*2-1+2:0] tmp02_0_24;
	wire [WIDTH*2-1+2:0] tmp02_0_25;
	wire [WIDTH*2-1+2:0] tmp02_0_26;
	wire [WIDTH*2-1+2:0] tmp02_0_27;
	wire [WIDTH*2-1+2:0] tmp02_0_28;
	wire [WIDTH*2-1+2:0] tmp02_0_29;
	wire [WIDTH*2-1+2:0] tmp02_0_30;
	wire [WIDTH*2-1+2:0] tmp02_0_31;
	wire [WIDTH*2-1+2:0] tmp02_0_32;
	wire [WIDTH*2-1+2:0] tmp02_0_33;
	wire [WIDTH*2-1+2:0] tmp02_0_34;
	wire [WIDTH*2-1+2:0] tmp02_0_35;
	wire [WIDTH*2-1+2:0] tmp02_0_36;
	wire [WIDTH*2-1+2:0] tmp02_0_37;
	wire [WIDTH*2-1+2:0] tmp02_0_38;
	wire [WIDTH*2-1+2:0] tmp02_0_39;
	wire [WIDTH*2-1+2:0] tmp02_0_40;
	wire [WIDTH*2-1+2:0] tmp02_0_41;
	wire [WIDTH*2-1+2:0] tmp02_0_42;
	wire [WIDTH*2-1+2:0] tmp02_0_43;
	wire [WIDTH*2-1+2:0] tmp02_0_44;
	wire [WIDTH*2-1+2:0] tmp02_0_45;
	wire [WIDTH*2-1+2:0] tmp02_0_46;
	wire [WIDTH*2-1+2:0] tmp02_0_47;
	wire [WIDTH*2-1+2:0] tmp02_0_48;
	wire [WIDTH*2-1+2:0] tmp02_0_49;
	wire [WIDTH*2-1+2:0] tmp02_0_50;
	wire [WIDTH*2-1+2:0] tmp02_0_51;
	wire [WIDTH*2-1+2:0] tmp02_0_52;
	wire [WIDTH*2-1+2:0] tmp02_0_53;
	wire [WIDTH*2-1+2:0] tmp02_0_54;
	wire [WIDTH*2-1+2:0] tmp02_0_55;
	wire [WIDTH*2-1+2:0] tmp02_0_56;
	wire [WIDTH*2-1+2:0] tmp02_0_57;
	wire [WIDTH*2-1+2:0] tmp02_0_58;
	wire [WIDTH*2-1+2:0] tmp02_0_59;
	wire [WIDTH*2-1+2:0] tmp02_0_60;
	wire [WIDTH*2-1+2:0] tmp02_0_61;
	wire [WIDTH*2-1+2:0] tmp02_0_62;
	wire [WIDTH*2-1+2:0] tmp02_0_63;
	wire [WIDTH*2-1+2:0] tmp02_0_64;
	wire [WIDTH*2-1+2:0] tmp02_0_65;
	wire [WIDTH*2-1+2:0] tmp02_0_66;
	wire [WIDTH*2-1+2:0] tmp02_0_67;
	wire [WIDTH*2-1+2:0] tmp02_0_68;
	wire [WIDTH*2-1+2:0] tmp02_0_69;
	wire [WIDTH*2-1+2:0] tmp02_0_70;
	wire [WIDTH*2-1+2:0] tmp02_0_71;
	wire [WIDTH*2-1+2:0] tmp02_0_72;
	wire [WIDTH*2-1+2:0] tmp02_0_73;
	wire [WIDTH*2-1+2:0] tmp02_0_74;
	wire [WIDTH*2-1+2:0] tmp02_0_75;
	wire [WIDTH*2-1+2:0] tmp02_0_76;
	wire [WIDTH*2-1+2:0] tmp02_0_77;
	wire [WIDTH*2-1+2:0] tmp02_0_78;
	wire [WIDTH*2-1+2:0] tmp02_0_79;
	wire [WIDTH*2-1+2:0] tmp02_0_80;
	wire [WIDTH*2-1+2:0] tmp02_0_81;
	wire [WIDTH*2-1+2:0] tmp02_0_82;
	wire [WIDTH*2-1+2:0] tmp02_0_83;
	wire [WIDTH*2-1+2:0] tmp02_1_0;
	wire [WIDTH*2-1+2:0] tmp02_1_1;
	wire [WIDTH*2-1+2:0] tmp02_1_2;
	wire [WIDTH*2-1+2:0] tmp02_1_3;
	wire [WIDTH*2-1+2:0] tmp02_1_4;
	wire [WIDTH*2-1+2:0] tmp02_1_5;
	wire [WIDTH*2-1+2:0] tmp02_1_6;
	wire [WIDTH*2-1+2:0] tmp02_1_7;
	wire [WIDTH*2-1+2:0] tmp02_1_8;
	wire [WIDTH*2-1+2:0] tmp02_1_9;
	wire [WIDTH*2-1+2:0] tmp02_1_10;
	wire [WIDTH*2-1+2:0] tmp02_1_11;
	wire [WIDTH*2-1+2:0] tmp02_1_12;
	wire [WIDTH*2-1+2:0] tmp02_1_13;
	wire [WIDTH*2-1+2:0] tmp02_1_14;
	wire [WIDTH*2-1+2:0] tmp02_1_15;
	wire [WIDTH*2-1+2:0] tmp02_1_16;
	wire [WIDTH*2-1+2:0] tmp02_1_17;
	wire [WIDTH*2-1+2:0] tmp02_1_18;
	wire [WIDTH*2-1+2:0] tmp02_1_19;
	wire [WIDTH*2-1+2:0] tmp02_1_20;
	wire [WIDTH*2-1+2:0] tmp02_1_21;
	wire [WIDTH*2-1+2:0] tmp02_1_22;
	wire [WIDTH*2-1+2:0] tmp02_1_23;
	wire [WIDTH*2-1+2:0] tmp02_1_24;
	wire [WIDTH*2-1+2:0] tmp02_1_25;
	wire [WIDTH*2-1+2:0] tmp02_1_26;
	wire [WIDTH*2-1+2:0] tmp02_1_27;
	wire [WIDTH*2-1+2:0] tmp02_1_28;
	wire [WIDTH*2-1+2:0] tmp02_1_29;
	wire [WIDTH*2-1+2:0] tmp02_1_30;
	wire [WIDTH*2-1+2:0] tmp02_1_31;
	wire [WIDTH*2-1+2:0] tmp02_1_32;
	wire [WIDTH*2-1+2:0] tmp02_1_33;
	wire [WIDTH*2-1+2:0] tmp02_1_34;
	wire [WIDTH*2-1+2:0] tmp02_1_35;
	wire [WIDTH*2-1+2:0] tmp02_1_36;
	wire [WIDTH*2-1+2:0] tmp02_1_37;
	wire [WIDTH*2-1+2:0] tmp02_1_38;
	wire [WIDTH*2-1+2:0] tmp02_1_39;
	wire [WIDTH*2-1+2:0] tmp02_1_40;
	wire [WIDTH*2-1+2:0] tmp02_1_41;
	wire [WIDTH*2-1+2:0] tmp02_1_42;
	wire [WIDTH*2-1+2:0] tmp02_1_43;
	wire [WIDTH*2-1+2:0] tmp02_1_44;
	wire [WIDTH*2-1+2:0] tmp02_1_45;
	wire [WIDTH*2-1+2:0] tmp02_1_46;
	wire [WIDTH*2-1+2:0] tmp02_1_47;
	wire [WIDTH*2-1+2:0] tmp02_1_48;
	wire [WIDTH*2-1+2:0] tmp02_1_49;
	wire [WIDTH*2-1+2:0] tmp02_1_50;
	wire [WIDTH*2-1+2:0] tmp02_1_51;
	wire [WIDTH*2-1+2:0] tmp02_1_52;
	wire [WIDTH*2-1+2:0] tmp02_1_53;
	wire [WIDTH*2-1+2:0] tmp02_1_54;
	wire [WIDTH*2-1+2:0] tmp02_1_55;
	wire [WIDTH*2-1+2:0] tmp02_1_56;
	wire [WIDTH*2-1+2:0] tmp02_1_57;
	wire [WIDTH*2-1+2:0] tmp02_1_58;
	wire [WIDTH*2-1+2:0] tmp02_1_59;
	wire [WIDTH*2-1+2:0] tmp02_1_60;
	wire [WIDTH*2-1+2:0] tmp02_1_61;
	wire [WIDTH*2-1+2:0] tmp02_1_62;
	wire [WIDTH*2-1+2:0] tmp02_1_63;
	wire [WIDTH*2-1+2:0] tmp02_1_64;
	wire [WIDTH*2-1+2:0] tmp02_1_65;
	wire [WIDTH*2-1+2:0] tmp02_1_66;
	wire [WIDTH*2-1+2:0] tmp02_1_67;
	wire [WIDTH*2-1+2:0] tmp02_1_68;
	wire [WIDTH*2-1+2:0] tmp02_1_69;
	wire [WIDTH*2-1+2:0] tmp02_1_70;
	wire [WIDTH*2-1+2:0] tmp02_1_71;
	wire [WIDTH*2-1+2:0] tmp02_1_72;
	wire [WIDTH*2-1+2:0] tmp02_1_73;
	wire [WIDTH*2-1+2:0] tmp02_1_74;
	wire [WIDTH*2-1+2:0] tmp02_1_75;
	wire [WIDTH*2-1+2:0] tmp02_1_76;
	wire [WIDTH*2-1+2:0] tmp02_1_77;
	wire [WIDTH*2-1+2:0] tmp02_1_78;
	wire [WIDTH*2-1+2:0] tmp02_1_79;
	wire [WIDTH*2-1+2:0] tmp02_1_80;
	wire [WIDTH*2-1+2:0] tmp02_1_81;
	wire [WIDTH*2-1+2:0] tmp02_1_82;
	wire [WIDTH*2-1+2:0] tmp02_1_83;
	wire [WIDTH*2-1+2:0] tmp02_2_0;
	wire [WIDTH*2-1+2:0] tmp02_2_1;
	wire [WIDTH*2-1+2:0] tmp02_2_2;
	wire [WIDTH*2-1+2:0] tmp02_2_3;
	wire [WIDTH*2-1+2:0] tmp02_2_4;
	wire [WIDTH*2-1+2:0] tmp02_2_5;
	wire [WIDTH*2-1+2:0] tmp02_2_6;
	wire [WIDTH*2-1+2:0] tmp02_2_7;
	wire [WIDTH*2-1+2:0] tmp02_2_8;
	wire [WIDTH*2-1+2:0] tmp02_2_9;
	wire [WIDTH*2-1+2:0] tmp02_2_10;
	wire [WIDTH*2-1+2:0] tmp02_2_11;
	wire [WIDTH*2-1+2:0] tmp02_2_12;
	wire [WIDTH*2-1+2:0] tmp02_2_13;
	wire [WIDTH*2-1+2:0] tmp02_2_14;
	wire [WIDTH*2-1+2:0] tmp02_2_15;
	wire [WIDTH*2-1+2:0] tmp02_2_16;
	wire [WIDTH*2-1+2:0] tmp02_2_17;
	wire [WIDTH*2-1+2:0] tmp02_2_18;
	wire [WIDTH*2-1+2:0] tmp02_2_19;
	wire [WIDTH*2-1+2:0] tmp02_2_20;
	wire [WIDTH*2-1+2:0] tmp02_2_21;
	wire [WIDTH*2-1+2:0] tmp02_2_22;
	wire [WIDTH*2-1+2:0] tmp02_2_23;
	wire [WIDTH*2-1+2:0] tmp02_2_24;
	wire [WIDTH*2-1+2:0] tmp02_2_25;
	wire [WIDTH*2-1+2:0] tmp02_2_26;
	wire [WIDTH*2-1+2:0] tmp02_2_27;
	wire [WIDTH*2-1+2:0] tmp02_2_28;
	wire [WIDTH*2-1+2:0] tmp02_2_29;
	wire [WIDTH*2-1+2:0] tmp02_2_30;
	wire [WIDTH*2-1+2:0] tmp02_2_31;
	wire [WIDTH*2-1+2:0] tmp02_2_32;
	wire [WIDTH*2-1+2:0] tmp02_2_33;
	wire [WIDTH*2-1+2:0] tmp02_2_34;
	wire [WIDTH*2-1+2:0] tmp02_2_35;
	wire [WIDTH*2-1+2:0] tmp02_2_36;
	wire [WIDTH*2-1+2:0] tmp02_2_37;
	wire [WIDTH*2-1+2:0] tmp02_2_38;
	wire [WIDTH*2-1+2:0] tmp02_2_39;
	wire [WIDTH*2-1+2:0] tmp02_2_40;
	wire [WIDTH*2-1+2:0] tmp02_2_41;
	wire [WIDTH*2-1+2:0] tmp02_2_42;
	wire [WIDTH*2-1+2:0] tmp02_2_43;
	wire [WIDTH*2-1+2:0] tmp02_2_44;
	wire [WIDTH*2-1+2:0] tmp02_2_45;
	wire [WIDTH*2-1+2:0] tmp02_2_46;
	wire [WIDTH*2-1+2:0] tmp02_2_47;
	wire [WIDTH*2-1+2:0] tmp02_2_48;
	wire [WIDTH*2-1+2:0] tmp02_2_49;
	wire [WIDTH*2-1+2:0] tmp02_2_50;
	wire [WIDTH*2-1+2:0] tmp02_2_51;
	wire [WIDTH*2-1+2:0] tmp02_2_52;
	wire [WIDTH*2-1+2:0] tmp02_2_53;
	wire [WIDTH*2-1+2:0] tmp02_2_54;
	wire [WIDTH*2-1+2:0] tmp02_2_55;
	wire [WIDTH*2-1+2:0] tmp02_2_56;
	wire [WIDTH*2-1+2:0] tmp02_2_57;
	wire [WIDTH*2-1+2:0] tmp02_2_58;
	wire [WIDTH*2-1+2:0] tmp02_2_59;
	wire [WIDTH*2-1+2:0] tmp02_2_60;
	wire [WIDTH*2-1+2:0] tmp02_2_61;
	wire [WIDTH*2-1+2:0] tmp02_2_62;
	wire [WIDTH*2-1+2:0] tmp02_2_63;
	wire [WIDTH*2-1+2:0] tmp02_2_64;
	wire [WIDTH*2-1+2:0] tmp02_2_65;
	wire [WIDTH*2-1+2:0] tmp02_2_66;
	wire [WIDTH*2-1+2:0] tmp02_2_67;
	wire [WIDTH*2-1+2:0] tmp02_2_68;
	wire [WIDTH*2-1+2:0] tmp02_2_69;
	wire [WIDTH*2-1+2:0] tmp02_2_70;
	wire [WIDTH*2-1+2:0] tmp02_2_71;
	wire [WIDTH*2-1+2:0] tmp02_2_72;
	wire [WIDTH*2-1+2:0] tmp02_2_73;
	wire [WIDTH*2-1+2:0] tmp02_2_74;
	wire [WIDTH*2-1+2:0] tmp02_2_75;
	wire [WIDTH*2-1+2:0] tmp02_2_76;
	wire [WIDTH*2-1+2:0] tmp02_2_77;
	wire [WIDTH*2-1+2:0] tmp02_2_78;
	wire [WIDTH*2-1+2:0] tmp02_2_79;
	wire [WIDTH*2-1+2:0] tmp02_2_80;
	wire [WIDTH*2-1+2:0] tmp02_2_81;
	wire [WIDTH*2-1+2:0] tmp02_2_82;
	wire [WIDTH*2-1+2:0] tmp02_2_83;
	wire [WIDTH*2-1+2:0] tmp02_3_0;
	wire [WIDTH*2-1+2:0] tmp02_3_1;
	wire [WIDTH*2-1+2:0] tmp02_3_2;
	wire [WIDTH*2-1+2:0] tmp02_3_3;
	wire [WIDTH*2-1+2:0] tmp02_3_4;
	wire [WIDTH*2-1+2:0] tmp02_3_5;
	wire [WIDTH*2-1+2:0] tmp02_3_6;
	wire [WIDTH*2-1+2:0] tmp02_3_7;
	wire [WIDTH*2-1+2:0] tmp02_3_8;
	wire [WIDTH*2-1+2:0] tmp02_3_9;
	wire [WIDTH*2-1+2:0] tmp02_3_10;
	wire [WIDTH*2-1+2:0] tmp02_3_11;
	wire [WIDTH*2-1+2:0] tmp02_3_12;
	wire [WIDTH*2-1+2:0] tmp02_3_13;
	wire [WIDTH*2-1+2:0] tmp02_3_14;
	wire [WIDTH*2-1+2:0] tmp02_3_15;
	wire [WIDTH*2-1+2:0] tmp02_3_16;
	wire [WIDTH*2-1+2:0] tmp02_3_17;
	wire [WIDTH*2-1+2:0] tmp02_3_18;
	wire [WIDTH*2-1+2:0] tmp02_3_19;
	wire [WIDTH*2-1+2:0] tmp02_3_20;
	wire [WIDTH*2-1+2:0] tmp02_3_21;
	wire [WIDTH*2-1+2:0] tmp02_3_22;
	wire [WIDTH*2-1+2:0] tmp02_3_23;
	wire [WIDTH*2-1+2:0] tmp02_3_24;
	wire [WIDTH*2-1+2:0] tmp02_3_25;
	wire [WIDTH*2-1+2:0] tmp02_3_26;
	wire [WIDTH*2-1+2:0] tmp02_3_27;
	wire [WIDTH*2-1+2:0] tmp02_3_28;
	wire [WIDTH*2-1+2:0] tmp02_3_29;
	wire [WIDTH*2-1+2:0] tmp02_3_30;
	wire [WIDTH*2-1+2:0] tmp02_3_31;
	wire [WIDTH*2-1+2:0] tmp02_3_32;
	wire [WIDTH*2-1+2:0] tmp02_3_33;
	wire [WIDTH*2-1+2:0] tmp02_3_34;
	wire [WIDTH*2-1+2:0] tmp02_3_35;
	wire [WIDTH*2-1+2:0] tmp02_3_36;
	wire [WIDTH*2-1+2:0] tmp02_3_37;
	wire [WIDTH*2-1+2:0] tmp02_3_38;
	wire [WIDTH*2-1+2:0] tmp02_3_39;
	wire [WIDTH*2-1+2:0] tmp02_3_40;
	wire [WIDTH*2-1+2:0] tmp02_3_41;
	wire [WIDTH*2-1+2:0] tmp02_3_42;
	wire [WIDTH*2-1+2:0] tmp02_3_43;
	wire [WIDTH*2-1+2:0] tmp02_3_44;
	wire [WIDTH*2-1+2:0] tmp02_3_45;
	wire [WIDTH*2-1+2:0] tmp02_3_46;
	wire [WIDTH*2-1+2:0] tmp02_3_47;
	wire [WIDTH*2-1+2:0] tmp02_3_48;
	wire [WIDTH*2-1+2:0] tmp02_3_49;
	wire [WIDTH*2-1+2:0] tmp02_3_50;
	wire [WIDTH*2-1+2:0] tmp02_3_51;
	wire [WIDTH*2-1+2:0] tmp02_3_52;
	wire [WIDTH*2-1+2:0] tmp02_3_53;
	wire [WIDTH*2-1+2:0] tmp02_3_54;
	wire [WIDTH*2-1+2:0] tmp02_3_55;
	wire [WIDTH*2-1+2:0] tmp02_3_56;
	wire [WIDTH*2-1+2:0] tmp02_3_57;
	wire [WIDTH*2-1+2:0] tmp02_3_58;
	wire [WIDTH*2-1+2:0] tmp02_3_59;
	wire [WIDTH*2-1+2:0] tmp02_3_60;
	wire [WIDTH*2-1+2:0] tmp02_3_61;
	wire [WIDTH*2-1+2:0] tmp02_3_62;
	wire [WIDTH*2-1+2:0] tmp02_3_63;
	wire [WIDTH*2-1+2:0] tmp02_3_64;
	wire [WIDTH*2-1+2:0] tmp02_3_65;
	wire [WIDTH*2-1+2:0] tmp02_3_66;
	wire [WIDTH*2-1+2:0] tmp02_3_67;
	wire [WIDTH*2-1+2:0] tmp02_3_68;
	wire [WIDTH*2-1+2:0] tmp02_3_69;
	wire [WIDTH*2-1+2:0] tmp02_3_70;
	wire [WIDTH*2-1+2:0] tmp02_3_71;
	wire [WIDTH*2-1+2:0] tmp02_3_72;
	wire [WIDTH*2-1+2:0] tmp02_3_73;
	wire [WIDTH*2-1+2:0] tmp02_3_74;
	wire [WIDTH*2-1+2:0] tmp02_3_75;
	wire [WIDTH*2-1+2:0] tmp02_3_76;
	wire [WIDTH*2-1+2:0] tmp02_3_77;
	wire [WIDTH*2-1+2:0] tmp02_3_78;
	wire [WIDTH*2-1+2:0] tmp02_3_79;
	wire [WIDTH*2-1+2:0] tmp02_3_80;
	wire [WIDTH*2-1+2:0] tmp02_3_81;
	wire [WIDTH*2-1+2:0] tmp02_3_82;
	wire [WIDTH*2-1+2:0] tmp02_3_83;
	wire [WIDTH*2-1+2:0] tmp02_4_0;
	wire [WIDTH*2-1+2:0] tmp02_4_1;
	wire [WIDTH*2-1+2:0] tmp02_4_2;
	wire [WIDTH*2-1+2:0] tmp02_4_3;
	wire [WIDTH*2-1+2:0] tmp02_4_4;
	wire [WIDTH*2-1+2:0] tmp02_4_5;
	wire [WIDTH*2-1+2:0] tmp02_4_6;
	wire [WIDTH*2-1+2:0] tmp02_4_7;
	wire [WIDTH*2-1+2:0] tmp02_4_8;
	wire [WIDTH*2-1+2:0] tmp02_4_9;
	wire [WIDTH*2-1+2:0] tmp02_4_10;
	wire [WIDTH*2-1+2:0] tmp02_4_11;
	wire [WIDTH*2-1+2:0] tmp02_4_12;
	wire [WIDTH*2-1+2:0] tmp02_4_13;
	wire [WIDTH*2-1+2:0] tmp02_4_14;
	wire [WIDTH*2-1+2:0] tmp02_4_15;
	wire [WIDTH*2-1+2:0] tmp02_4_16;
	wire [WIDTH*2-1+2:0] tmp02_4_17;
	wire [WIDTH*2-1+2:0] tmp02_4_18;
	wire [WIDTH*2-1+2:0] tmp02_4_19;
	wire [WIDTH*2-1+2:0] tmp02_4_20;
	wire [WIDTH*2-1+2:0] tmp02_4_21;
	wire [WIDTH*2-1+2:0] tmp02_4_22;
	wire [WIDTH*2-1+2:0] tmp02_4_23;
	wire [WIDTH*2-1+2:0] tmp02_4_24;
	wire [WIDTH*2-1+2:0] tmp02_4_25;
	wire [WIDTH*2-1+2:0] tmp02_4_26;
	wire [WIDTH*2-1+2:0] tmp02_4_27;
	wire [WIDTH*2-1+2:0] tmp02_4_28;
	wire [WIDTH*2-1+2:0] tmp02_4_29;
	wire [WIDTH*2-1+2:0] tmp02_4_30;
	wire [WIDTH*2-1+2:0] tmp02_4_31;
	wire [WIDTH*2-1+2:0] tmp02_4_32;
	wire [WIDTH*2-1+2:0] tmp02_4_33;
	wire [WIDTH*2-1+2:0] tmp02_4_34;
	wire [WIDTH*2-1+2:0] tmp02_4_35;
	wire [WIDTH*2-1+2:0] tmp02_4_36;
	wire [WIDTH*2-1+2:0] tmp02_4_37;
	wire [WIDTH*2-1+2:0] tmp02_4_38;
	wire [WIDTH*2-1+2:0] tmp02_4_39;
	wire [WIDTH*2-1+2:0] tmp02_4_40;
	wire [WIDTH*2-1+2:0] tmp02_4_41;
	wire [WIDTH*2-1+2:0] tmp02_4_42;
	wire [WIDTH*2-1+2:0] tmp02_4_43;
	wire [WIDTH*2-1+2:0] tmp02_4_44;
	wire [WIDTH*2-1+2:0] tmp02_4_45;
	wire [WIDTH*2-1+2:0] tmp02_4_46;
	wire [WIDTH*2-1+2:0] tmp02_4_47;
	wire [WIDTH*2-1+2:0] tmp02_4_48;
	wire [WIDTH*2-1+2:0] tmp02_4_49;
	wire [WIDTH*2-1+2:0] tmp02_4_50;
	wire [WIDTH*2-1+2:0] tmp02_4_51;
	wire [WIDTH*2-1+2:0] tmp02_4_52;
	wire [WIDTH*2-1+2:0] tmp02_4_53;
	wire [WIDTH*2-1+2:0] tmp02_4_54;
	wire [WIDTH*2-1+2:0] tmp02_4_55;
	wire [WIDTH*2-1+2:0] tmp02_4_56;
	wire [WIDTH*2-1+2:0] tmp02_4_57;
	wire [WIDTH*2-1+2:0] tmp02_4_58;
	wire [WIDTH*2-1+2:0] tmp02_4_59;
	wire [WIDTH*2-1+2:0] tmp02_4_60;
	wire [WIDTH*2-1+2:0] tmp02_4_61;
	wire [WIDTH*2-1+2:0] tmp02_4_62;
	wire [WIDTH*2-1+2:0] tmp02_4_63;
	wire [WIDTH*2-1+2:0] tmp02_4_64;
	wire [WIDTH*2-1+2:0] tmp02_4_65;
	wire [WIDTH*2-1+2:0] tmp02_4_66;
	wire [WIDTH*2-1+2:0] tmp02_4_67;
	wire [WIDTH*2-1+2:0] tmp02_4_68;
	wire [WIDTH*2-1+2:0] tmp02_4_69;
	wire [WIDTH*2-1+2:0] tmp02_4_70;
	wire [WIDTH*2-1+2:0] tmp02_4_71;
	wire [WIDTH*2-1+2:0] tmp02_4_72;
	wire [WIDTH*2-1+2:0] tmp02_4_73;
	wire [WIDTH*2-1+2:0] tmp02_4_74;
	wire [WIDTH*2-1+2:0] tmp02_4_75;
	wire [WIDTH*2-1+2:0] tmp02_4_76;
	wire [WIDTH*2-1+2:0] tmp02_4_77;
	wire [WIDTH*2-1+2:0] tmp02_4_78;
	wire [WIDTH*2-1+2:0] tmp02_4_79;
	wire [WIDTH*2-1+2:0] tmp02_4_80;
	wire [WIDTH*2-1+2:0] tmp02_4_81;
	wire [WIDTH*2-1+2:0] tmp02_4_82;
	wire [WIDTH*2-1+2:0] tmp02_4_83;
	wire [WIDTH*2-1+2:0] tmp02_5_0;
	wire [WIDTH*2-1+2:0] tmp02_5_1;
	wire [WIDTH*2-1+2:0] tmp02_5_2;
	wire [WIDTH*2-1+2:0] tmp02_5_3;
	wire [WIDTH*2-1+2:0] tmp02_5_4;
	wire [WIDTH*2-1+2:0] tmp02_5_5;
	wire [WIDTH*2-1+2:0] tmp02_5_6;
	wire [WIDTH*2-1+2:0] tmp02_5_7;
	wire [WIDTH*2-1+2:0] tmp02_5_8;
	wire [WIDTH*2-1+2:0] tmp02_5_9;
	wire [WIDTH*2-1+2:0] tmp02_5_10;
	wire [WIDTH*2-1+2:0] tmp02_5_11;
	wire [WIDTH*2-1+2:0] tmp02_5_12;
	wire [WIDTH*2-1+2:0] tmp02_5_13;
	wire [WIDTH*2-1+2:0] tmp02_5_14;
	wire [WIDTH*2-1+2:0] tmp02_5_15;
	wire [WIDTH*2-1+2:0] tmp02_5_16;
	wire [WIDTH*2-1+2:0] tmp02_5_17;
	wire [WIDTH*2-1+2:0] tmp02_5_18;
	wire [WIDTH*2-1+2:0] tmp02_5_19;
	wire [WIDTH*2-1+2:0] tmp02_5_20;
	wire [WIDTH*2-1+2:0] tmp02_5_21;
	wire [WIDTH*2-1+2:0] tmp02_5_22;
	wire [WIDTH*2-1+2:0] tmp02_5_23;
	wire [WIDTH*2-1+2:0] tmp02_5_24;
	wire [WIDTH*2-1+2:0] tmp02_5_25;
	wire [WIDTH*2-1+2:0] tmp02_5_26;
	wire [WIDTH*2-1+2:0] tmp02_5_27;
	wire [WIDTH*2-1+2:0] tmp02_5_28;
	wire [WIDTH*2-1+2:0] tmp02_5_29;
	wire [WIDTH*2-1+2:0] tmp02_5_30;
	wire [WIDTH*2-1+2:0] tmp02_5_31;
	wire [WIDTH*2-1+2:0] tmp02_5_32;
	wire [WIDTH*2-1+2:0] tmp02_5_33;
	wire [WIDTH*2-1+2:0] tmp02_5_34;
	wire [WIDTH*2-1+2:0] tmp02_5_35;
	wire [WIDTH*2-1+2:0] tmp02_5_36;
	wire [WIDTH*2-1+2:0] tmp02_5_37;
	wire [WIDTH*2-1+2:0] tmp02_5_38;
	wire [WIDTH*2-1+2:0] tmp02_5_39;
	wire [WIDTH*2-1+2:0] tmp02_5_40;
	wire [WIDTH*2-1+2:0] tmp02_5_41;
	wire [WIDTH*2-1+2:0] tmp02_5_42;
	wire [WIDTH*2-1+2:0] tmp02_5_43;
	wire [WIDTH*2-1+2:0] tmp02_5_44;
	wire [WIDTH*2-1+2:0] tmp02_5_45;
	wire [WIDTH*2-1+2:0] tmp02_5_46;
	wire [WIDTH*2-1+2:0] tmp02_5_47;
	wire [WIDTH*2-1+2:0] tmp02_5_48;
	wire [WIDTH*2-1+2:0] tmp02_5_49;
	wire [WIDTH*2-1+2:0] tmp02_5_50;
	wire [WIDTH*2-1+2:0] tmp02_5_51;
	wire [WIDTH*2-1+2:0] tmp02_5_52;
	wire [WIDTH*2-1+2:0] tmp02_5_53;
	wire [WIDTH*2-1+2:0] tmp02_5_54;
	wire [WIDTH*2-1+2:0] tmp02_5_55;
	wire [WIDTH*2-1+2:0] tmp02_5_56;
	wire [WIDTH*2-1+2:0] tmp02_5_57;
	wire [WIDTH*2-1+2:0] tmp02_5_58;
	wire [WIDTH*2-1+2:0] tmp02_5_59;
	wire [WIDTH*2-1+2:0] tmp02_5_60;
	wire [WIDTH*2-1+2:0] tmp02_5_61;
	wire [WIDTH*2-1+2:0] tmp02_5_62;
	wire [WIDTH*2-1+2:0] tmp02_5_63;
	wire [WIDTH*2-1+2:0] tmp02_5_64;
	wire [WIDTH*2-1+2:0] tmp02_5_65;
	wire [WIDTH*2-1+2:0] tmp02_5_66;
	wire [WIDTH*2-1+2:0] tmp02_5_67;
	wire [WIDTH*2-1+2:0] tmp02_5_68;
	wire [WIDTH*2-1+2:0] tmp02_5_69;
	wire [WIDTH*2-1+2:0] tmp02_5_70;
	wire [WIDTH*2-1+2:0] tmp02_5_71;
	wire [WIDTH*2-1+2:0] tmp02_5_72;
	wire [WIDTH*2-1+2:0] tmp02_5_73;
	wire [WIDTH*2-1+2:0] tmp02_5_74;
	wire [WIDTH*2-1+2:0] tmp02_5_75;
	wire [WIDTH*2-1+2:0] tmp02_5_76;
	wire [WIDTH*2-1+2:0] tmp02_5_77;
	wire [WIDTH*2-1+2:0] tmp02_5_78;
	wire [WIDTH*2-1+2:0] tmp02_5_79;
	wire [WIDTH*2-1+2:0] tmp02_5_80;
	wire [WIDTH*2-1+2:0] tmp02_5_81;
	wire [WIDTH*2-1+2:0] tmp02_5_82;
	wire [WIDTH*2-1+2:0] tmp02_5_83;
	wire [WIDTH*2-1+2:0] tmp02_6_0;
	wire [WIDTH*2-1+2:0] tmp02_6_1;
	wire [WIDTH*2-1+2:0] tmp02_6_2;
	wire [WIDTH*2-1+2:0] tmp02_6_3;
	wire [WIDTH*2-1+2:0] tmp02_6_4;
	wire [WIDTH*2-1+2:0] tmp02_6_5;
	wire [WIDTH*2-1+2:0] tmp02_6_6;
	wire [WIDTH*2-1+2:0] tmp02_6_7;
	wire [WIDTH*2-1+2:0] tmp02_6_8;
	wire [WIDTH*2-1+2:0] tmp02_6_9;
	wire [WIDTH*2-1+2:0] tmp02_6_10;
	wire [WIDTH*2-1+2:0] tmp02_6_11;
	wire [WIDTH*2-1+2:0] tmp02_6_12;
	wire [WIDTH*2-1+2:0] tmp02_6_13;
	wire [WIDTH*2-1+2:0] tmp02_6_14;
	wire [WIDTH*2-1+2:0] tmp02_6_15;
	wire [WIDTH*2-1+2:0] tmp02_6_16;
	wire [WIDTH*2-1+2:0] tmp02_6_17;
	wire [WIDTH*2-1+2:0] tmp02_6_18;
	wire [WIDTH*2-1+2:0] tmp02_6_19;
	wire [WIDTH*2-1+2:0] tmp02_6_20;
	wire [WIDTH*2-1+2:0] tmp02_6_21;
	wire [WIDTH*2-1+2:0] tmp02_6_22;
	wire [WIDTH*2-1+2:0] tmp02_6_23;
	wire [WIDTH*2-1+2:0] tmp02_6_24;
	wire [WIDTH*2-1+2:0] tmp02_6_25;
	wire [WIDTH*2-1+2:0] tmp02_6_26;
	wire [WIDTH*2-1+2:0] tmp02_6_27;
	wire [WIDTH*2-1+2:0] tmp02_6_28;
	wire [WIDTH*2-1+2:0] tmp02_6_29;
	wire [WIDTH*2-1+2:0] tmp02_6_30;
	wire [WIDTH*2-1+2:0] tmp02_6_31;
	wire [WIDTH*2-1+2:0] tmp02_6_32;
	wire [WIDTH*2-1+2:0] tmp02_6_33;
	wire [WIDTH*2-1+2:0] tmp02_6_34;
	wire [WIDTH*2-1+2:0] tmp02_6_35;
	wire [WIDTH*2-1+2:0] tmp02_6_36;
	wire [WIDTH*2-1+2:0] tmp02_6_37;
	wire [WIDTH*2-1+2:0] tmp02_6_38;
	wire [WIDTH*2-1+2:0] tmp02_6_39;
	wire [WIDTH*2-1+2:0] tmp02_6_40;
	wire [WIDTH*2-1+2:0] tmp02_6_41;
	wire [WIDTH*2-1+2:0] tmp02_6_42;
	wire [WIDTH*2-1+2:0] tmp02_6_43;
	wire [WIDTH*2-1+2:0] tmp02_6_44;
	wire [WIDTH*2-1+2:0] tmp02_6_45;
	wire [WIDTH*2-1+2:0] tmp02_6_46;
	wire [WIDTH*2-1+2:0] tmp02_6_47;
	wire [WIDTH*2-1+2:0] tmp02_6_48;
	wire [WIDTH*2-1+2:0] tmp02_6_49;
	wire [WIDTH*2-1+2:0] tmp02_6_50;
	wire [WIDTH*2-1+2:0] tmp02_6_51;
	wire [WIDTH*2-1+2:0] tmp02_6_52;
	wire [WIDTH*2-1+2:0] tmp02_6_53;
	wire [WIDTH*2-1+2:0] tmp02_6_54;
	wire [WIDTH*2-1+2:0] tmp02_6_55;
	wire [WIDTH*2-1+2:0] tmp02_6_56;
	wire [WIDTH*2-1+2:0] tmp02_6_57;
	wire [WIDTH*2-1+2:0] tmp02_6_58;
	wire [WIDTH*2-1+2:0] tmp02_6_59;
	wire [WIDTH*2-1+2:0] tmp02_6_60;
	wire [WIDTH*2-1+2:0] tmp02_6_61;
	wire [WIDTH*2-1+2:0] tmp02_6_62;
	wire [WIDTH*2-1+2:0] tmp02_6_63;
	wire [WIDTH*2-1+2:0] tmp02_6_64;
	wire [WIDTH*2-1+2:0] tmp02_6_65;
	wire [WIDTH*2-1+2:0] tmp02_6_66;
	wire [WIDTH*2-1+2:0] tmp02_6_67;
	wire [WIDTH*2-1+2:0] tmp02_6_68;
	wire [WIDTH*2-1+2:0] tmp02_6_69;
	wire [WIDTH*2-1+2:0] tmp02_6_70;
	wire [WIDTH*2-1+2:0] tmp02_6_71;
	wire [WIDTH*2-1+2:0] tmp02_6_72;
	wire [WIDTH*2-1+2:0] tmp02_6_73;
	wire [WIDTH*2-1+2:0] tmp02_6_74;
	wire [WIDTH*2-1+2:0] tmp02_6_75;
	wire [WIDTH*2-1+2:0] tmp02_6_76;
	wire [WIDTH*2-1+2:0] tmp02_6_77;
	wire [WIDTH*2-1+2:0] tmp02_6_78;
	wire [WIDTH*2-1+2:0] tmp02_6_79;
	wire [WIDTH*2-1+2:0] tmp02_6_80;
	wire [WIDTH*2-1+2:0] tmp02_6_81;
	wire [WIDTH*2-1+2:0] tmp02_6_82;
	wire [WIDTH*2-1+2:0] tmp02_6_83;
	wire [WIDTH*2-1+2:0] tmp02_7_0;
	wire [WIDTH*2-1+2:0] tmp02_7_1;
	wire [WIDTH*2-1+2:0] tmp02_7_2;
	wire [WIDTH*2-1+2:0] tmp02_7_3;
	wire [WIDTH*2-1+2:0] tmp02_7_4;
	wire [WIDTH*2-1+2:0] tmp02_7_5;
	wire [WIDTH*2-1+2:0] tmp02_7_6;
	wire [WIDTH*2-1+2:0] tmp02_7_7;
	wire [WIDTH*2-1+2:0] tmp02_7_8;
	wire [WIDTH*2-1+2:0] tmp02_7_9;
	wire [WIDTH*2-1+2:0] tmp02_7_10;
	wire [WIDTH*2-1+2:0] tmp02_7_11;
	wire [WIDTH*2-1+2:0] tmp02_7_12;
	wire [WIDTH*2-1+2:0] tmp02_7_13;
	wire [WIDTH*2-1+2:0] tmp02_7_14;
	wire [WIDTH*2-1+2:0] tmp02_7_15;
	wire [WIDTH*2-1+2:0] tmp02_7_16;
	wire [WIDTH*2-1+2:0] tmp02_7_17;
	wire [WIDTH*2-1+2:0] tmp02_7_18;
	wire [WIDTH*2-1+2:0] tmp02_7_19;
	wire [WIDTH*2-1+2:0] tmp02_7_20;
	wire [WIDTH*2-1+2:0] tmp02_7_21;
	wire [WIDTH*2-1+2:0] tmp02_7_22;
	wire [WIDTH*2-1+2:0] tmp02_7_23;
	wire [WIDTH*2-1+2:0] tmp02_7_24;
	wire [WIDTH*2-1+2:0] tmp02_7_25;
	wire [WIDTH*2-1+2:0] tmp02_7_26;
	wire [WIDTH*2-1+2:0] tmp02_7_27;
	wire [WIDTH*2-1+2:0] tmp02_7_28;
	wire [WIDTH*2-1+2:0] tmp02_7_29;
	wire [WIDTH*2-1+2:0] tmp02_7_30;
	wire [WIDTH*2-1+2:0] tmp02_7_31;
	wire [WIDTH*2-1+2:0] tmp02_7_32;
	wire [WIDTH*2-1+2:0] tmp02_7_33;
	wire [WIDTH*2-1+2:0] tmp02_7_34;
	wire [WIDTH*2-1+2:0] tmp02_7_35;
	wire [WIDTH*2-1+2:0] tmp02_7_36;
	wire [WIDTH*2-1+2:0] tmp02_7_37;
	wire [WIDTH*2-1+2:0] tmp02_7_38;
	wire [WIDTH*2-1+2:0] tmp02_7_39;
	wire [WIDTH*2-1+2:0] tmp02_7_40;
	wire [WIDTH*2-1+2:0] tmp02_7_41;
	wire [WIDTH*2-1+2:0] tmp02_7_42;
	wire [WIDTH*2-1+2:0] tmp02_7_43;
	wire [WIDTH*2-1+2:0] tmp02_7_44;
	wire [WIDTH*2-1+2:0] tmp02_7_45;
	wire [WIDTH*2-1+2:0] tmp02_7_46;
	wire [WIDTH*2-1+2:0] tmp02_7_47;
	wire [WIDTH*2-1+2:0] tmp02_7_48;
	wire [WIDTH*2-1+2:0] tmp02_7_49;
	wire [WIDTH*2-1+2:0] tmp02_7_50;
	wire [WIDTH*2-1+2:0] tmp02_7_51;
	wire [WIDTH*2-1+2:0] tmp02_7_52;
	wire [WIDTH*2-1+2:0] tmp02_7_53;
	wire [WIDTH*2-1+2:0] tmp02_7_54;
	wire [WIDTH*2-1+2:0] tmp02_7_55;
	wire [WIDTH*2-1+2:0] tmp02_7_56;
	wire [WIDTH*2-1+2:0] tmp02_7_57;
	wire [WIDTH*2-1+2:0] tmp02_7_58;
	wire [WIDTH*2-1+2:0] tmp02_7_59;
	wire [WIDTH*2-1+2:0] tmp02_7_60;
	wire [WIDTH*2-1+2:0] tmp02_7_61;
	wire [WIDTH*2-1+2:0] tmp02_7_62;
	wire [WIDTH*2-1+2:0] tmp02_7_63;
	wire [WIDTH*2-1+2:0] tmp02_7_64;
	wire [WIDTH*2-1+2:0] tmp02_7_65;
	wire [WIDTH*2-1+2:0] tmp02_7_66;
	wire [WIDTH*2-1+2:0] tmp02_7_67;
	wire [WIDTH*2-1+2:0] tmp02_7_68;
	wire [WIDTH*2-1+2:0] tmp02_7_69;
	wire [WIDTH*2-1+2:0] tmp02_7_70;
	wire [WIDTH*2-1+2:0] tmp02_7_71;
	wire [WIDTH*2-1+2:0] tmp02_7_72;
	wire [WIDTH*2-1+2:0] tmp02_7_73;
	wire [WIDTH*2-1+2:0] tmp02_7_74;
	wire [WIDTH*2-1+2:0] tmp02_7_75;
	wire [WIDTH*2-1+2:0] tmp02_7_76;
	wire [WIDTH*2-1+2:0] tmp02_7_77;
	wire [WIDTH*2-1+2:0] tmp02_7_78;
	wire [WIDTH*2-1+2:0] tmp02_7_79;
	wire [WIDTH*2-1+2:0] tmp02_7_80;
	wire [WIDTH*2-1+2:0] tmp02_7_81;
	wire [WIDTH*2-1+2:0] tmp02_7_82;
	wire [WIDTH*2-1+2:0] tmp02_7_83;
	wire [WIDTH*2-1+2:0] tmp02_8_0;
	wire [WIDTH*2-1+2:0] tmp02_8_1;
	wire [WIDTH*2-1+2:0] tmp02_8_2;
	wire [WIDTH*2-1+2:0] tmp02_8_3;
	wire [WIDTH*2-1+2:0] tmp02_8_4;
	wire [WIDTH*2-1+2:0] tmp02_8_5;
	wire [WIDTH*2-1+2:0] tmp02_8_6;
	wire [WIDTH*2-1+2:0] tmp02_8_7;
	wire [WIDTH*2-1+2:0] tmp02_8_8;
	wire [WIDTH*2-1+2:0] tmp02_8_9;
	wire [WIDTH*2-1+2:0] tmp02_8_10;
	wire [WIDTH*2-1+2:0] tmp02_8_11;
	wire [WIDTH*2-1+2:0] tmp02_8_12;
	wire [WIDTH*2-1+2:0] tmp02_8_13;
	wire [WIDTH*2-1+2:0] tmp02_8_14;
	wire [WIDTH*2-1+2:0] tmp02_8_15;
	wire [WIDTH*2-1+2:0] tmp02_8_16;
	wire [WIDTH*2-1+2:0] tmp02_8_17;
	wire [WIDTH*2-1+2:0] tmp02_8_18;
	wire [WIDTH*2-1+2:0] tmp02_8_19;
	wire [WIDTH*2-1+2:0] tmp02_8_20;
	wire [WIDTH*2-1+2:0] tmp02_8_21;
	wire [WIDTH*2-1+2:0] tmp02_8_22;
	wire [WIDTH*2-1+2:0] tmp02_8_23;
	wire [WIDTH*2-1+2:0] tmp02_8_24;
	wire [WIDTH*2-1+2:0] tmp02_8_25;
	wire [WIDTH*2-1+2:0] tmp02_8_26;
	wire [WIDTH*2-1+2:0] tmp02_8_27;
	wire [WIDTH*2-1+2:0] tmp02_8_28;
	wire [WIDTH*2-1+2:0] tmp02_8_29;
	wire [WIDTH*2-1+2:0] tmp02_8_30;
	wire [WIDTH*2-1+2:0] tmp02_8_31;
	wire [WIDTH*2-1+2:0] tmp02_8_32;
	wire [WIDTH*2-1+2:0] tmp02_8_33;
	wire [WIDTH*2-1+2:0] tmp02_8_34;
	wire [WIDTH*2-1+2:0] tmp02_8_35;
	wire [WIDTH*2-1+2:0] tmp02_8_36;
	wire [WIDTH*2-1+2:0] tmp02_8_37;
	wire [WIDTH*2-1+2:0] tmp02_8_38;
	wire [WIDTH*2-1+2:0] tmp02_8_39;
	wire [WIDTH*2-1+2:0] tmp02_8_40;
	wire [WIDTH*2-1+2:0] tmp02_8_41;
	wire [WIDTH*2-1+2:0] tmp02_8_42;
	wire [WIDTH*2-1+2:0] tmp02_8_43;
	wire [WIDTH*2-1+2:0] tmp02_8_44;
	wire [WIDTH*2-1+2:0] tmp02_8_45;
	wire [WIDTH*2-1+2:0] tmp02_8_46;
	wire [WIDTH*2-1+2:0] tmp02_8_47;
	wire [WIDTH*2-1+2:0] tmp02_8_48;
	wire [WIDTH*2-1+2:0] tmp02_8_49;
	wire [WIDTH*2-1+2:0] tmp02_8_50;
	wire [WIDTH*2-1+2:0] tmp02_8_51;
	wire [WIDTH*2-1+2:0] tmp02_8_52;
	wire [WIDTH*2-1+2:0] tmp02_8_53;
	wire [WIDTH*2-1+2:0] tmp02_8_54;
	wire [WIDTH*2-1+2:0] tmp02_8_55;
	wire [WIDTH*2-1+2:0] tmp02_8_56;
	wire [WIDTH*2-1+2:0] tmp02_8_57;
	wire [WIDTH*2-1+2:0] tmp02_8_58;
	wire [WIDTH*2-1+2:0] tmp02_8_59;
	wire [WIDTH*2-1+2:0] tmp02_8_60;
	wire [WIDTH*2-1+2:0] tmp02_8_61;
	wire [WIDTH*2-1+2:0] tmp02_8_62;
	wire [WIDTH*2-1+2:0] tmp02_8_63;
	wire [WIDTH*2-1+2:0] tmp02_8_64;
	wire [WIDTH*2-1+2:0] tmp02_8_65;
	wire [WIDTH*2-1+2:0] tmp02_8_66;
	wire [WIDTH*2-1+2:0] tmp02_8_67;
	wire [WIDTH*2-1+2:0] tmp02_8_68;
	wire [WIDTH*2-1+2:0] tmp02_8_69;
	wire [WIDTH*2-1+2:0] tmp02_8_70;
	wire [WIDTH*2-1+2:0] tmp02_8_71;
	wire [WIDTH*2-1+2:0] tmp02_8_72;
	wire [WIDTH*2-1+2:0] tmp02_8_73;
	wire [WIDTH*2-1+2:0] tmp02_8_74;
	wire [WIDTH*2-1+2:0] tmp02_8_75;
	wire [WIDTH*2-1+2:0] tmp02_8_76;
	wire [WIDTH*2-1+2:0] tmp02_8_77;
	wire [WIDTH*2-1+2:0] tmp02_8_78;
	wire [WIDTH*2-1+2:0] tmp02_8_79;
	wire [WIDTH*2-1+2:0] tmp02_8_80;
	wire [WIDTH*2-1+2:0] tmp02_8_81;
	wire [WIDTH*2-1+2:0] tmp02_8_82;
	wire [WIDTH*2-1+2:0] tmp02_8_83;
	wire [WIDTH*2-1+2:0] tmp02_9_0;
	wire [WIDTH*2-1+2:0] tmp02_9_1;
	wire [WIDTH*2-1+2:0] tmp02_9_2;
	wire [WIDTH*2-1+2:0] tmp02_9_3;
	wire [WIDTH*2-1+2:0] tmp02_9_4;
	wire [WIDTH*2-1+2:0] tmp02_9_5;
	wire [WIDTH*2-1+2:0] tmp02_9_6;
	wire [WIDTH*2-1+2:0] tmp02_9_7;
	wire [WIDTH*2-1+2:0] tmp02_9_8;
	wire [WIDTH*2-1+2:0] tmp02_9_9;
	wire [WIDTH*2-1+2:0] tmp02_9_10;
	wire [WIDTH*2-1+2:0] tmp02_9_11;
	wire [WIDTH*2-1+2:0] tmp02_9_12;
	wire [WIDTH*2-1+2:0] tmp02_9_13;
	wire [WIDTH*2-1+2:0] tmp02_9_14;
	wire [WIDTH*2-1+2:0] tmp02_9_15;
	wire [WIDTH*2-1+2:0] tmp02_9_16;
	wire [WIDTH*2-1+2:0] tmp02_9_17;
	wire [WIDTH*2-1+2:0] tmp02_9_18;
	wire [WIDTH*2-1+2:0] tmp02_9_19;
	wire [WIDTH*2-1+2:0] tmp02_9_20;
	wire [WIDTH*2-1+2:0] tmp02_9_21;
	wire [WIDTH*2-1+2:0] tmp02_9_22;
	wire [WIDTH*2-1+2:0] tmp02_9_23;
	wire [WIDTH*2-1+2:0] tmp02_9_24;
	wire [WIDTH*2-1+2:0] tmp02_9_25;
	wire [WIDTH*2-1+2:0] tmp02_9_26;
	wire [WIDTH*2-1+2:0] tmp02_9_27;
	wire [WIDTH*2-1+2:0] tmp02_9_28;
	wire [WIDTH*2-1+2:0] tmp02_9_29;
	wire [WIDTH*2-1+2:0] tmp02_9_30;
	wire [WIDTH*2-1+2:0] tmp02_9_31;
	wire [WIDTH*2-1+2:0] tmp02_9_32;
	wire [WIDTH*2-1+2:0] tmp02_9_33;
	wire [WIDTH*2-1+2:0] tmp02_9_34;
	wire [WIDTH*2-1+2:0] tmp02_9_35;
	wire [WIDTH*2-1+2:0] tmp02_9_36;
	wire [WIDTH*2-1+2:0] tmp02_9_37;
	wire [WIDTH*2-1+2:0] tmp02_9_38;
	wire [WIDTH*2-1+2:0] tmp02_9_39;
	wire [WIDTH*2-1+2:0] tmp02_9_40;
	wire [WIDTH*2-1+2:0] tmp02_9_41;
	wire [WIDTH*2-1+2:0] tmp02_9_42;
	wire [WIDTH*2-1+2:0] tmp02_9_43;
	wire [WIDTH*2-1+2:0] tmp02_9_44;
	wire [WIDTH*2-1+2:0] tmp02_9_45;
	wire [WIDTH*2-1+2:0] tmp02_9_46;
	wire [WIDTH*2-1+2:0] tmp02_9_47;
	wire [WIDTH*2-1+2:0] tmp02_9_48;
	wire [WIDTH*2-1+2:0] tmp02_9_49;
	wire [WIDTH*2-1+2:0] tmp02_9_50;
	wire [WIDTH*2-1+2:0] tmp02_9_51;
	wire [WIDTH*2-1+2:0] tmp02_9_52;
	wire [WIDTH*2-1+2:0] tmp02_9_53;
	wire [WIDTH*2-1+2:0] tmp02_9_54;
	wire [WIDTH*2-1+2:0] tmp02_9_55;
	wire [WIDTH*2-1+2:0] tmp02_9_56;
	wire [WIDTH*2-1+2:0] tmp02_9_57;
	wire [WIDTH*2-1+2:0] tmp02_9_58;
	wire [WIDTH*2-1+2:0] tmp02_9_59;
	wire [WIDTH*2-1+2:0] tmp02_9_60;
	wire [WIDTH*2-1+2:0] tmp02_9_61;
	wire [WIDTH*2-1+2:0] tmp02_9_62;
	wire [WIDTH*2-1+2:0] tmp02_9_63;
	wire [WIDTH*2-1+2:0] tmp02_9_64;
	wire [WIDTH*2-1+2:0] tmp02_9_65;
	wire [WIDTH*2-1+2:0] tmp02_9_66;
	wire [WIDTH*2-1+2:0] tmp02_9_67;
	wire [WIDTH*2-1+2:0] tmp02_9_68;
	wire [WIDTH*2-1+2:0] tmp02_9_69;
	wire [WIDTH*2-1+2:0] tmp02_9_70;
	wire [WIDTH*2-1+2:0] tmp02_9_71;
	wire [WIDTH*2-1+2:0] tmp02_9_72;
	wire [WIDTH*2-1+2:0] tmp02_9_73;
	wire [WIDTH*2-1+2:0] tmp02_9_74;
	wire [WIDTH*2-1+2:0] tmp02_9_75;
	wire [WIDTH*2-1+2:0] tmp02_9_76;
	wire [WIDTH*2-1+2:0] tmp02_9_77;
	wire [WIDTH*2-1+2:0] tmp02_9_78;
	wire [WIDTH*2-1+2:0] tmp02_9_79;
	wire [WIDTH*2-1+2:0] tmp02_9_80;
	wire [WIDTH*2-1+2:0] tmp02_9_81;
	wire [WIDTH*2-1+2:0] tmp02_9_82;
	wire [WIDTH*2-1+2:0] tmp02_9_83;
	wire [WIDTH*2-1+2:0] tmp02_10_0;
	wire [WIDTH*2-1+2:0] tmp02_10_1;
	wire [WIDTH*2-1+2:0] tmp02_10_2;
	wire [WIDTH*2-1+2:0] tmp02_10_3;
	wire [WIDTH*2-1+2:0] tmp02_10_4;
	wire [WIDTH*2-1+2:0] tmp02_10_5;
	wire [WIDTH*2-1+2:0] tmp02_10_6;
	wire [WIDTH*2-1+2:0] tmp02_10_7;
	wire [WIDTH*2-1+2:0] tmp02_10_8;
	wire [WIDTH*2-1+2:0] tmp02_10_9;
	wire [WIDTH*2-1+2:0] tmp02_10_10;
	wire [WIDTH*2-1+2:0] tmp02_10_11;
	wire [WIDTH*2-1+2:0] tmp02_10_12;
	wire [WIDTH*2-1+2:0] tmp02_10_13;
	wire [WIDTH*2-1+2:0] tmp02_10_14;
	wire [WIDTH*2-1+2:0] tmp02_10_15;
	wire [WIDTH*2-1+2:0] tmp02_10_16;
	wire [WIDTH*2-1+2:0] tmp02_10_17;
	wire [WIDTH*2-1+2:0] tmp02_10_18;
	wire [WIDTH*2-1+2:0] tmp02_10_19;
	wire [WIDTH*2-1+2:0] tmp02_10_20;
	wire [WIDTH*2-1+2:0] tmp02_10_21;
	wire [WIDTH*2-1+2:0] tmp02_10_22;
	wire [WIDTH*2-1+2:0] tmp02_10_23;
	wire [WIDTH*2-1+2:0] tmp02_10_24;
	wire [WIDTH*2-1+2:0] tmp02_10_25;
	wire [WIDTH*2-1+2:0] tmp02_10_26;
	wire [WIDTH*2-1+2:0] tmp02_10_27;
	wire [WIDTH*2-1+2:0] tmp02_10_28;
	wire [WIDTH*2-1+2:0] tmp02_10_29;
	wire [WIDTH*2-1+2:0] tmp02_10_30;
	wire [WIDTH*2-1+2:0] tmp02_10_31;
	wire [WIDTH*2-1+2:0] tmp02_10_32;
	wire [WIDTH*2-1+2:0] tmp02_10_33;
	wire [WIDTH*2-1+2:0] tmp02_10_34;
	wire [WIDTH*2-1+2:0] tmp02_10_35;
	wire [WIDTH*2-1+2:0] tmp02_10_36;
	wire [WIDTH*2-1+2:0] tmp02_10_37;
	wire [WIDTH*2-1+2:0] tmp02_10_38;
	wire [WIDTH*2-1+2:0] tmp02_10_39;
	wire [WIDTH*2-1+2:0] tmp02_10_40;
	wire [WIDTH*2-1+2:0] tmp02_10_41;
	wire [WIDTH*2-1+2:0] tmp02_10_42;
	wire [WIDTH*2-1+2:0] tmp02_10_43;
	wire [WIDTH*2-1+2:0] tmp02_10_44;
	wire [WIDTH*2-1+2:0] tmp02_10_45;
	wire [WIDTH*2-1+2:0] tmp02_10_46;
	wire [WIDTH*2-1+2:0] tmp02_10_47;
	wire [WIDTH*2-1+2:0] tmp02_10_48;
	wire [WIDTH*2-1+2:0] tmp02_10_49;
	wire [WIDTH*2-1+2:0] tmp02_10_50;
	wire [WIDTH*2-1+2:0] tmp02_10_51;
	wire [WIDTH*2-1+2:0] tmp02_10_52;
	wire [WIDTH*2-1+2:0] tmp02_10_53;
	wire [WIDTH*2-1+2:0] tmp02_10_54;
	wire [WIDTH*2-1+2:0] tmp02_10_55;
	wire [WIDTH*2-1+2:0] tmp02_10_56;
	wire [WIDTH*2-1+2:0] tmp02_10_57;
	wire [WIDTH*2-1+2:0] tmp02_10_58;
	wire [WIDTH*2-1+2:0] tmp02_10_59;
	wire [WIDTH*2-1+2:0] tmp02_10_60;
	wire [WIDTH*2-1+2:0] tmp02_10_61;
	wire [WIDTH*2-1+2:0] tmp02_10_62;
	wire [WIDTH*2-1+2:0] tmp02_10_63;
	wire [WIDTH*2-1+2:0] tmp02_10_64;
	wire [WIDTH*2-1+2:0] tmp02_10_65;
	wire [WIDTH*2-1+2:0] tmp02_10_66;
	wire [WIDTH*2-1+2:0] tmp02_10_67;
	wire [WIDTH*2-1+2:0] tmp02_10_68;
	wire [WIDTH*2-1+2:0] tmp02_10_69;
	wire [WIDTH*2-1+2:0] tmp02_10_70;
	wire [WIDTH*2-1+2:0] tmp02_10_71;
	wire [WIDTH*2-1+2:0] tmp02_10_72;
	wire [WIDTH*2-1+2:0] tmp02_10_73;
	wire [WIDTH*2-1+2:0] tmp02_10_74;
	wire [WIDTH*2-1+2:0] tmp02_10_75;
	wire [WIDTH*2-1+2:0] tmp02_10_76;
	wire [WIDTH*2-1+2:0] tmp02_10_77;
	wire [WIDTH*2-1+2:0] tmp02_10_78;
	wire [WIDTH*2-1+2:0] tmp02_10_79;
	wire [WIDTH*2-1+2:0] tmp02_10_80;
	wire [WIDTH*2-1+2:0] tmp02_10_81;
	wire [WIDTH*2-1+2:0] tmp02_10_82;
	wire [WIDTH*2-1+2:0] tmp02_10_83;
	wire [WIDTH*2-1+2:0] tmp02_11_0;
	wire [WIDTH*2-1+2:0] tmp02_11_1;
	wire [WIDTH*2-1+2:0] tmp02_11_2;
	wire [WIDTH*2-1+2:0] tmp02_11_3;
	wire [WIDTH*2-1+2:0] tmp02_11_4;
	wire [WIDTH*2-1+2:0] tmp02_11_5;
	wire [WIDTH*2-1+2:0] tmp02_11_6;
	wire [WIDTH*2-1+2:0] tmp02_11_7;
	wire [WIDTH*2-1+2:0] tmp02_11_8;
	wire [WIDTH*2-1+2:0] tmp02_11_9;
	wire [WIDTH*2-1+2:0] tmp02_11_10;
	wire [WIDTH*2-1+2:0] tmp02_11_11;
	wire [WIDTH*2-1+2:0] tmp02_11_12;
	wire [WIDTH*2-1+2:0] tmp02_11_13;
	wire [WIDTH*2-1+2:0] tmp02_11_14;
	wire [WIDTH*2-1+2:0] tmp02_11_15;
	wire [WIDTH*2-1+2:0] tmp02_11_16;
	wire [WIDTH*2-1+2:0] tmp02_11_17;
	wire [WIDTH*2-1+2:0] tmp02_11_18;
	wire [WIDTH*2-1+2:0] tmp02_11_19;
	wire [WIDTH*2-1+2:0] tmp02_11_20;
	wire [WIDTH*2-1+2:0] tmp02_11_21;
	wire [WIDTH*2-1+2:0] tmp02_11_22;
	wire [WIDTH*2-1+2:0] tmp02_11_23;
	wire [WIDTH*2-1+2:0] tmp02_11_24;
	wire [WIDTH*2-1+2:0] tmp02_11_25;
	wire [WIDTH*2-1+2:0] tmp02_11_26;
	wire [WIDTH*2-1+2:0] tmp02_11_27;
	wire [WIDTH*2-1+2:0] tmp02_11_28;
	wire [WIDTH*2-1+2:0] tmp02_11_29;
	wire [WIDTH*2-1+2:0] tmp02_11_30;
	wire [WIDTH*2-1+2:0] tmp02_11_31;
	wire [WIDTH*2-1+2:0] tmp02_11_32;
	wire [WIDTH*2-1+2:0] tmp02_11_33;
	wire [WIDTH*2-1+2:0] tmp02_11_34;
	wire [WIDTH*2-1+2:0] tmp02_11_35;
	wire [WIDTH*2-1+2:0] tmp02_11_36;
	wire [WIDTH*2-1+2:0] tmp02_11_37;
	wire [WIDTH*2-1+2:0] tmp02_11_38;
	wire [WIDTH*2-1+2:0] tmp02_11_39;
	wire [WIDTH*2-1+2:0] tmp02_11_40;
	wire [WIDTH*2-1+2:0] tmp02_11_41;
	wire [WIDTH*2-1+2:0] tmp02_11_42;
	wire [WIDTH*2-1+2:0] tmp02_11_43;
	wire [WIDTH*2-1+2:0] tmp02_11_44;
	wire [WIDTH*2-1+2:0] tmp02_11_45;
	wire [WIDTH*2-1+2:0] tmp02_11_46;
	wire [WIDTH*2-1+2:0] tmp02_11_47;
	wire [WIDTH*2-1+2:0] tmp02_11_48;
	wire [WIDTH*2-1+2:0] tmp02_11_49;
	wire [WIDTH*2-1+2:0] tmp02_11_50;
	wire [WIDTH*2-1+2:0] tmp02_11_51;
	wire [WIDTH*2-1+2:0] tmp02_11_52;
	wire [WIDTH*2-1+2:0] tmp02_11_53;
	wire [WIDTH*2-1+2:0] tmp02_11_54;
	wire [WIDTH*2-1+2:0] tmp02_11_55;
	wire [WIDTH*2-1+2:0] tmp02_11_56;
	wire [WIDTH*2-1+2:0] tmp02_11_57;
	wire [WIDTH*2-1+2:0] tmp02_11_58;
	wire [WIDTH*2-1+2:0] tmp02_11_59;
	wire [WIDTH*2-1+2:0] tmp02_11_60;
	wire [WIDTH*2-1+2:0] tmp02_11_61;
	wire [WIDTH*2-1+2:0] tmp02_11_62;
	wire [WIDTH*2-1+2:0] tmp02_11_63;
	wire [WIDTH*2-1+2:0] tmp02_11_64;
	wire [WIDTH*2-1+2:0] tmp02_11_65;
	wire [WIDTH*2-1+2:0] tmp02_11_66;
	wire [WIDTH*2-1+2:0] tmp02_11_67;
	wire [WIDTH*2-1+2:0] tmp02_11_68;
	wire [WIDTH*2-1+2:0] tmp02_11_69;
	wire [WIDTH*2-1+2:0] tmp02_11_70;
	wire [WIDTH*2-1+2:0] tmp02_11_71;
	wire [WIDTH*2-1+2:0] tmp02_11_72;
	wire [WIDTH*2-1+2:0] tmp02_11_73;
	wire [WIDTH*2-1+2:0] tmp02_11_74;
	wire [WIDTH*2-1+2:0] tmp02_11_75;
	wire [WIDTH*2-1+2:0] tmp02_11_76;
	wire [WIDTH*2-1+2:0] tmp02_11_77;
	wire [WIDTH*2-1+2:0] tmp02_11_78;
	wire [WIDTH*2-1+2:0] tmp02_11_79;
	wire [WIDTH*2-1+2:0] tmp02_11_80;
	wire [WIDTH*2-1+2:0] tmp02_11_81;
	wire [WIDTH*2-1+2:0] tmp02_11_82;
	wire [WIDTH*2-1+2:0] tmp02_11_83;
	wire [WIDTH*2-1+2:0] tmp02_12_0;
	wire [WIDTH*2-1+2:0] tmp02_12_1;
	wire [WIDTH*2-1+2:0] tmp02_12_2;
	wire [WIDTH*2-1+2:0] tmp02_12_3;
	wire [WIDTH*2-1+2:0] tmp02_12_4;
	wire [WIDTH*2-1+2:0] tmp02_12_5;
	wire [WIDTH*2-1+2:0] tmp02_12_6;
	wire [WIDTH*2-1+2:0] tmp02_12_7;
	wire [WIDTH*2-1+2:0] tmp02_12_8;
	wire [WIDTH*2-1+2:0] tmp02_12_9;
	wire [WIDTH*2-1+2:0] tmp02_12_10;
	wire [WIDTH*2-1+2:0] tmp02_12_11;
	wire [WIDTH*2-1+2:0] tmp02_12_12;
	wire [WIDTH*2-1+2:0] tmp02_12_13;
	wire [WIDTH*2-1+2:0] tmp02_12_14;
	wire [WIDTH*2-1+2:0] tmp02_12_15;
	wire [WIDTH*2-1+2:0] tmp02_12_16;
	wire [WIDTH*2-1+2:0] tmp02_12_17;
	wire [WIDTH*2-1+2:0] tmp02_12_18;
	wire [WIDTH*2-1+2:0] tmp02_12_19;
	wire [WIDTH*2-1+2:0] tmp02_12_20;
	wire [WIDTH*2-1+2:0] tmp02_12_21;
	wire [WIDTH*2-1+2:0] tmp02_12_22;
	wire [WIDTH*2-1+2:0] tmp02_12_23;
	wire [WIDTH*2-1+2:0] tmp02_12_24;
	wire [WIDTH*2-1+2:0] tmp02_12_25;
	wire [WIDTH*2-1+2:0] tmp02_12_26;
	wire [WIDTH*2-1+2:0] tmp02_12_27;
	wire [WIDTH*2-1+2:0] tmp02_12_28;
	wire [WIDTH*2-1+2:0] tmp02_12_29;
	wire [WIDTH*2-1+2:0] tmp02_12_30;
	wire [WIDTH*2-1+2:0] tmp02_12_31;
	wire [WIDTH*2-1+2:0] tmp02_12_32;
	wire [WIDTH*2-1+2:0] tmp02_12_33;
	wire [WIDTH*2-1+2:0] tmp02_12_34;
	wire [WIDTH*2-1+2:0] tmp02_12_35;
	wire [WIDTH*2-1+2:0] tmp02_12_36;
	wire [WIDTH*2-1+2:0] tmp02_12_37;
	wire [WIDTH*2-1+2:0] tmp02_12_38;
	wire [WIDTH*2-1+2:0] tmp02_12_39;
	wire [WIDTH*2-1+2:0] tmp02_12_40;
	wire [WIDTH*2-1+2:0] tmp02_12_41;
	wire [WIDTH*2-1+2:0] tmp02_12_42;
	wire [WIDTH*2-1+2:0] tmp02_12_43;
	wire [WIDTH*2-1+2:0] tmp02_12_44;
	wire [WIDTH*2-1+2:0] tmp02_12_45;
	wire [WIDTH*2-1+2:0] tmp02_12_46;
	wire [WIDTH*2-1+2:0] tmp02_12_47;
	wire [WIDTH*2-1+2:0] tmp02_12_48;
	wire [WIDTH*2-1+2:0] tmp02_12_49;
	wire [WIDTH*2-1+2:0] tmp02_12_50;
	wire [WIDTH*2-1+2:0] tmp02_12_51;
	wire [WIDTH*2-1+2:0] tmp02_12_52;
	wire [WIDTH*2-1+2:0] tmp02_12_53;
	wire [WIDTH*2-1+2:0] tmp02_12_54;
	wire [WIDTH*2-1+2:0] tmp02_12_55;
	wire [WIDTH*2-1+2:0] tmp02_12_56;
	wire [WIDTH*2-1+2:0] tmp02_12_57;
	wire [WIDTH*2-1+2:0] tmp02_12_58;
	wire [WIDTH*2-1+2:0] tmp02_12_59;
	wire [WIDTH*2-1+2:0] tmp02_12_60;
	wire [WIDTH*2-1+2:0] tmp02_12_61;
	wire [WIDTH*2-1+2:0] tmp02_12_62;
	wire [WIDTH*2-1+2:0] tmp02_12_63;
	wire [WIDTH*2-1+2:0] tmp02_12_64;
	wire [WIDTH*2-1+2:0] tmp02_12_65;
	wire [WIDTH*2-1+2:0] tmp02_12_66;
	wire [WIDTH*2-1+2:0] tmp02_12_67;
	wire [WIDTH*2-1+2:0] tmp02_12_68;
	wire [WIDTH*2-1+2:0] tmp02_12_69;
	wire [WIDTH*2-1+2:0] tmp02_12_70;
	wire [WIDTH*2-1+2:0] tmp02_12_71;
	wire [WIDTH*2-1+2:0] tmp02_12_72;
	wire [WIDTH*2-1+2:0] tmp02_12_73;
	wire [WIDTH*2-1+2:0] tmp02_12_74;
	wire [WIDTH*2-1+2:0] tmp02_12_75;
	wire [WIDTH*2-1+2:0] tmp02_12_76;
	wire [WIDTH*2-1+2:0] tmp02_12_77;
	wire [WIDTH*2-1+2:0] tmp02_12_78;
	wire [WIDTH*2-1+2:0] tmp02_12_79;
	wire [WIDTH*2-1+2:0] tmp02_12_80;
	wire [WIDTH*2-1+2:0] tmp02_12_81;
	wire [WIDTH*2-1+2:0] tmp02_12_82;
	wire [WIDTH*2-1+2:0] tmp02_12_83;
	wire [WIDTH*2-1+2:0] tmp02_13_0;
	wire [WIDTH*2-1+2:0] tmp02_13_1;
	wire [WIDTH*2-1+2:0] tmp02_13_2;
	wire [WIDTH*2-1+2:0] tmp02_13_3;
	wire [WIDTH*2-1+2:0] tmp02_13_4;
	wire [WIDTH*2-1+2:0] tmp02_13_5;
	wire [WIDTH*2-1+2:0] tmp02_13_6;
	wire [WIDTH*2-1+2:0] tmp02_13_7;
	wire [WIDTH*2-1+2:0] tmp02_13_8;
	wire [WIDTH*2-1+2:0] tmp02_13_9;
	wire [WIDTH*2-1+2:0] tmp02_13_10;
	wire [WIDTH*2-1+2:0] tmp02_13_11;
	wire [WIDTH*2-1+2:0] tmp02_13_12;
	wire [WIDTH*2-1+2:0] tmp02_13_13;
	wire [WIDTH*2-1+2:0] tmp02_13_14;
	wire [WIDTH*2-1+2:0] tmp02_13_15;
	wire [WIDTH*2-1+2:0] tmp02_13_16;
	wire [WIDTH*2-1+2:0] tmp02_13_17;
	wire [WIDTH*2-1+2:0] tmp02_13_18;
	wire [WIDTH*2-1+2:0] tmp02_13_19;
	wire [WIDTH*2-1+2:0] tmp02_13_20;
	wire [WIDTH*2-1+2:0] tmp02_13_21;
	wire [WIDTH*2-1+2:0] tmp02_13_22;
	wire [WIDTH*2-1+2:0] tmp02_13_23;
	wire [WIDTH*2-1+2:0] tmp02_13_24;
	wire [WIDTH*2-1+2:0] tmp02_13_25;
	wire [WIDTH*2-1+2:0] tmp02_13_26;
	wire [WIDTH*2-1+2:0] tmp02_13_27;
	wire [WIDTH*2-1+2:0] tmp02_13_28;
	wire [WIDTH*2-1+2:0] tmp02_13_29;
	wire [WIDTH*2-1+2:0] tmp02_13_30;
	wire [WIDTH*2-1+2:0] tmp02_13_31;
	wire [WIDTH*2-1+2:0] tmp02_13_32;
	wire [WIDTH*2-1+2:0] tmp02_13_33;
	wire [WIDTH*2-1+2:0] tmp02_13_34;
	wire [WIDTH*2-1+2:0] tmp02_13_35;
	wire [WIDTH*2-1+2:0] tmp02_13_36;
	wire [WIDTH*2-1+2:0] tmp02_13_37;
	wire [WIDTH*2-1+2:0] tmp02_13_38;
	wire [WIDTH*2-1+2:0] tmp02_13_39;
	wire [WIDTH*2-1+2:0] tmp02_13_40;
	wire [WIDTH*2-1+2:0] tmp02_13_41;
	wire [WIDTH*2-1+2:0] tmp02_13_42;
	wire [WIDTH*2-1+2:0] tmp02_13_43;
	wire [WIDTH*2-1+2:0] tmp02_13_44;
	wire [WIDTH*2-1+2:0] tmp02_13_45;
	wire [WIDTH*2-1+2:0] tmp02_13_46;
	wire [WIDTH*2-1+2:0] tmp02_13_47;
	wire [WIDTH*2-1+2:0] tmp02_13_48;
	wire [WIDTH*2-1+2:0] tmp02_13_49;
	wire [WIDTH*2-1+2:0] tmp02_13_50;
	wire [WIDTH*2-1+2:0] tmp02_13_51;
	wire [WIDTH*2-1+2:0] tmp02_13_52;
	wire [WIDTH*2-1+2:0] tmp02_13_53;
	wire [WIDTH*2-1+2:0] tmp02_13_54;
	wire [WIDTH*2-1+2:0] tmp02_13_55;
	wire [WIDTH*2-1+2:0] tmp02_13_56;
	wire [WIDTH*2-1+2:0] tmp02_13_57;
	wire [WIDTH*2-1+2:0] tmp02_13_58;
	wire [WIDTH*2-1+2:0] tmp02_13_59;
	wire [WIDTH*2-1+2:0] tmp02_13_60;
	wire [WIDTH*2-1+2:0] tmp02_13_61;
	wire [WIDTH*2-1+2:0] tmp02_13_62;
	wire [WIDTH*2-1+2:0] tmp02_13_63;
	wire [WIDTH*2-1+2:0] tmp02_13_64;
	wire [WIDTH*2-1+2:0] tmp02_13_65;
	wire [WIDTH*2-1+2:0] tmp02_13_66;
	wire [WIDTH*2-1+2:0] tmp02_13_67;
	wire [WIDTH*2-1+2:0] tmp02_13_68;
	wire [WIDTH*2-1+2:0] tmp02_13_69;
	wire [WIDTH*2-1+2:0] tmp02_13_70;
	wire [WIDTH*2-1+2:0] tmp02_13_71;
	wire [WIDTH*2-1+2:0] tmp02_13_72;
	wire [WIDTH*2-1+2:0] tmp02_13_73;
	wire [WIDTH*2-1+2:0] tmp02_13_74;
	wire [WIDTH*2-1+2:0] tmp02_13_75;
	wire [WIDTH*2-1+2:0] tmp02_13_76;
	wire [WIDTH*2-1+2:0] tmp02_13_77;
	wire [WIDTH*2-1+2:0] tmp02_13_78;
	wire [WIDTH*2-1+2:0] tmp02_13_79;
	wire [WIDTH*2-1+2:0] tmp02_13_80;
	wire [WIDTH*2-1+2:0] tmp02_13_81;
	wire [WIDTH*2-1+2:0] tmp02_13_82;
	wire [WIDTH*2-1+2:0] tmp02_13_83;
	wire [WIDTH*2-1+2:0] tmp02_14_0;
	wire [WIDTH*2-1+2:0] tmp02_14_1;
	wire [WIDTH*2-1+2:0] tmp02_14_2;
	wire [WIDTH*2-1+2:0] tmp02_14_3;
	wire [WIDTH*2-1+2:0] tmp02_14_4;
	wire [WIDTH*2-1+2:0] tmp02_14_5;
	wire [WIDTH*2-1+2:0] tmp02_14_6;
	wire [WIDTH*2-1+2:0] tmp02_14_7;
	wire [WIDTH*2-1+2:0] tmp02_14_8;
	wire [WIDTH*2-1+2:0] tmp02_14_9;
	wire [WIDTH*2-1+2:0] tmp02_14_10;
	wire [WIDTH*2-1+2:0] tmp02_14_11;
	wire [WIDTH*2-1+2:0] tmp02_14_12;
	wire [WIDTH*2-1+2:0] tmp02_14_13;
	wire [WIDTH*2-1+2:0] tmp02_14_14;
	wire [WIDTH*2-1+2:0] tmp02_14_15;
	wire [WIDTH*2-1+2:0] tmp02_14_16;
	wire [WIDTH*2-1+2:0] tmp02_14_17;
	wire [WIDTH*2-1+2:0] tmp02_14_18;
	wire [WIDTH*2-1+2:0] tmp02_14_19;
	wire [WIDTH*2-1+2:0] tmp02_14_20;
	wire [WIDTH*2-1+2:0] tmp02_14_21;
	wire [WIDTH*2-1+2:0] tmp02_14_22;
	wire [WIDTH*2-1+2:0] tmp02_14_23;
	wire [WIDTH*2-1+2:0] tmp02_14_24;
	wire [WIDTH*2-1+2:0] tmp02_14_25;
	wire [WIDTH*2-1+2:0] tmp02_14_26;
	wire [WIDTH*2-1+2:0] tmp02_14_27;
	wire [WIDTH*2-1+2:0] tmp02_14_28;
	wire [WIDTH*2-1+2:0] tmp02_14_29;
	wire [WIDTH*2-1+2:0] tmp02_14_30;
	wire [WIDTH*2-1+2:0] tmp02_14_31;
	wire [WIDTH*2-1+2:0] tmp02_14_32;
	wire [WIDTH*2-1+2:0] tmp02_14_33;
	wire [WIDTH*2-1+2:0] tmp02_14_34;
	wire [WIDTH*2-1+2:0] tmp02_14_35;
	wire [WIDTH*2-1+2:0] tmp02_14_36;
	wire [WIDTH*2-1+2:0] tmp02_14_37;
	wire [WIDTH*2-1+2:0] tmp02_14_38;
	wire [WIDTH*2-1+2:0] tmp02_14_39;
	wire [WIDTH*2-1+2:0] tmp02_14_40;
	wire [WIDTH*2-1+2:0] tmp02_14_41;
	wire [WIDTH*2-1+2:0] tmp02_14_42;
	wire [WIDTH*2-1+2:0] tmp02_14_43;
	wire [WIDTH*2-1+2:0] tmp02_14_44;
	wire [WIDTH*2-1+2:0] tmp02_14_45;
	wire [WIDTH*2-1+2:0] tmp02_14_46;
	wire [WIDTH*2-1+2:0] tmp02_14_47;
	wire [WIDTH*2-1+2:0] tmp02_14_48;
	wire [WIDTH*2-1+2:0] tmp02_14_49;
	wire [WIDTH*2-1+2:0] tmp02_14_50;
	wire [WIDTH*2-1+2:0] tmp02_14_51;
	wire [WIDTH*2-1+2:0] tmp02_14_52;
	wire [WIDTH*2-1+2:0] tmp02_14_53;
	wire [WIDTH*2-1+2:0] tmp02_14_54;
	wire [WIDTH*2-1+2:0] tmp02_14_55;
	wire [WIDTH*2-1+2:0] tmp02_14_56;
	wire [WIDTH*2-1+2:0] tmp02_14_57;
	wire [WIDTH*2-1+2:0] tmp02_14_58;
	wire [WIDTH*2-1+2:0] tmp02_14_59;
	wire [WIDTH*2-1+2:0] tmp02_14_60;
	wire [WIDTH*2-1+2:0] tmp02_14_61;
	wire [WIDTH*2-1+2:0] tmp02_14_62;
	wire [WIDTH*2-1+2:0] tmp02_14_63;
	wire [WIDTH*2-1+2:0] tmp02_14_64;
	wire [WIDTH*2-1+2:0] tmp02_14_65;
	wire [WIDTH*2-1+2:0] tmp02_14_66;
	wire [WIDTH*2-1+2:0] tmp02_14_67;
	wire [WIDTH*2-1+2:0] tmp02_14_68;
	wire [WIDTH*2-1+2:0] tmp02_14_69;
	wire [WIDTH*2-1+2:0] tmp02_14_70;
	wire [WIDTH*2-1+2:0] tmp02_14_71;
	wire [WIDTH*2-1+2:0] tmp02_14_72;
	wire [WIDTH*2-1+2:0] tmp02_14_73;
	wire [WIDTH*2-1+2:0] tmp02_14_74;
	wire [WIDTH*2-1+2:0] tmp02_14_75;
	wire [WIDTH*2-1+2:0] tmp02_14_76;
	wire [WIDTH*2-1+2:0] tmp02_14_77;
	wire [WIDTH*2-1+2:0] tmp02_14_78;
	wire [WIDTH*2-1+2:0] tmp02_14_79;
	wire [WIDTH*2-1+2:0] tmp02_14_80;
	wire [WIDTH*2-1+2:0] tmp02_14_81;
	wire [WIDTH*2-1+2:0] tmp02_14_82;
	wire [WIDTH*2-1+2:0] tmp02_14_83;
	wire [WIDTH*2-1+2:0] tmp02_15_0;
	wire [WIDTH*2-1+2:0] tmp02_15_1;
	wire [WIDTH*2-1+2:0] tmp02_15_2;
	wire [WIDTH*2-1+2:0] tmp02_15_3;
	wire [WIDTH*2-1+2:0] tmp02_15_4;
	wire [WIDTH*2-1+2:0] tmp02_15_5;
	wire [WIDTH*2-1+2:0] tmp02_15_6;
	wire [WIDTH*2-1+2:0] tmp02_15_7;
	wire [WIDTH*2-1+2:0] tmp02_15_8;
	wire [WIDTH*2-1+2:0] tmp02_15_9;
	wire [WIDTH*2-1+2:0] tmp02_15_10;
	wire [WIDTH*2-1+2:0] tmp02_15_11;
	wire [WIDTH*2-1+2:0] tmp02_15_12;
	wire [WIDTH*2-1+2:0] tmp02_15_13;
	wire [WIDTH*2-1+2:0] tmp02_15_14;
	wire [WIDTH*2-1+2:0] tmp02_15_15;
	wire [WIDTH*2-1+2:0] tmp02_15_16;
	wire [WIDTH*2-1+2:0] tmp02_15_17;
	wire [WIDTH*2-1+2:0] tmp02_15_18;
	wire [WIDTH*2-1+2:0] tmp02_15_19;
	wire [WIDTH*2-1+2:0] tmp02_15_20;
	wire [WIDTH*2-1+2:0] tmp02_15_21;
	wire [WIDTH*2-1+2:0] tmp02_15_22;
	wire [WIDTH*2-1+2:0] tmp02_15_23;
	wire [WIDTH*2-1+2:0] tmp02_15_24;
	wire [WIDTH*2-1+2:0] tmp02_15_25;
	wire [WIDTH*2-1+2:0] tmp02_15_26;
	wire [WIDTH*2-1+2:0] tmp02_15_27;
	wire [WIDTH*2-1+2:0] tmp02_15_28;
	wire [WIDTH*2-1+2:0] tmp02_15_29;
	wire [WIDTH*2-1+2:0] tmp02_15_30;
	wire [WIDTH*2-1+2:0] tmp02_15_31;
	wire [WIDTH*2-1+2:0] tmp02_15_32;
	wire [WIDTH*2-1+2:0] tmp02_15_33;
	wire [WIDTH*2-1+2:0] tmp02_15_34;
	wire [WIDTH*2-1+2:0] tmp02_15_35;
	wire [WIDTH*2-1+2:0] tmp02_15_36;
	wire [WIDTH*2-1+2:0] tmp02_15_37;
	wire [WIDTH*2-1+2:0] tmp02_15_38;
	wire [WIDTH*2-1+2:0] tmp02_15_39;
	wire [WIDTH*2-1+2:0] tmp02_15_40;
	wire [WIDTH*2-1+2:0] tmp02_15_41;
	wire [WIDTH*2-1+2:0] tmp02_15_42;
	wire [WIDTH*2-1+2:0] tmp02_15_43;
	wire [WIDTH*2-1+2:0] tmp02_15_44;
	wire [WIDTH*2-1+2:0] tmp02_15_45;
	wire [WIDTH*2-1+2:0] tmp02_15_46;
	wire [WIDTH*2-1+2:0] tmp02_15_47;
	wire [WIDTH*2-1+2:0] tmp02_15_48;
	wire [WIDTH*2-1+2:0] tmp02_15_49;
	wire [WIDTH*2-1+2:0] tmp02_15_50;
	wire [WIDTH*2-1+2:0] tmp02_15_51;
	wire [WIDTH*2-1+2:0] tmp02_15_52;
	wire [WIDTH*2-1+2:0] tmp02_15_53;
	wire [WIDTH*2-1+2:0] tmp02_15_54;
	wire [WIDTH*2-1+2:0] tmp02_15_55;
	wire [WIDTH*2-1+2:0] tmp02_15_56;
	wire [WIDTH*2-1+2:0] tmp02_15_57;
	wire [WIDTH*2-1+2:0] tmp02_15_58;
	wire [WIDTH*2-1+2:0] tmp02_15_59;
	wire [WIDTH*2-1+2:0] tmp02_15_60;
	wire [WIDTH*2-1+2:0] tmp02_15_61;
	wire [WIDTH*2-1+2:0] tmp02_15_62;
	wire [WIDTH*2-1+2:0] tmp02_15_63;
	wire [WIDTH*2-1+2:0] tmp02_15_64;
	wire [WIDTH*2-1+2:0] tmp02_15_65;
	wire [WIDTH*2-1+2:0] tmp02_15_66;
	wire [WIDTH*2-1+2:0] tmp02_15_67;
	wire [WIDTH*2-1+2:0] tmp02_15_68;
	wire [WIDTH*2-1+2:0] tmp02_15_69;
	wire [WIDTH*2-1+2:0] tmp02_15_70;
	wire [WIDTH*2-1+2:0] tmp02_15_71;
	wire [WIDTH*2-1+2:0] tmp02_15_72;
	wire [WIDTH*2-1+2:0] tmp02_15_73;
	wire [WIDTH*2-1+2:0] tmp02_15_74;
	wire [WIDTH*2-1+2:0] tmp02_15_75;
	wire [WIDTH*2-1+2:0] tmp02_15_76;
	wire [WIDTH*2-1+2:0] tmp02_15_77;
	wire [WIDTH*2-1+2:0] tmp02_15_78;
	wire [WIDTH*2-1+2:0] tmp02_15_79;
	wire [WIDTH*2-1+2:0] tmp02_15_80;
	wire [WIDTH*2-1+2:0] tmp02_15_81;
	wire [WIDTH*2-1+2:0] tmp02_15_82;
	wire [WIDTH*2-1+2:0] tmp02_15_83;
	wire [WIDTH*2-1+2:0] tmp02_16_0;
	wire [WIDTH*2-1+2:0] tmp02_16_1;
	wire [WIDTH*2-1+2:0] tmp02_16_2;
	wire [WIDTH*2-1+2:0] tmp02_16_3;
	wire [WIDTH*2-1+2:0] tmp02_16_4;
	wire [WIDTH*2-1+2:0] tmp02_16_5;
	wire [WIDTH*2-1+2:0] tmp02_16_6;
	wire [WIDTH*2-1+2:0] tmp02_16_7;
	wire [WIDTH*2-1+2:0] tmp02_16_8;
	wire [WIDTH*2-1+2:0] tmp02_16_9;
	wire [WIDTH*2-1+2:0] tmp02_16_10;
	wire [WIDTH*2-1+2:0] tmp02_16_11;
	wire [WIDTH*2-1+2:0] tmp02_16_12;
	wire [WIDTH*2-1+2:0] tmp02_16_13;
	wire [WIDTH*2-1+2:0] tmp02_16_14;
	wire [WIDTH*2-1+2:0] tmp02_16_15;
	wire [WIDTH*2-1+2:0] tmp02_16_16;
	wire [WIDTH*2-1+2:0] tmp02_16_17;
	wire [WIDTH*2-1+2:0] tmp02_16_18;
	wire [WIDTH*2-1+2:0] tmp02_16_19;
	wire [WIDTH*2-1+2:0] tmp02_16_20;
	wire [WIDTH*2-1+2:0] tmp02_16_21;
	wire [WIDTH*2-1+2:0] tmp02_16_22;
	wire [WIDTH*2-1+2:0] tmp02_16_23;
	wire [WIDTH*2-1+2:0] tmp02_16_24;
	wire [WIDTH*2-1+2:0] tmp02_16_25;
	wire [WIDTH*2-1+2:0] tmp02_16_26;
	wire [WIDTH*2-1+2:0] tmp02_16_27;
	wire [WIDTH*2-1+2:0] tmp02_16_28;
	wire [WIDTH*2-1+2:0] tmp02_16_29;
	wire [WIDTH*2-1+2:0] tmp02_16_30;
	wire [WIDTH*2-1+2:0] tmp02_16_31;
	wire [WIDTH*2-1+2:0] tmp02_16_32;
	wire [WIDTH*2-1+2:0] tmp02_16_33;
	wire [WIDTH*2-1+2:0] tmp02_16_34;
	wire [WIDTH*2-1+2:0] tmp02_16_35;
	wire [WIDTH*2-1+2:0] tmp02_16_36;
	wire [WIDTH*2-1+2:0] tmp02_16_37;
	wire [WIDTH*2-1+2:0] tmp02_16_38;
	wire [WIDTH*2-1+2:0] tmp02_16_39;
	wire [WIDTH*2-1+2:0] tmp02_16_40;
	wire [WIDTH*2-1+2:0] tmp02_16_41;
	wire [WIDTH*2-1+2:0] tmp02_16_42;
	wire [WIDTH*2-1+2:0] tmp02_16_43;
	wire [WIDTH*2-1+2:0] tmp02_16_44;
	wire [WIDTH*2-1+2:0] tmp02_16_45;
	wire [WIDTH*2-1+2:0] tmp02_16_46;
	wire [WIDTH*2-1+2:0] tmp02_16_47;
	wire [WIDTH*2-1+2:0] tmp02_16_48;
	wire [WIDTH*2-1+2:0] tmp02_16_49;
	wire [WIDTH*2-1+2:0] tmp02_16_50;
	wire [WIDTH*2-1+2:0] tmp02_16_51;
	wire [WIDTH*2-1+2:0] tmp02_16_52;
	wire [WIDTH*2-1+2:0] tmp02_16_53;
	wire [WIDTH*2-1+2:0] tmp02_16_54;
	wire [WIDTH*2-1+2:0] tmp02_16_55;
	wire [WIDTH*2-1+2:0] tmp02_16_56;
	wire [WIDTH*2-1+2:0] tmp02_16_57;
	wire [WIDTH*2-1+2:0] tmp02_16_58;
	wire [WIDTH*2-1+2:0] tmp02_16_59;
	wire [WIDTH*2-1+2:0] tmp02_16_60;
	wire [WIDTH*2-1+2:0] tmp02_16_61;
	wire [WIDTH*2-1+2:0] tmp02_16_62;
	wire [WIDTH*2-1+2:0] tmp02_16_63;
	wire [WIDTH*2-1+2:0] tmp02_16_64;
	wire [WIDTH*2-1+2:0] tmp02_16_65;
	wire [WIDTH*2-1+2:0] tmp02_16_66;
	wire [WIDTH*2-1+2:0] tmp02_16_67;
	wire [WIDTH*2-1+2:0] tmp02_16_68;
	wire [WIDTH*2-1+2:0] tmp02_16_69;
	wire [WIDTH*2-1+2:0] tmp02_16_70;
	wire [WIDTH*2-1+2:0] tmp02_16_71;
	wire [WIDTH*2-1+2:0] tmp02_16_72;
	wire [WIDTH*2-1+2:0] tmp02_16_73;
	wire [WIDTH*2-1+2:0] tmp02_16_74;
	wire [WIDTH*2-1+2:0] tmp02_16_75;
	wire [WIDTH*2-1+2:0] tmp02_16_76;
	wire [WIDTH*2-1+2:0] tmp02_16_77;
	wire [WIDTH*2-1+2:0] tmp02_16_78;
	wire [WIDTH*2-1+2:0] tmp02_16_79;
	wire [WIDTH*2-1+2:0] tmp02_16_80;
	wire [WIDTH*2-1+2:0] tmp02_16_81;
	wire [WIDTH*2-1+2:0] tmp02_16_82;
	wire [WIDTH*2-1+2:0] tmp02_16_83;
	wire [WIDTH*2-1+2:0] tmp02_17_0;
	wire [WIDTH*2-1+2:0] tmp02_17_1;
	wire [WIDTH*2-1+2:0] tmp02_17_2;
	wire [WIDTH*2-1+2:0] tmp02_17_3;
	wire [WIDTH*2-1+2:0] tmp02_17_4;
	wire [WIDTH*2-1+2:0] tmp02_17_5;
	wire [WIDTH*2-1+2:0] tmp02_17_6;
	wire [WIDTH*2-1+2:0] tmp02_17_7;
	wire [WIDTH*2-1+2:0] tmp02_17_8;
	wire [WIDTH*2-1+2:0] tmp02_17_9;
	wire [WIDTH*2-1+2:0] tmp02_17_10;
	wire [WIDTH*2-1+2:0] tmp02_17_11;
	wire [WIDTH*2-1+2:0] tmp02_17_12;
	wire [WIDTH*2-1+2:0] tmp02_17_13;
	wire [WIDTH*2-1+2:0] tmp02_17_14;
	wire [WIDTH*2-1+2:0] tmp02_17_15;
	wire [WIDTH*2-1+2:0] tmp02_17_16;
	wire [WIDTH*2-1+2:0] tmp02_17_17;
	wire [WIDTH*2-1+2:0] tmp02_17_18;
	wire [WIDTH*2-1+2:0] tmp02_17_19;
	wire [WIDTH*2-1+2:0] tmp02_17_20;
	wire [WIDTH*2-1+2:0] tmp02_17_21;
	wire [WIDTH*2-1+2:0] tmp02_17_22;
	wire [WIDTH*2-1+2:0] tmp02_17_23;
	wire [WIDTH*2-1+2:0] tmp02_17_24;
	wire [WIDTH*2-1+2:0] tmp02_17_25;
	wire [WIDTH*2-1+2:0] tmp02_17_26;
	wire [WIDTH*2-1+2:0] tmp02_17_27;
	wire [WIDTH*2-1+2:0] tmp02_17_28;
	wire [WIDTH*2-1+2:0] tmp02_17_29;
	wire [WIDTH*2-1+2:0] tmp02_17_30;
	wire [WIDTH*2-1+2:0] tmp02_17_31;
	wire [WIDTH*2-1+2:0] tmp02_17_32;
	wire [WIDTH*2-1+2:0] tmp02_17_33;
	wire [WIDTH*2-1+2:0] tmp02_17_34;
	wire [WIDTH*2-1+2:0] tmp02_17_35;
	wire [WIDTH*2-1+2:0] tmp02_17_36;
	wire [WIDTH*2-1+2:0] tmp02_17_37;
	wire [WIDTH*2-1+2:0] tmp02_17_38;
	wire [WIDTH*2-1+2:0] tmp02_17_39;
	wire [WIDTH*2-1+2:0] tmp02_17_40;
	wire [WIDTH*2-1+2:0] tmp02_17_41;
	wire [WIDTH*2-1+2:0] tmp02_17_42;
	wire [WIDTH*2-1+2:0] tmp02_17_43;
	wire [WIDTH*2-1+2:0] tmp02_17_44;
	wire [WIDTH*2-1+2:0] tmp02_17_45;
	wire [WIDTH*2-1+2:0] tmp02_17_46;
	wire [WIDTH*2-1+2:0] tmp02_17_47;
	wire [WIDTH*2-1+2:0] tmp02_17_48;
	wire [WIDTH*2-1+2:0] tmp02_17_49;
	wire [WIDTH*2-1+2:0] tmp02_17_50;
	wire [WIDTH*2-1+2:0] tmp02_17_51;
	wire [WIDTH*2-1+2:0] tmp02_17_52;
	wire [WIDTH*2-1+2:0] tmp02_17_53;
	wire [WIDTH*2-1+2:0] tmp02_17_54;
	wire [WIDTH*2-1+2:0] tmp02_17_55;
	wire [WIDTH*2-1+2:0] tmp02_17_56;
	wire [WIDTH*2-1+2:0] tmp02_17_57;
	wire [WIDTH*2-1+2:0] tmp02_17_58;
	wire [WIDTH*2-1+2:0] tmp02_17_59;
	wire [WIDTH*2-1+2:0] tmp02_17_60;
	wire [WIDTH*2-1+2:0] tmp02_17_61;
	wire [WIDTH*2-1+2:0] tmp02_17_62;
	wire [WIDTH*2-1+2:0] tmp02_17_63;
	wire [WIDTH*2-1+2:0] tmp02_17_64;
	wire [WIDTH*2-1+2:0] tmp02_17_65;
	wire [WIDTH*2-1+2:0] tmp02_17_66;
	wire [WIDTH*2-1+2:0] tmp02_17_67;
	wire [WIDTH*2-1+2:0] tmp02_17_68;
	wire [WIDTH*2-1+2:0] tmp02_17_69;
	wire [WIDTH*2-1+2:0] tmp02_17_70;
	wire [WIDTH*2-1+2:0] tmp02_17_71;
	wire [WIDTH*2-1+2:0] tmp02_17_72;
	wire [WIDTH*2-1+2:0] tmp02_17_73;
	wire [WIDTH*2-1+2:0] tmp02_17_74;
	wire [WIDTH*2-1+2:0] tmp02_17_75;
	wire [WIDTH*2-1+2:0] tmp02_17_76;
	wire [WIDTH*2-1+2:0] tmp02_17_77;
	wire [WIDTH*2-1+2:0] tmp02_17_78;
	wire [WIDTH*2-1+2:0] tmp02_17_79;
	wire [WIDTH*2-1+2:0] tmp02_17_80;
	wire [WIDTH*2-1+2:0] tmp02_17_81;
	wire [WIDTH*2-1+2:0] tmp02_17_82;
	wire [WIDTH*2-1+2:0] tmp02_17_83;
	wire [WIDTH*2-1+2:0] tmp02_18_0;
	wire [WIDTH*2-1+2:0] tmp02_18_1;
	wire [WIDTH*2-1+2:0] tmp02_18_2;
	wire [WIDTH*2-1+2:0] tmp02_18_3;
	wire [WIDTH*2-1+2:0] tmp02_18_4;
	wire [WIDTH*2-1+2:0] tmp02_18_5;
	wire [WIDTH*2-1+2:0] tmp02_18_6;
	wire [WIDTH*2-1+2:0] tmp02_18_7;
	wire [WIDTH*2-1+2:0] tmp02_18_8;
	wire [WIDTH*2-1+2:0] tmp02_18_9;
	wire [WIDTH*2-1+2:0] tmp02_18_10;
	wire [WIDTH*2-1+2:0] tmp02_18_11;
	wire [WIDTH*2-1+2:0] tmp02_18_12;
	wire [WIDTH*2-1+2:0] tmp02_18_13;
	wire [WIDTH*2-1+2:0] tmp02_18_14;
	wire [WIDTH*2-1+2:0] tmp02_18_15;
	wire [WIDTH*2-1+2:0] tmp02_18_16;
	wire [WIDTH*2-1+2:0] tmp02_18_17;
	wire [WIDTH*2-1+2:0] tmp02_18_18;
	wire [WIDTH*2-1+2:0] tmp02_18_19;
	wire [WIDTH*2-1+2:0] tmp02_18_20;
	wire [WIDTH*2-1+2:0] tmp02_18_21;
	wire [WIDTH*2-1+2:0] tmp02_18_22;
	wire [WIDTH*2-1+2:0] tmp02_18_23;
	wire [WIDTH*2-1+2:0] tmp02_18_24;
	wire [WIDTH*2-1+2:0] tmp02_18_25;
	wire [WIDTH*2-1+2:0] tmp02_18_26;
	wire [WIDTH*2-1+2:0] tmp02_18_27;
	wire [WIDTH*2-1+2:0] tmp02_18_28;
	wire [WIDTH*2-1+2:0] tmp02_18_29;
	wire [WIDTH*2-1+2:0] tmp02_18_30;
	wire [WIDTH*2-1+2:0] tmp02_18_31;
	wire [WIDTH*2-1+2:0] tmp02_18_32;
	wire [WIDTH*2-1+2:0] tmp02_18_33;
	wire [WIDTH*2-1+2:0] tmp02_18_34;
	wire [WIDTH*2-1+2:0] tmp02_18_35;
	wire [WIDTH*2-1+2:0] tmp02_18_36;
	wire [WIDTH*2-1+2:0] tmp02_18_37;
	wire [WIDTH*2-1+2:0] tmp02_18_38;
	wire [WIDTH*2-1+2:0] tmp02_18_39;
	wire [WIDTH*2-1+2:0] tmp02_18_40;
	wire [WIDTH*2-1+2:0] tmp02_18_41;
	wire [WIDTH*2-1+2:0] tmp02_18_42;
	wire [WIDTH*2-1+2:0] tmp02_18_43;
	wire [WIDTH*2-1+2:0] tmp02_18_44;
	wire [WIDTH*2-1+2:0] tmp02_18_45;
	wire [WIDTH*2-1+2:0] tmp02_18_46;
	wire [WIDTH*2-1+2:0] tmp02_18_47;
	wire [WIDTH*2-1+2:0] tmp02_18_48;
	wire [WIDTH*2-1+2:0] tmp02_18_49;
	wire [WIDTH*2-1+2:0] tmp02_18_50;
	wire [WIDTH*2-1+2:0] tmp02_18_51;
	wire [WIDTH*2-1+2:0] tmp02_18_52;
	wire [WIDTH*2-1+2:0] tmp02_18_53;
	wire [WIDTH*2-1+2:0] tmp02_18_54;
	wire [WIDTH*2-1+2:0] tmp02_18_55;
	wire [WIDTH*2-1+2:0] tmp02_18_56;
	wire [WIDTH*2-1+2:0] tmp02_18_57;
	wire [WIDTH*2-1+2:0] tmp02_18_58;
	wire [WIDTH*2-1+2:0] tmp02_18_59;
	wire [WIDTH*2-1+2:0] tmp02_18_60;
	wire [WIDTH*2-1+2:0] tmp02_18_61;
	wire [WIDTH*2-1+2:0] tmp02_18_62;
	wire [WIDTH*2-1+2:0] tmp02_18_63;
	wire [WIDTH*2-1+2:0] tmp02_18_64;
	wire [WIDTH*2-1+2:0] tmp02_18_65;
	wire [WIDTH*2-1+2:0] tmp02_18_66;
	wire [WIDTH*2-1+2:0] tmp02_18_67;
	wire [WIDTH*2-1+2:0] tmp02_18_68;
	wire [WIDTH*2-1+2:0] tmp02_18_69;
	wire [WIDTH*2-1+2:0] tmp02_18_70;
	wire [WIDTH*2-1+2:0] tmp02_18_71;
	wire [WIDTH*2-1+2:0] tmp02_18_72;
	wire [WIDTH*2-1+2:0] tmp02_18_73;
	wire [WIDTH*2-1+2:0] tmp02_18_74;
	wire [WIDTH*2-1+2:0] tmp02_18_75;
	wire [WIDTH*2-1+2:0] tmp02_18_76;
	wire [WIDTH*2-1+2:0] tmp02_18_77;
	wire [WIDTH*2-1+2:0] tmp02_18_78;
	wire [WIDTH*2-1+2:0] tmp02_18_79;
	wire [WIDTH*2-1+2:0] tmp02_18_80;
	wire [WIDTH*2-1+2:0] tmp02_18_81;
	wire [WIDTH*2-1+2:0] tmp02_18_82;
	wire [WIDTH*2-1+2:0] tmp02_18_83;
	wire [WIDTH*2-1+2:0] tmp02_19_0;
	wire [WIDTH*2-1+2:0] tmp02_19_1;
	wire [WIDTH*2-1+2:0] tmp02_19_2;
	wire [WIDTH*2-1+2:0] tmp02_19_3;
	wire [WIDTH*2-1+2:0] tmp02_19_4;
	wire [WIDTH*2-1+2:0] tmp02_19_5;
	wire [WIDTH*2-1+2:0] tmp02_19_6;
	wire [WIDTH*2-1+2:0] tmp02_19_7;
	wire [WIDTH*2-1+2:0] tmp02_19_8;
	wire [WIDTH*2-1+2:0] tmp02_19_9;
	wire [WIDTH*2-1+2:0] tmp02_19_10;
	wire [WIDTH*2-1+2:0] tmp02_19_11;
	wire [WIDTH*2-1+2:0] tmp02_19_12;
	wire [WIDTH*2-1+2:0] tmp02_19_13;
	wire [WIDTH*2-1+2:0] tmp02_19_14;
	wire [WIDTH*2-1+2:0] tmp02_19_15;
	wire [WIDTH*2-1+2:0] tmp02_19_16;
	wire [WIDTH*2-1+2:0] tmp02_19_17;
	wire [WIDTH*2-1+2:0] tmp02_19_18;
	wire [WIDTH*2-1+2:0] tmp02_19_19;
	wire [WIDTH*2-1+2:0] tmp02_19_20;
	wire [WIDTH*2-1+2:0] tmp02_19_21;
	wire [WIDTH*2-1+2:0] tmp02_19_22;
	wire [WIDTH*2-1+2:0] tmp02_19_23;
	wire [WIDTH*2-1+2:0] tmp02_19_24;
	wire [WIDTH*2-1+2:0] tmp02_19_25;
	wire [WIDTH*2-1+2:0] tmp02_19_26;
	wire [WIDTH*2-1+2:0] tmp02_19_27;
	wire [WIDTH*2-1+2:0] tmp02_19_28;
	wire [WIDTH*2-1+2:0] tmp02_19_29;
	wire [WIDTH*2-1+2:0] tmp02_19_30;
	wire [WIDTH*2-1+2:0] tmp02_19_31;
	wire [WIDTH*2-1+2:0] tmp02_19_32;
	wire [WIDTH*2-1+2:0] tmp02_19_33;
	wire [WIDTH*2-1+2:0] tmp02_19_34;
	wire [WIDTH*2-1+2:0] tmp02_19_35;
	wire [WIDTH*2-1+2:0] tmp02_19_36;
	wire [WIDTH*2-1+2:0] tmp02_19_37;
	wire [WIDTH*2-1+2:0] tmp02_19_38;
	wire [WIDTH*2-1+2:0] tmp02_19_39;
	wire [WIDTH*2-1+2:0] tmp02_19_40;
	wire [WIDTH*2-1+2:0] tmp02_19_41;
	wire [WIDTH*2-1+2:0] tmp02_19_42;
	wire [WIDTH*2-1+2:0] tmp02_19_43;
	wire [WIDTH*2-1+2:0] tmp02_19_44;
	wire [WIDTH*2-1+2:0] tmp02_19_45;
	wire [WIDTH*2-1+2:0] tmp02_19_46;
	wire [WIDTH*2-1+2:0] tmp02_19_47;
	wire [WIDTH*2-1+2:0] tmp02_19_48;
	wire [WIDTH*2-1+2:0] tmp02_19_49;
	wire [WIDTH*2-1+2:0] tmp02_19_50;
	wire [WIDTH*2-1+2:0] tmp02_19_51;
	wire [WIDTH*2-1+2:0] tmp02_19_52;
	wire [WIDTH*2-1+2:0] tmp02_19_53;
	wire [WIDTH*2-1+2:0] tmp02_19_54;
	wire [WIDTH*2-1+2:0] tmp02_19_55;
	wire [WIDTH*2-1+2:0] tmp02_19_56;
	wire [WIDTH*2-1+2:0] tmp02_19_57;
	wire [WIDTH*2-1+2:0] tmp02_19_58;
	wire [WIDTH*2-1+2:0] tmp02_19_59;
	wire [WIDTH*2-1+2:0] tmp02_19_60;
	wire [WIDTH*2-1+2:0] tmp02_19_61;
	wire [WIDTH*2-1+2:0] tmp02_19_62;
	wire [WIDTH*2-1+2:0] tmp02_19_63;
	wire [WIDTH*2-1+2:0] tmp02_19_64;
	wire [WIDTH*2-1+2:0] tmp02_19_65;
	wire [WIDTH*2-1+2:0] tmp02_19_66;
	wire [WIDTH*2-1+2:0] tmp02_19_67;
	wire [WIDTH*2-1+2:0] tmp02_19_68;
	wire [WIDTH*2-1+2:0] tmp02_19_69;
	wire [WIDTH*2-1+2:0] tmp02_19_70;
	wire [WIDTH*2-1+2:0] tmp02_19_71;
	wire [WIDTH*2-1+2:0] tmp02_19_72;
	wire [WIDTH*2-1+2:0] tmp02_19_73;
	wire [WIDTH*2-1+2:0] tmp02_19_74;
	wire [WIDTH*2-1+2:0] tmp02_19_75;
	wire [WIDTH*2-1+2:0] tmp02_19_76;
	wire [WIDTH*2-1+2:0] tmp02_19_77;
	wire [WIDTH*2-1+2:0] tmp02_19_78;
	wire [WIDTH*2-1+2:0] tmp02_19_79;
	wire [WIDTH*2-1+2:0] tmp02_19_80;
	wire [WIDTH*2-1+2:0] tmp02_19_81;
	wire [WIDTH*2-1+2:0] tmp02_19_82;
	wire [WIDTH*2-1+2:0] tmp02_19_83;
	wire [WIDTH*2-1+2:0] tmp02_20_0;
	wire [WIDTH*2-1+2:0] tmp02_20_1;
	wire [WIDTH*2-1+2:0] tmp02_20_2;
	wire [WIDTH*2-1+2:0] tmp02_20_3;
	wire [WIDTH*2-1+2:0] tmp02_20_4;
	wire [WIDTH*2-1+2:0] tmp02_20_5;
	wire [WIDTH*2-1+2:0] tmp02_20_6;
	wire [WIDTH*2-1+2:0] tmp02_20_7;
	wire [WIDTH*2-1+2:0] tmp02_20_8;
	wire [WIDTH*2-1+2:0] tmp02_20_9;
	wire [WIDTH*2-1+2:0] tmp02_20_10;
	wire [WIDTH*2-1+2:0] tmp02_20_11;
	wire [WIDTH*2-1+2:0] tmp02_20_12;
	wire [WIDTH*2-1+2:0] tmp02_20_13;
	wire [WIDTH*2-1+2:0] tmp02_20_14;
	wire [WIDTH*2-1+2:0] tmp02_20_15;
	wire [WIDTH*2-1+2:0] tmp02_20_16;
	wire [WIDTH*2-1+2:0] tmp02_20_17;
	wire [WIDTH*2-1+2:0] tmp02_20_18;
	wire [WIDTH*2-1+2:0] tmp02_20_19;
	wire [WIDTH*2-1+2:0] tmp02_20_20;
	wire [WIDTH*2-1+2:0] tmp02_20_21;
	wire [WIDTH*2-1+2:0] tmp02_20_22;
	wire [WIDTH*2-1+2:0] tmp02_20_23;
	wire [WIDTH*2-1+2:0] tmp02_20_24;
	wire [WIDTH*2-1+2:0] tmp02_20_25;
	wire [WIDTH*2-1+2:0] tmp02_20_26;
	wire [WIDTH*2-1+2:0] tmp02_20_27;
	wire [WIDTH*2-1+2:0] tmp02_20_28;
	wire [WIDTH*2-1+2:0] tmp02_20_29;
	wire [WIDTH*2-1+2:0] tmp02_20_30;
	wire [WIDTH*2-1+2:0] tmp02_20_31;
	wire [WIDTH*2-1+2:0] tmp02_20_32;
	wire [WIDTH*2-1+2:0] tmp02_20_33;
	wire [WIDTH*2-1+2:0] tmp02_20_34;
	wire [WIDTH*2-1+2:0] tmp02_20_35;
	wire [WIDTH*2-1+2:0] tmp02_20_36;
	wire [WIDTH*2-1+2:0] tmp02_20_37;
	wire [WIDTH*2-1+2:0] tmp02_20_38;
	wire [WIDTH*2-1+2:0] tmp02_20_39;
	wire [WIDTH*2-1+2:0] tmp02_20_40;
	wire [WIDTH*2-1+2:0] tmp02_20_41;
	wire [WIDTH*2-1+2:0] tmp02_20_42;
	wire [WIDTH*2-1+2:0] tmp02_20_43;
	wire [WIDTH*2-1+2:0] tmp02_20_44;
	wire [WIDTH*2-1+2:0] tmp02_20_45;
	wire [WIDTH*2-1+2:0] tmp02_20_46;
	wire [WIDTH*2-1+2:0] tmp02_20_47;
	wire [WIDTH*2-1+2:0] tmp02_20_48;
	wire [WIDTH*2-1+2:0] tmp02_20_49;
	wire [WIDTH*2-1+2:0] tmp02_20_50;
	wire [WIDTH*2-1+2:0] tmp02_20_51;
	wire [WIDTH*2-1+2:0] tmp02_20_52;
	wire [WIDTH*2-1+2:0] tmp02_20_53;
	wire [WIDTH*2-1+2:0] tmp02_20_54;
	wire [WIDTH*2-1+2:0] tmp02_20_55;
	wire [WIDTH*2-1+2:0] tmp02_20_56;
	wire [WIDTH*2-1+2:0] tmp02_20_57;
	wire [WIDTH*2-1+2:0] tmp02_20_58;
	wire [WIDTH*2-1+2:0] tmp02_20_59;
	wire [WIDTH*2-1+2:0] tmp02_20_60;
	wire [WIDTH*2-1+2:0] tmp02_20_61;
	wire [WIDTH*2-1+2:0] tmp02_20_62;
	wire [WIDTH*2-1+2:0] tmp02_20_63;
	wire [WIDTH*2-1+2:0] tmp02_20_64;
	wire [WIDTH*2-1+2:0] tmp02_20_65;
	wire [WIDTH*2-1+2:0] tmp02_20_66;
	wire [WIDTH*2-1+2:0] tmp02_20_67;
	wire [WIDTH*2-1+2:0] tmp02_20_68;
	wire [WIDTH*2-1+2:0] tmp02_20_69;
	wire [WIDTH*2-1+2:0] tmp02_20_70;
	wire [WIDTH*2-1+2:0] tmp02_20_71;
	wire [WIDTH*2-1+2:0] tmp02_20_72;
	wire [WIDTH*2-1+2:0] tmp02_20_73;
	wire [WIDTH*2-1+2:0] tmp02_20_74;
	wire [WIDTH*2-1+2:0] tmp02_20_75;
	wire [WIDTH*2-1+2:0] tmp02_20_76;
	wire [WIDTH*2-1+2:0] tmp02_20_77;
	wire [WIDTH*2-1+2:0] tmp02_20_78;
	wire [WIDTH*2-1+2:0] tmp02_20_79;
	wire [WIDTH*2-1+2:0] tmp02_20_80;
	wire [WIDTH*2-1+2:0] tmp02_20_81;
	wire [WIDTH*2-1+2:0] tmp02_20_82;
	wire [WIDTH*2-1+2:0] tmp02_20_83;
	wire [WIDTH*2-1+2:0] tmp02_21_0;
	wire [WIDTH*2-1+2:0] tmp02_21_1;
	wire [WIDTH*2-1+2:0] tmp02_21_2;
	wire [WIDTH*2-1+2:0] tmp02_21_3;
	wire [WIDTH*2-1+2:0] tmp02_21_4;
	wire [WIDTH*2-1+2:0] tmp02_21_5;
	wire [WIDTH*2-1+2:0] tmp02_21_6;
	wire [WIDTH*2-1+2:0] tmp02_21_7;
	wire [WIDTH*2-1+2:0] tmp02_21_8;
	wire [WIDTH*2-1+2:0] tmp02_21_9;
	wire [WIDTH*2-1+2:0] tmp02_21_10;
	wire [WIDTH*2-1+2:0] tmp02_21_11;
	wire [WIDTH*2-1+2:0] tmp02_21_12;
	wire [WIDTH*2-1+2:0] tmp02_21_13;
	wire [WIDTH*2-1+2:0] tmp02_21_14;
	wire [WIDTH*2-1+2:0] tmp02_21_15;
	wire [WIDTH*2-1+2:0] tmp02_21_16;
	wire [WIDTH*2-1+2:0] tmp02_21_17;
	wire [WIDTH*2-1+2:0] tmp02_21_18;
	wire [WIDTH*2-1+2:0] tmp02_21_19;
	wire [WIDTH*2-1+2:0] tmp02_21_20;
	wire [WIDTH*2-1+2:0] tmp02_21_21;
	wire [WIDTH*2-1+2:0] tmp02_21_22;
	wire [WIDTH*2-1+2:0] tmp02_21_23;
	wire [WIDTH*2-1+2:0] tmp02_21_24;
	wire [WIDTH*2-1+2:0] tmp02_21_25;
	wire [WIDTH*2-1+2:0] tmp02_21_26;
	wire [WIDTH*2-1+2:0] tmp02_21_27;
	wire [WIDTH*2-1+2:0] tmp02_21_28;
	wire [WIDTH*2-1+2:0] tmp02_21_29;
	wire [WIDTH*2-1+2:0] tmp02_21_30;
	wire [WIDTH*2-1+2:0] tmp02_21_31;
	wire [WIDTH*2-1+2:0] tmp02_21_32;
	wire [WIDTH*2-1+2:0] tmp02_21_33;
	wire [WIDTH*2-1+2:0] tmp02_21_34;
	wire [WIDTH*2-1+2:0] tmp02_21_35;
	wire [WIDTH*2-1+2:0] tmp02_21_36;
	wire [WIDTH*2-1+2:0] tmp02_21_37;
	wire [WIDTH*2-1+2:0] tmp02_21_38;
	wire [WIDTH*2-1+2:0] tmp02_21_39;
	wire [WIDTH*2-1+2:0] tmp02_21_40;
	wire [WIDTH*2-1+2:0] tmp02_21_41;
	wire [WIDTH*2-1+2:0] tmp02_21_42;
	wire [WIDTH*2-1+2:0] tmp02_21_43;
	wire [WIDTH*2-1+2:0] tmp02_21_44;
	wire [WIDTH*2-1+2:0] tmp02_21_45;
	wire [WIDTH*2-1+2:0] tmp02_21_46;
	wire [WIDTH*2-1+2:0] tmp02_21_47;
	wire [WIDTH*2-1+2:0] tmp02_21_48;
	wire [WIDTH*2-1+2:0] tmp02_21_49;
	wire [WIDTH*2-1+2:0] tmp02_21_50;
	wire [WIDTH*2-1+2:0] tmp02_21_51;
	wire [WIDTH*2-1+2:0] tmp02_21_52;
	wire [WIDTH*2-1+2:0] tmp02_21_53;
	wire [WIDTH*2-1+2:0] tmp02_21_54;
	wire [WIDTH*2-1+2:0] tmp02_21_55;
	wire [WIDTH*2-1+2:0] tmp02_21_56;
	wire [WIDTH*2-1+2:0] tmp02_21_57;
	wire [WIDTH*2-1+2:0] tmp02_21_58;
	wire [WIDTH*2-1+2:0] tmp02_21_59;
	wire [WIDTH*2-1+2:0] tmp02_21_60;
	wire [WIDTH*2-1+2:0] tmp02_21_61;
	wire [WIDTH*2-1+2:0] tmp02_21_62;
	wire [WIDTH*2-1+2:0] tmp02_21_63;
	wire [WIDTH*2-1+2:0] tmp02_21_64;
	wire [WIDTH*2-1+2:0] tmp02_21_65;
	wire [WIDTH*2-1+2:0] tmp02_21_66;
	wire [WIDTH*2-1+2:0] tmp02_21_67;
	wire [WIDTH*2-1+2:0] tmp02_21_68;
	wire [WIDTH*2-1+2:0] tmp02_21_69;
	wire [WIDTH*2-1+2:0] tmp02_21_70;
	wire [WIDTH*2-1+2:0] tmp02_21_71;
	wire [WIDTH*2-1+2:0] tmp02_21_72;
	wire [WIDTH*2-1+2:0] tmp02_21_73;
	wire [WIDTH*2-1+2:0] tmp02_21_74;
	wire [WIDTH*2-1+2:0] tmp02_21_75;
	wire [WIDTH*2-1+2:0] tmp02_21_76;
	wire [WIDTH*2-1+2:0] tmp02_21_77;
	wire [WIDTH*2-1+2:0] tmp02_21_78;
	wire [WIDTH*2-1+2:0] tmp02_21_79;
	wire [WIDTH*2-1+2:0] tmp02_21_80;
	wire [WIDTH*2-1+2:0] tmp02_21_81;
	wire [WIDTH*2-1+2:0] tmp02_21_82;
	wire [WIDTH*2-1+2:0] tmp02_21_83;
	wire [WIDTH*2-1+2:0] tmp02_22_0;
	wire [WIDTH*2-1+2:0] tmp02_22_1;
	wire [WIDTH*2-1+2:0] tmp02_22_2;
	wire [WIDTH*2-1+2:0] tmp02_22_3;
	wire [WIDTH*2-1+2:0] tmp02_22_4;
	wire [WIDTH*2-1+2:0] tmp02_22_5;
	wire [WIDTH*2-1+2:0] tmp02_22_6;
	wire [WIDTH*2-1+2:0] tmp02_22_7;
	wire [WIDTH*2-1+2:0] tmp02_22_8;
	wire [WIDTH*2-1+2:0] tmp02_22_9;
	wire [WIDTH*2-1+2:0] tmp02_22_10;
	wire [WIDTH*2-1+2:0] tmp02_22_11;
	wire [WIDTH*2-1+2:0] tmp02_22_12;
	wire [WIDTH*2-1+2:0] tmp02_22_13;
	wire [WIDTH*2-1+2:0] tmp02_22_14;
	wire [WIDTH*2-1+2:0] tmp02_22_15;
	wire [WIDTH*2-1+2:0] tmp02_22_16;
	wire [WIDTH*2-1+2:0] tmp02_22_17;
	wire [WIDTH*2-1+2:0] tmp02_22_18;
	wire [WIDTH*2-1+2:0] tmp02_22_19;
	wire [WIDTH*2-1+2:0] tmp02_22_20;
	wire [WIDTH*2-1+2:0] tmp02_22_21;
	wire [WIDTH*2-1+2:0] tmp02_22_22;
	wire [WIDTH*2-1+2:0] tmp02_22_23;
	wire [WIDTH*2-1+2:0] tmp02_22_24;
	wire [WIDTH*2-1+2:0] tmp02_22_25;
	wire [WIDTH*2-1+2:0] tmp02_22_26;
	wire [WIDTH*2-1+2:0] tmp02_22_27;
	wire [WIDTH*2-1+2:0] tmp02_22_28;
	wire [WIDTH*2-1+2:0] tmp02_22_29;
	wire [WIDTH*2-1+2:0] tmp02_22_30;
	wire [WIDTH*2-1+2:0] tmp02_22_31;
	wire [WIDTH*2-1+2:0] tmp02_22_32;
	wire [WIDTH*2-1+2:0] tmp02_22_33;
	wire [WIDTH*2-1+2:0] tmp02_22_34;
	wire [WIDTH*2-1+2:0] tmp02_22_35;
	wire [WIDTH*2-1+2:0] tmp02_22_36;
	wire [WIDTH*2-1+2:0] tmp02_22_37;
	wire [WIDTH*2-1+2:0] tmp02_22_38;
	wire [WIDTH*2-1+2:0] tmp02_22_39;
	wire [WIDTH*2-1+2:0] tmp02_22_40;
	wire [WIDTH*2-1+2:0] tmp02_22_41;
	wire [WIDTH*2-1+2:0] tmp02_22_42;
	wire [WIDTH*2-1+2:0] tmp02_22_43;
	wire [WIDTH*2-1+2:0] tmp02_22_44;
	wire [WIDTH*2-1+2:0] tmp02_22_45;
	wire [WIDTH*2-1+2:0] tmp02_22_46;
	wire [WIDTH*2-1+2:0] tmp02_22_47;
	wire [WIDTH*2-1+2:0] tmp02_22_48;
	wire [WIDTH*2-1+2:0] tmp02_22_49;
	wire [WIDTH*2-1+2:0] tmp02_22_50;
	wire [WIDTH*2-1+2:0] tmp02_22_51;
	wire [WIDTH*2-1+2:0] tmp02_22_52;
	wire [WIDTH*2-1+2:0] tmp02_22_53;
	wire [WIDTH*2-1+2:0] tmp02_22_54;
	wire [WIDTH*2-1+2:0] tmp02_22_55;
	wire [WIDTH*2-1+2:0] tmp02_22_56;
	wire [WIDTH*2-1+2:0] tmp02_22_57;
	wire [WIDTH*2-1+2:0] tmp02_22_58;
	wire [WIDTH*2-1+2:0] tmp02_22_59;
	wire [WIDTH*2-1+2:0] tmp02_22_60;
	wire [WIDTH*2-1+2:0] tmp02_22_61;
	wire [WIDTH*2-1+2:0] tmp02_22_62;
	wire [WIDTH*2-1+2:0] tmp02_22_63;
	wire [WIDTH*2-1+2:0] tmp02_22_64;
	wire [WIDTH*2-1+2:0] tmp02_22_65;
	wire [WIDTH*2-1+2:0] tmp02_22_66;
	wire [WIDTH*2-1+2:0] tmp02_22_67;
	wire [WIDTH*2-1+2:0] tmp02_22_68;
	wire [WIDTH*2-1+2:0] tmp02_22_69;
	wire [WIDTH*2-1+2:0] tmp02_22_70;
	wire [WIDTH*2-1+2:0] tmp02_22_71;
	wire [WIDTH*2-1+2:0] tmp02_22_72;
	wire [WIDTH*2-1+2:0] tmp02_22_73;
	wire [WIDTH*2-1+2:0] tmp02_22_74;
	wire [WIDTH*2-1+2:0] tmp02_22_75;
	wire [WIDTH*2-1+2:0] tmp02_22_76;
	wire [WIDTH*2-1+2:0] tmp02_22_77;
	wire [WIDTH*2-1+2:0] tmp02_22_78;
	wire [WIDTH*2-1+2:0] tmp02_22_79;
	wire [WIDTH*2-1+2:0] tmp02_22_80;
	wire [WIDTH*2-1+2:0] tmp02_22_81;
	wire [WIDTH*2-1+2:0] tmp02_22_82;
	wire [WIDTH*2-1+2:0] tmp02_22_83;
	wire [WIDTH*2-1+2:0] tmp02_23_0;
	wire [WIDTH*2-1+2:0] tmp02_23_1;
	wire [WIDTH*2-1+2:0] tmp02_23_2;
	wire [WIDTH*2-1+2:0] tmp02_23_3;
	wire [WIDTH*2-1+2:0] tmp02_23_4;
	wire [WIDTH*2-1+2:0] tmp02_23_5;
	wire [WIDTH*2-1+2:0] tmp02_23_6;
	wire [WIDTH*2-1+2:0] tmp02_23_7;
	wire [WIDTH*2-1+2:0] tmp02_23_8;
	wire [WIDTH*2-1+2:0] tmp02_23_9;
	wire [WIDTH*2-1+2:0] tmp02_23_10;
	wire [WIDTH*2-1+2:0] tmp02_23_11;
	wire [WIDTH*2-1+2:0] tmp02_23_12;
	wire [WIDTH*2-1+2:0] tmp02_23_13;
	wire [WIDTH*2-1+2:0] tmp02_23_14;
	wire [WIDTH*2-1+2:0] tmp02_23_15;
	wire [WIDTH*2-1+2:0] tmp02_23_16;
	wire [WIDTH*2-1+2:0] tmp02_23_17;
	wire [WIDTH*2-1+2:0] tmp02_23_18;
	wire [WIDTH*2-1+2:0] tmp02_23_19;
	wire [WIDTH*2-1+2:0] tmp02_23_20;
	wire [WIDTH*2-1+2:0] tmp02_23_21;
	wire [WIDTH*2-1+2:0] tmp02_23_22;
	wire [WIDTH*2-1+2:0] tmp02_23_23;
	wire [WIDTH*2-1+2:0] tmp02_23_24;
	wire [WIDTH*2-1+2:0] tmp02_23_25;
	wire [WIDTH*2-1+2:0] tmp02_23_26;
	wire [WIDTH*2-1+2:0] tmp02_23_27;
	wire [WIDTH*2-1+2:0] tmp02_23_28;
	wire [WIDTH*2-1+2:0] tmp02_23_29;
	wire [WIDTH*2-1+2:0] tmp02_23_30;
	wire [WIDTH*2-1+2:0] tmp02_23_31;
	wire [WIDTH*2-1+2:0] tmp02_23_32;
	wire [WIDTH*2-1+2:0] tmp02_23_33;
	wire [WIDTH*2-1+2:0] tmp02_23_34;
	wire [WIDTH*2-1+2:0] tmp02_23_35;
	wire [WIDTH*2-1+2:0] tmp02_23_36;
	wire [WIDTH*2-1+2:0] tmp02_23_37;
	wire [WIDTH*2-1+2:0] tmp02_23_38;
	wire [WIDTH*2-1+2:0] tmp02_23_39;
	wire [WIDTH*2-1+2:0] tmp02_23_40;
	wire [WIDTH*2-1+2:0] tmp02_23_41;
	wire [WIDTH*2-1+2:0] tmp02_23_42;
	wire [WIDTH*2-1+2:0] tmp02_23_43;
	wire [WIDTH*2-1+2:0] tmp02_23_44;
	wire [WIDTH*2-1+2:0] tmp02_23_45;
	wire [WIDTH*2-1+2:0] tmp02_23_46;
	wire [WIDTH*2-1+2:0] tmp02_23_47;
	wire [WIDTH*2-1+2:0] tmp02_23_48;
	wire [WIDTH*2-1+2:0] tmp02_23_49;
	wire [WIDTH*2-1+2:0] tmp02_23_50;
	wire [WIDTH*2-1+2:0] tmp02_23_51;
	wire [WIDTH*2-1+2:0] tmp02_23_52;
	wire [WIDTH*2-1+2:0] tmp02_23_53;
	wire [WIDTH*2-1+2:0] tmp02_23_54;
	wire [WIDTH*2-1+2:0] tmp02_23_55;
	wire [WIDTH*2-1+2:0] tmp02_23_56;
	wire [WIDTH*2-1+2:0] tmp02_23_57;
	wire [WIDTH*2-1+2:0] tmp02_23_58;
	wire [WIDTH*2-1+2:0] tmp02_23_59;
	wire [WIDTH*2-1+2:0] tmp02_23_60;
	wire [WIDTH*2-1+2:0] tmp02_23_61;
	wire [WIDTH*2-1+2:0] tmp02_23_62;
	wire [WIDTH*2-1+2:0] tmp02_23_63;
	wire [WIDTH*2-1+2:0] tmp02_23_64;
	wire [WIDTH*2-1+2:0] tmp02_23_65;
	wire [WIDTH*2-1+2:0] tmp02_23_66;
	wire [WIDTH*2-1+2:0] tmp02_23_67;
	wire [WIDTH*2-1+2:0] tmp02_23_68;
	wire [WIDTH*2-1+2:0] tmp02_23_69;
	wire [WIDTH*2-1+2:0] tmp02_23_70;
	wire [WIDTH*2-1+2:0] tmp02_23_71;
	wire [WIDTH*2-1+2:0] tmp02_23_72;
	wire [WIDTH*2-1+2:0] tmp02_23_73;
	wire [WIDTH*2-1+2:0] tmp02_23_74;
	wire [WIDTH*2-1+2:0] tmp02_23_75;
	wire [WIDTH*2-1+2:0] tmp02_23_76;
	wire [WIDTH*2-1+2:0] tmp02_23_77;
	wire [WIDTH*2-1+2:0] tmp02_23_78;
	wire [WIDTH*2-1+2:0] tmp02_23_79;
	wire [WIDTH*2-1+2:0] tmp02_23_80;
	wire [WIDTH*2-1+2:0] tmp02_23_81;
	wire [WIDTH*2-1+2:0] tmp02_23_82;
	wire [WIDTH*2-1+2:0] tmp02_23_83;
	wire [WIDTH*2-1+2:0] tmp02_24_0;
	wire [WIDTH*2-1+2:0] tmp02_24_1;
	wire [WIDTH*2-1+2:0] tmp02_24_2;
	wire [WIDTH*2-1+2:0] tmp02_24_3;
	wire [WIDTH*2-1+2:0] tmp02_24_4;
	wire [WIDTH*2-1+2:0] tmp02_24_5;
	wire [WIDTH*2-1+2:0] tmp02_24_6;
	wire [WIDTH*2-1+2:0] tmp02_24_7;
	wire [WIDTH*2-1+2:0] tmp02_24_8;
	wire [WIDTH*2-1+2:0] tmp02_24_9;
	wire [WIDTH*2-1+2:0] tmp02_24_10;
	wire [WIDTH*2-1+2:0] tmp02_24_11;
	wire [WIDTH*2-1+2:0] tmp02_24_12;
	wire [WIDTH*2-1+2:0] tmp02_24_13;
	wire [WIDTH*2-1+2:0] tmp02_24_14;
	wire [WIDTH*2-1+2:0] tmp02_24_15;
	wire [WIDTH*2-1+2:0] tmp02_24_16;
	wire [WIDTH*2-1+2:0] tmp02_24_17;
	wire [WIDTH*2-1+2:0] tmp02_24_18;
	wire [WIDTH*2-1+2:0] tmp02_24_19;
	wire [WIDTH*2-1+2:0] tmp02_24_20;
	wire [WIDTH*2-1+2:0] tmp02_24_21;
	wire [WIDTH*2-1+2:0] tmp02_24_22;
	wire [WIDTH*2-1+2:0] tmp02_24_23;
	wire [WIDTH*2-1+2:0] tmp02_24_24;
	wire [WIDTH*2-1+2:0] tmp02_24_25;
	wire [WIDTH*2-1+2:0] tmp02_24_26;
	wire [WIDTH*2-1+2:0] tmp02_24_27;
	wire [WIDTH*2-1+2:0] tmp02_24_28;
	wire [WIDTH*2-1+2:0] tmp02_24_29;
	wire [WIDTH*2-1+2:0] tmp02_24_30;
	wire [WIDTH*2-1+2:0] tmp02_24_31;
	wire [WIDTH*2-1+2:0] tmp02_24_32;
	wire [WIDTH*2-1+2:0] tmp02_24_33;
	wire [WIDTH*2-1+2:0] tmp02_24_34;
	wire [WIDTH*2-1+2:0] tmp02_24_35;
	wire [WIDTH*2-1+2:0] tmp02_24_36;
	wire [WIDTH*2-1+2:0] tmp02_24_37;
	wire [WIDTH*2-1+2:0] tmp02_24_38;
	wire [WIDTH*2-1+2:0] tmp02_24_39;
	wire [WIDTH*2-1+2:0] tmp02_24_40;
	wire [WIDTH*2-1+2:0] tmp02_24_41;
	wire [WIDTH*2-1+2:0] tmp02_24_42;
	wire [WIDTH*2-1+2:0] tmp02_24_43;
	wire [WIDTH*2-1+2:0] tmp02_24_44;
	wire [WIDTH*2-1+2:0] tmp02_24_45;
	wire [WIDTH*2-1+2:0] tmp02_24_46;
	wire [WIDTH*2-1+2:0] tmp02_24_47;
	wire [WIDTH*2-1+2:0] tmp02_24_48;
	wire [WIDTH*2-1+2:0] tmp02_24_49;
	wire [WIDTH*2-1+2:0] tmp02_24_50;
	wire [WIDTH*2-1+2:0] tmp02_24_51;
	wire [WIDTH*2-1+2:0] tmp02_24_52;
	wire [WIDTH*2-1+2:0] tmp02_24_53;
	wire [WIDTH*2-1+2:0] tmp02_24_54;
	wire [WIDTH*2-1+2:0] tmp02_24_55;
	wire [WIDTH*2-1+2:0] tmp02_24_56;
	wire [WIDTH*2-1+2:0] tmp02_24_57;
	wire [WIDTH*2-1+2:0] tmp02_24_58;
	wire [WIDTH*2-1+2:0] tmp02_24_59;
	wire [WIDTH*2-1+2:0] tmp02_24_60;
	wire [WIDTH*2-1+2:0] tmp02_24_61;
	wire [WIDTH*2-1+2:0] tmp02_24_62;
	wire [WIDTH*2-1+2:0] tmp02_24_63;
	wire [WIDTH*2-1+2:0] tmp02_24_64;
	wire [WIDTH*2-1+2:0] tmp02_24_65;
	wire [WIDTH*2-1+2:0] tmp02_24_66;
	wire [WIDTH*2-1+2:0] tmp02_24_67;
	wire [WIDTH*2-1+2:0] tmp02_24_68;
	wire [WIDTH*2-1+2:0] tmp02_24_69;
	wire [WIDTH*2-1+2:0] tmp02_24_70;
	wire [WIDTH*2-1+2:0] tmp02_24_71;
	wire [WIDTH*2-1+2:0] tmp02_24_72;
	wire [WIDTH*2-1+2:0] tmp02_24_73;
	wire [WIDTH*2-1+2:0] tmp02_24_74;
	wire [WIDTH*2-1+2:0] tmp02_24_75;
	wire [WIDTH*2-1+2:0] tmp02_24_76;
	wire [WIDTH*2-1+2:0] tmp02_24_77;
	wire [WIDTH*2-1+2:0] tmp02_24_78;
	wire [WIDTH*2-1+2:0] tmp02_24_79;
	wire [WIDTH*2-1+2:0] tmp02_24_80;
	wire [WIDTH*2-1+2:0] tmp02_24_81;
	wire [WIDTH*2-1+2:0] tmp02_24_82;
	wire [WIDTH*2-1+2:0] tmp02_24_83;
	wire [WIDTH*2-1+2:0] tmp02_25_0;
	wire [WIDTH*2-1+2:0] tmp02_25_1;
	wire [WIDTH*2-1+2:0] tmp02_25_2;
	wire [WIDTH*2-1+2:0] tmp02_25_3;
	wire [WIDTH*2-1+2:0] tmp02_25_4;
	wire [WIDTH*2-1+2:0] tmp02_25_5;
	wire [WIDTH*2-1+2:0] tmp02_25_6;
	wire [WIDTH*2-1+2:0] tmp02_25_7;
	wire [WIDTH*2-1+2:0] tmp02_25_8;
	wire [WIDTH*2-1+2:0] tmp02_25_9;
	wire [WIDTH*2-1+2:0] tmp02_25_10;
	wire [WIDTH*2-1+2:0] tmp02_25_11;
	wire [WIDTH*2-1+2:0] tmp02_25_12;
	wire [WIDTH*2-1+2:0] tmp02_25_13;
	wire [WIDTH*2-1+2:0] tmp02_25_14;
	wire [WIDTH*2-1+2:0] tmp02_25_15;
	wire [WIDTH*2-1+2:0] tmp02_25_16;
	wire [WIDTH*2-1+2:0] tmp02_25_17;
	wire [WIDTH*2-1+2:0] tmp02_25_18;
	wire [WIDTH*2-1+2:0] tmp02_25_19;
	wire [WIDTH*2-1+2:0] tmp02_25_20;
	wire [WIDTH*2-1+2:0] tmp02_25_21;
	wire [WIDTH*2-1+2:0] tmp02_25_22;
	wire [WIDTH*2-1+2:0] tmp02_25_23;
	wire [WIDTH*2-1+2:0] tmp02_25_24;
	wire [WIDTH*2-1+2:0] tmp02_25_25;
	wire [WIDTH*2-1+2:0] tmp02_25_26;
	wire [WIDTH*2-1+2:0] tmp02_25_27;
	wire [WIDTH*2-1+2:0] tmp02_25_28;
	wire [WIDTH*2-1+2:0] tmp02_25_29;
	wire [WIDTH*2-1+2:0] tmp02_25_30;
	wire [WIDTH*2-1+2:0] tmp02_25_31;
	wire [WIDTH*2-1+2:0] tmp02_25_32;
	wire [WIDTH*2-1+2:0] tmp02_25_33;
	wire [WIDTH*2-1+2:0] tmp02_25_34;
	wire [WIDTH*2-1+2:0] tmp02_25_35;
	wire [WIDTH*2-1+2:0] tmp02_25_36;
	wire [WIDTH*2-1+2:0] tmp02_25_37;
	wire [WIDTH*2-1+2:0] tmp02_25_38;
	wire [WIDTH*2-1+2:0] tmp02_25_39;
	wire [WIDTH*2-1+2:0] tmp02_25_40;
	wire [WIDTH*2-1+2:0] tmp02_25_41;
	wire [WIDTH*2-1+2:0] tmp02_25_42;
	wire [WIDTH*2-1+2:0] tmp02_25_43;
	wire [WIDTH*2-1+2:0] tmp02_25_44;
	wire [WIDTH*2-1+2:0] tmp02_25_45;
	wire [WIDTH*2-1+2:0] tmp02_25_46;
	wire [WIDTH*2-1+2:0] tmp02_25_47;
	wire [WIDTH*2-1+2:0] tmp02_25_48;
	wire [WIDTH*2-1+2:0] tmp02_25_49;
	wire [WIDTH*2-1+2:0] tmp02_25_50;
	wire [WIDTH*2-1+2:0] tmp02_25_51;
	wire [WIDTH*2-1+2:0] tmp02_25_52;
	wire [WIDTH*2-1+2:0] tmp02_25_53;
	wire [WIDTH*2-1+2:0] tmp02_25_54;
	wire [WIDTH*2-1+2:0] tmp02_25_55;
	wire [WIDTH*2-1+2:0] tmp02_25_56;
	wire [WIDTH*2-1+2:0] tmp02_25_57;
	wire [WIDTH*2-1+2:0] tmp02_25_58;
	wire [WIDTH*2-1+2:0] tmp02_25_59;
	wire [WIDTH*2-1+2:0] tmp02_25_60;
	wire [WIDTH*2-1+2:0] tmp02_25_61;
	wire [WIDTH*2-1+2:0] tmp02_25_62;
	wire [WIDTH*2-1+2:0] tmp02_25_63;
	wire [WIDTH*2-1+2:0] tmp02_25_64;
	wire [WIDTH*2-1+2:0] tmp02_25_65;
	wire [WIDTH*2-1+2:0] tmp02_25_66;
	wire [WIDTH*2-1+2:0] tmp02_25_67;
	wire [WIDTH*2-1+2:0] tmp02_25_68;
	wire [WIDTH*2-1+2:0] tmp02_25_69;
	wire [WIDTH*2-1+2:0] tmp02_25_70;
	wire [WIDTH*2-1+2:0] tmp02_25_71;
	wire [WIDTH*2-1+2:0] tmp02_25_72;
	wire [WIDTH*2-1+2:0] tmp02_25_73;
	wire [WIDTH*2-1+2:0] tmp02_25_74;
	wire [WIDTH*2-1+2:0] tmp02_25_75;
	wire [WIDTH*2-1+2:0] tmp02_25_76;
	wire [WIDTH*2-1+2:0] tmp02_25_77;
	wire [WIDTH*2-1+2:0] tmp02_25_78;
	wire [WIDTH*2-1+2:0] tmp02_25_79;
	wire [WIDTH*2-1+2:0] tmp02_25_80;
	wire [WIDTH*2-1+2:0] tmp02_25_81;
	wire [WIDTH*2-1+2:0] tmp02_25_82;
	wire [WIDTH*2-1+2:0] tmp02_25_83;
	wire [WIDTH*2-1+2:0] tmp02_26_0;
	wire [WIDTH*2-1+2:0] tmp02_26_1;
	wire [WIDTH*2-1+2:0] tmp02_26_2;
	wire [WIDTH*2-1+2:0] tmp02_26_3;
	wire [WIDTH*2-1+2:0] tmp02_26_4;
	wire [WIDTH*2-1+2:0] tmp02_26_5;
	wire [WIDTH*2-1+2:0] tmp02_26_6;
	wire [WIDTH*2-1+2:0] tmp02_26_7;
	wire [WIDTH*2-1+2:0] tmp02_26_8;
	wire [WIDTH*2-1+2:0] tmp02_26_9;
	wire [WIDTH*2-1+2:0] tmp02_26_10;
	wire [WIDTH*2-1+2:0] tmp02_26_11;
	wire [WIDTH*2-1+2:0] tmp02_26_12;
	wire [WIDTH*2-1+2:0] tmp02_26_13;
	wire [WIDTH*2-1+2:0] tmp02_26_14;
	wire [WIDTH*2-1+2:0] tmp02_26_15;
	wire [WIDTH*2-1+2:0] tmp02_26_16;
	wire [WIDTH*2-1+2:0] tmp02_26_17;
	wire [WIDTH*2-1+2:0] tmp02_26_18;
	wire [WIDTH*2-1+2:0] tmp02_26_19;
	wire [WIDTH*2-1+2:0] tmp02_26_20;
	wire [WIDTH*2-1+2:0] tmp02_26_21;
	wire [WIDTH*2-1+2:0] tmp02_26_22;
	wire [WIDTH*2-1+2:0] tmp02_26_23;
	wire [WIDTH*2-1+2:0] tmp02_26_24;
	wire [WIDTH*2-1+2:0] tmp02_26_25;
	wire [WIDTH*2-1+2:0] tmp02_26_26;
	wire [WIDTH*2-1+2:0] tmp02_26_27;
	wire [WIDTH*2-1+2:0] tmp02_26_28;
	wire [WIDTH*2-1+2:0] tmp02_26_29;
	wire [WIDTH*2-1+2:0] tmp02_26_30;
	wire [WIDTH*2-1+2:0] tmp02_26_31;
	wire [WIDTH*2-1+2:0] tmp02_26_32;
	wire [WIDTH*2-1+2:0] tmp02_26_33;
	wire [WIDTH*2-1+2:0] tmp02_26_34;
	wire [WIDTH*2-1+2:0] tmp02_26_35;
	wire [WIDTH*2-1+2:0] tmp02_26_36;
	wire [WIDTH*2-1+2:0] tmp02_26_37;
	wire [WIDTH*2-1+2:0] tmp02_26_38;
	wire [WIDTH*2-1+2:0] tmp02_26_39;
	wire [WIDTH*2-1+2:0] tmp02_26_40;
	wire [WIDTH*2-1+2:0] tmp02_26_41;
	wire [WIDTH*2-1+2:0] tmp02_26_42;
	wire [WIDTH*2-1+2:0] tmp02_26_43;
	wire [WIDTH*2-1+2:0] tmp02_26_44;
	wire [WIDTH*2-1+2:0] tmp02_26_45;
	wire [WIDTH*2-1+2:0] tmp02_26_46;
	wire [WIDTH*2-1+2:0] tmp02_26_47;
	wire [WIDTH*2-1+2:0] tmp02_26_48;
	wire [WIDTH*2-1+2:0] tmp02_26_49;
	wire [WIDTH*2-1+2:0] tmp02_26_50;
	wire [WIDTH*2-1+2:0] tmp02_26_51;
	wire [WIDTH*2-1+2:0] tmp02_26_52;
	wire [WIDTH*2-1+2:0] tmp02_26_53;
	wire [WIDTH*2-1+2:0] tmp02_26_54;
	wire [WIDTH*2-1+2:0] tmp02_26_55;
	wire [WIDTH*2-1+2:0] tmp02_26_56;
	wire [WIDTH*2-1+2:0] tmp02_26_57;
	wire [WIDTH*2-1+2:0] tmp02_26_58;
	wire [WIDTH*2-1+2:0] tmp02_26_59;
	wire [WIDTH*2-1+2:0] tmp02_26_60;
	wire [WIDTH*2-1+2:0] tmp02_26_61;
	wire [WIDTH*2-1+2:0] tmp02_26_62;
	wire [WIDTH*2-1+2:0] tmp02_26_63;
	wire [WIDTH*2-1+2:0] tmp02_26_64;
	wire [WIDTH*2-1+2:0] tmp02_26_65;
	wire [WIDTH*2-1+2:0] tmp02_26_66;
	wire [WIDTH*2-1+2:0] tmp02_26_67;
	wire [WIDTH*2-1+2:0] tmp02_26_68;
	wire [WIDTH*2-1+2:0] tmp02_26_69;
	wire [WIDTH*2-1+2:0] tmp02_26_70;
	wire [WIDTH*2-1+2:0] tmp02_26_71;
	wire [WIDTH*2-1+2:0] tmp02_26_72;
	wire [WIDTH*2-1+2:0] tmp02_26_73;
	wire [WIDTH*2-1+2:0] tmp02_26_74;
	wire [WIDTH*2-1+2:0] tmp02_26_75;
	wire [WIDTH*2-1+2:0] tmp02_26_76;
	wire [WIDTH*2-1+2:0] tmp02_26_77;
	wire [WIDTH*2-1+2:0] tmp02_26_78;
	wire [WIDTH*2-1+2:0] tmp02_26_79;
	wire [WIDTH*2-1+2:0] tmp02_26_80;
	wire [WIDTH*2-1+2:0] tmp02_26_81;
	wire [WIDTH*2-1+2:0] tmp02_26_82;
	wire [WIDTH*2-1+2:0] tmp02_26_83;
	wire [WIDTH*2-1+2:0] tmp02_27_0;
	wire [WIDTH*2-1+2:0] tmp02_27_1;
	wire [WIDTH*2-1+2:0] tmp02_27_2;
	wire [WIDTH*2-1+2:0] tmp02_27_3;
	wire [WIDTH*2-1+2:0] tmp02_27_4;
	wire [WIDTH*2-1+2:0] tmp02_27_5;
	wire [WIDTH*2-1+2:0] tmp02_27_6;
	wire [WIDTH*2-1+2:0] tmp02_27_7;
	wire [WIDTH*2-1+2:0] tmp02_27_8;
	wire [WIDTH*2-1+2:0] tmp02_27_9;
	wire [WIDTH*2-1+2:0] tmp02_27_10;
	wire [WIDTH*2-1+2:0] tmp02_27_11;
	wire [WIDTH*2-1+2:0] tmp02_27_12;
	wire [WIDTH*2-1+2:0] tmp02_27_13;
	wire [WIDTH*2-1+2:0] tmp02_27_14;
	wire [WIDTH*2-1+2:0] tmp02_27_15;
	wire [WIDTH*2-1+2:0] tmp02_27_16;
	wire [WIDTH*2-1+2:0] tmp02_27_17;
	wire [WIDTH*2-1+2:0] tmp02_27_18;
	wire [WIDTH*2-1+2:0] tmp02_27_19;
	wire [WIDTH*2-1+2:0] tmp02_27_20;
	wire [WIDTH*2-1+2:0] tmp02_27_21;
	wire [WIDTH*2-1+2:0] tmp02_27_22;
	wire [WIDTH*2-1+2:0] tmp02_27_23;
	wire [WIDTH*2-1+2:0] tmp02_27_24;
	wire [WIDTH*2-1+2:0] tmp02_27_25;
	wire [WIDTH*2-1+2:0] tmp02_27_26;
	wire [WIDTH*2-1+2:0] tmp02_27_27;
	wire [WIDTH*2-1+2:0] tmp02_27_28;
	wire [WIDTH*2-1+2:0] tmp02_27_29;
	wire [WIDTH*2-1+2:0] tmp02_27_30;
	wire [WIDTH*2-1+2:0] tmp02_27_31;
	wire [WIDTH*2-1+2:0] tmp02_27_32;
	wire [WIDTH*2-1+2:0] tmp02_27_33;
	wire [WIDTH*2-1+2:0] tmp02_27_34;
	wire [WIDTH*2-1+2:0] tmp02_27_35;
	wire [WIDTH*2-1+2:0] tmp02_27_36;
	wire [WIDTH*2-1+2:0] tmp02_27_37;
	wire [WIDTH*2-1+2:0] tmp02_27_38;
	wire [WIDTH*2-1+2:0] tmp02_27_39;
	wire [WIDTH*2-1+2:0] tmp02_27_40;
	wire [WIDTH*2-1+2:0] tmp02_27_41;
	wire [WIDTH*2-1+2:0] tmp02_27_42;
	wire [WIDTH*2-1+2:0] tmp02_27_43;
	wire [WIDTH*2-1+2:0] tmp02_27_44;
	wire [WIDTH*2-1+2:0] tmp02_27_45;
	wire [WIDTH*2-1+2:0] tmp02_27_46;
	wire [WIDTH*2-1+2:0] tmp02_27_47;
	wire [WIDTH*2-1+2:0] tmp02_27_48;
	wire [WIDTH*2-1+2:0] tmp02_27_49;
	wire [WIDTH*2-1+2:0] tmp02_27_50;
	wire [WIDTH*2-1+2:0] tmp02_27_51;
	wire [WIDTH*2-1+2:0] tmp02_27_52;
	wire [WIDTH*2-1+2:0] tmp02_27_53;
	wire [WIDTH*2-1+2:0] tmp02_27_54;
	wire [WIDTH*2-1+2:0] tmp02_27_55;
	wire [WIDTH*2-1+2:0] tmp02_27_56;
	wire [WIDTH*2-1+2:0] tmp02_27_57;
	wire [WIDTH*2-1+2:0] tmp02_27_58;
	wire [WIDTH*2-1+2:0] tmp02_27_59;
	wire [WIDTH*2-1+2:0] tmp02_27_60;
	wire [WIDTH*2-1+2:0] tmp02_27_61;
	wire [WIDTH*2-1+2:0] tmp02_27_62;
	wire [WIDTH*2-1+2:0] tmp02_27_63;
	wire [WIDTH*2-1+2:0] tmp02_27_64;
	wire [WIDTH*2-1+2:0] tmp02_27_65;
	wire [WIDTH*2-1+2:0] tmp02_27_66;
	wire [WIDTH*2-1+2:0] tmp02_27_67;
	wire [WIDTH*2-1+2:0] tmp02_27_68;
	wire [WIDTH*2-1+2:0] tmp02_27_69;
	wire [WIDTH*2-1+2:0] tmp02_27_70;
	wire [WIDTH*2-1+2:0] tmp02_27_71;
	wire [WIDTH*2-1+2:0] tmp02_27_72;
	wire [WIDTH*2-1+2:0] tmp02_27_73;
	wire [WIDTH*2-1+2:0] tmp02_27_74;
	wire [WIDTH*2-1+2:0] tmp02_27_75;
	wire [WIDTH*2-1+2:0] tmp02_27_76;
	wire [WIDTH*2-1+2:0] tmp02_27_77;
	wire [WIDTH*2-1+2:0] tmp02_27_78;
	wire [WIDTH*2-1+2:0] tmp02_27_79;
	wire [WIDTH*2-1+2:0] tmp02_27_80;
	wire [WIDTH*2-1+2:0] tmp02_27_81;
	wire [WIDTH*2-1+2:0] tmp02_27_82;
	wire [WIDTH*2-1+2:0] tmp02_27_83;
	wire [WIDTH*2-1+2:0] tmp02_28_0;
	wire [WIDTH*2-1+2:0] tmp02_28_1;
	wire [WIDTH*2-1+2:0] tmp02_28_2;
	wire [WIDTH*2-1+2:0] tmp02_28_3;
	wire [WIDTH*2-1+2:0] tmp02_28_4;
	wire [WIDTH*2-1+2:0] tmp02_28_5;
	wire [WIDTH*2-1+2:0] tmp02_28_6;
	wire [WIDTH*2-1+2:0] tmp02_28_7;
	wire [WIDTH*2-1+2:0] tmp02_28_8;
	wire [WIDTH*2-1+2:0] tmp02_28_9;
	wire [WIDTH*2-1+2:0] tmp02_28_10;
	wire [WIDTH*2-1+2:0] tmp02_28_11;
	wire [WIDTH*2-1+2:0] tmp02_28_12;
	wire [WIDTH*2-1+2:0] tmp02_28_13;
	wire [WIDTH*2-1+2:0] tmp02_28_14;
	wire [WIDTH*2-1+2:0] tmp02_28_15;
	wire [WIDTH*2-1+2:0] tmp02_28_16;
	wire [WIDTH*2-1+2:0] tmp02_28_17;
	wire [WIDTH*2-1+2:0] tmp02_28_18;
	wire [WIDTH*2-1+2:0] tmp02_28_19;
	wire [WIDTH*2-1+2:0] tmp02_28_20;
	wire [WIDTH*2-1+2:0] tmp02_28_21;
	wire [WIDTH*2-1+2:0] tmp02_28_22;
	wire [WIDTH*2-1+2:0] tmp02_28_23;
	wire [WIDTH*2-1+2:0] tmp02_28_24;
	wire [WIDTH*2-1+2:0] tmp02_28_25;
	wire [WIDTH*2-1+2:0] tmp02_28_26;
	wire [WIDTH*2-1+2:0] tmp02_28_27;
	wire [WIDTH*2-1+2:0] tmp02_28_28;
	wire [WIDTH*2-1+2:0] tmp02_28_29;
	wire [WIDTH*2-1+2:0] tmp02_28_30;
	wire [WIDTH*2-1+2:0] tmp02_28_31;
	wire [WIDTH*2-1+2:0] tmp02_28_32;
	wire [WIDTH*2-1+2:0] tmp02_28_33;
	wire [WIDTH*2-1+2:0] tmp02_28_34;
	wire [WIDTH*2-1+2:0] tmp02_28_35;
	wire [WIDTH*2-1+2:0] tmp02_28_36;
	wire [WIDTH*2-1+2:0] tmp02_28_37;
	wire [WIDTH*2-1+2:0] tmp02_28_38;
	wire [WIDTH*2-1+2:0] tmp02_28_39;
	wire [WIDTH*2-1+2:0] tmp02_28_40;
	wire [WIDTH*2-1+2:0] tmp02_28_41;
	wire [WIDTH*2-1+2:0] tmp02_28_42;
	wire [WIDTH*2-1+2:0] tmp02_28_43;
	wire [WIDTH*2-1+2:0] tmp02_28_44;
	wire [WIDTH*2-1+2:0] tmp02_28_45;
	wire [WIDTH*2-1+2:0] tmp02_28_46;
	wire [WIDTH*2-1+2:0] tmp02_28_47;
	wire [WIDTH*2-1+2:0] tmp02_28_48;
	wire [WIDTH*2-1+2:0] tmp02_28_49;
	wire [WIDTH*2-1+2:0] tmp02_28_50;
	wire [WIDTH*2-1+2:0] tmp02_28_51;
	wire [WIDTH*2-1+2:0] tmp02_28_52;
	wire [WIDTH*2-1+2:0] tmp02_28_53;
	wire [WIDTH*2-1+2:0] tmp02_28_54;
	wire [WIDTH*2-1+2:0] tmp02_28_55;
	wire [WIDTH*2-1+2:0] tmp02_28_56;
	wire [WIDTH*2-1+2:0] tmp02_28_57;
	wire [WIDTH*2-1+2:0] tmp02_28_58;
	wire [WIDTH*2-1+2:0] tmp02_28_59;
	wire [WIDTH*2-1+2:0] tmp02_28_60;
	wire [WIDTH*2-1+2:0] tmp02_28_61;
	wire [WIDTH*2-1+2:0] tmp02_28_62;
	wire [WIDTH*2-1+2:0] tmp02_28_63;
	wire [WIDTH*2-1+2:0] tmp02_28_64;
	wire [WIDTH*2-1+2:0] tmp02_28_65;
	wire [WIDTH*2-1+2:0] tmp02_28_66;
	wire [WIDTH*2-1+2:0] tmp02_28_67;
	wire [WIDTH*2-1+2:0] tmp02_28_68;
	wire [WIDTH*2-1+2:0] tmp02_28_69;
	wire [WIDTH*2-1+2:0] tmp02_28_70;
	wire [WIDTH*2-1+2:0] tmp02_28_71;
	wire [WIDTH*2-1+2:0] tmp02_28_72;
	wire [WIDTH*2-1+2:0] tmp02_28_73;
	wire [WIDTH*2-1+2:0] tmp02_28_74;
	wire [WIDTH*2-1+2:0] tmp02_28_75;
	wire [WIDTH*2-1+2:0] tmp02_28_76;
	wire [WIDTH*2-1+2:0] tmp02_28_77;
	wire [WIDTH*2-1+2:0] tmp02_28_78;
	wire [WIDTH*2-1+2:0] tmp02_28_79;
	wire [WIDTH*2-1+2:0] tmp02_28_80;
	wire [WIDTH*2-1+2:0] tmp02_28_81;
	wire [WIDTH*2-1+2:0] tmp02_28_82;
	wire [WIDTH*2-1+2:0] tmp02_28_83;
	wire [WIDTH*2-1+2:0] tmp02_29_0;
	wire [WIDTH*2-1+2:0] tmp02_29_1;
	wire [WIDTH*2-1+2:0] tmp02_29_2;
	wire [WIDTH*2-1+2:0] tmp02_29_3;
	wire [WIDTH*2-1+2:0] tmp02_29_4;
	wire [WIDTH*2-1+2:0] tmp02_29_5;
	wire [WIDTH*2-1+2:0] tmp02_29_6;
	wire [WIDTH*2-1+2:0] tmp02_29_7;
	wire [WIDTH*2-1+2:0] tmp02_29_8;
	wire [WIDTH*2-1+2:0] tmp02_29_9;
	wire [WIDTH*2-1+2:0] tmp02_29_10;
	wire [WIDTH*2-1+2:0] tmp02_29_11;
	wire [WIDTH*2-1+2:0] tmp02_29_12;
	wire [WIDTH*2-1+2:0] tmp02_29_13;
	wire [WIDTH*2-1+2:0] tmp02_29_14;
	wire [WIDTH*2-1+2:0] tmp02_29_15;
	wire [WIDTH*2-1+2:0] tmp02_29_16;
	wire [WIDTH*2-1+2:0] tmp02_29_17;
	wire [WIDTH*2-1+2:0] tmp02_29_18;
	wire [WIDTH*2-1+2:0] tmp02_29_19;
	wire [WIDTH*2-1+2:0] tmp02_29_20;
	wire [WIDTH*2-1+2:0] tmp02_29_21;
	wire [WIDTH*2-1+2:0] tmp02_29_22;
	wire [WIDTH*2-1+2:0] tmp02_29_23;
	wire [WIDTH*2-1+2:0] tmp02_29_24;
	wire [WIDTH*2-1+2:0] tmp02_29_25;
	wire [WIDTH*2-1+2:0] tmp02_29_26;
	wire [WIDTH*2-1+2:0] tmp02_29_27;
	wire [WIDTH*2-1+2:0] tmp02_29_28;
	wire [WIDTH*2-1+2:0] tmp02_29_29;
	wire [WIDTH*2-1+2:0] tmp02_29_30;
	wire [WIDTH*2-1+2:0] tmp02_29_31;
	wire [WIDTH*2-1+2:0] tmp02_29_32;
	wire [WIDTH*2-1+2:0] tmp02_29_33;
	wire [WIDTH*2-1+2:0] tmp02_29_34;
	wire [WIDTH*2-1+2:0] tmp02_29_35;
	wire [WIDTH*2-1+2:0] tmp02_29_36;
	wire [WIDTH*2-1+2:0] tmp02_29_37;
	wire [WIDTH*2-1+2:0] tmp02_29_38;
	wire [WIDTH*2-1+2:0] tmp02_29_39;
	wire [WIDTH*2-1+2:0] tmp02_29_40;
	wire [WIDTH*2-1+2:0] tmp02_29_41;
	wire [WIDTH*2-1+2:0] tmp02_29_42;
	wire [WIDTH*2-1+2:0] tmp02_29_43;
	wire [WIDTH*2-1+2:0] tmp02_29_44;
	wire [WIDTH*2-1+2:0] tmp02_29_45;
	wire [WIDTH*2-1+2:0] tmp02_29_46;
	wire [WIDTH*2-1+2:0] tmp02_29_47;
	wire [WIDTH*2-1+2:0] tmp02_29_48;
	wire [WIDTH*2-1+2:0] tmp02_29_49;
	wire [WIDTH*2-1+2:0] tmp02_29_50;
	wire [WIDTH*2-1+2:0] tmp02_29_51;
	wire [WIDTH*2-1+2:0] tmp02_29_52;
	wire [WIDTH*2-1+2:0] tmp02_29_53;
	wire [WIDTH*2-1+2:0] tmp02_29_54;
	wire [WIDTH*2-1+2:0] tmp02_29_55;
	wire [WIDTH*2-1+2:0] tmp02_29_56;
	wire [WIDTH*2-1+2:0] tmp02_29_57;
	wire [WIDTH*2-1+2:0] tmp02_29_58;
	wire [WIDTH*2-1+2:0] tmp02_29_59;
	wire [WIDTH*2-1+2:0] tmp02_29_60;
	wire [WIDTH*2-1+2:0] tmp02_29_61;
	wire [WIDTH*2-1+2:0] tmp02_29_62;
	wire [WIDTH*2-1+2:0] tmp02_29_63;
	wire [WIDTH*2-1+2:0] tmp02_29_64;
	wire [WIDTH*2-1+2:0] tmp02_29_65;
	wire [WIDTH*2-1+2:0] tmp02_29_66;
	wire [WIDTH*2-1+2:0] tmp02_29_67;
	wire [WIDTH*2-1+2:0] tmp02_29_68;
	wire [WIDTH*2-1+2:0] tmp02_29_69;
	wire [WIDTH*2-1+2:0] tmp02_29_70;
	wire [WIDTH*2-1+2:0] tmp02_29_71;
	wire [WIDTH*2-1+2:0] tmp02_29_72;
	wire [WIDTH*2-1+2:0] tmp02_29_73;
	wire [WIDTH*2-1+2:0] tmp02_29_74;
	wire [WIDTH*2-1+2:0] tmp02_29_75;
	wire [WIDTH*2-1+2:0] tmp02_29_76;
	wire [WIDTH*2-1+2:0] tmp02_29_77;
	wire [WIDTH*2-1+2:0] tmp02_29_78;
	wire [WIDTH*2-1+2:0] tmp02_29_79;
	wire [WIDTH*2-1+2:0] tmp02_29_80;
	wire [WIDTH*2-1+2:0] tmp02_29_81;
	wire [WIDTH*2-1+2:0] tmp02_29_82;
	wire [WIDTH*2-1+2:0] tmp02_29_83;
	wire [WIDTH*2-1+2:0] tmp02_30_0;
	wire [WIDTH*2-1+2:0] tmp02_30_1;
	wire [WIDTH*2-1+2:0] tmp02_30_2;
	wire [WIDTH*2-1+2:0] tmp02_30_3;
	wire [WIDTH*2-1+2:0] tmp02_30_4;
	wire [WIDTH*2-1+2:0] tmp02_30_5;
	wire [WIDTH*2-1+2:0] tmp02_30_6;
	wire [WIDTH*2-1+2:0] tmp02_30_7;
	wire [WIDTH*2-1+2:0] tmp02_30_8;
	wire [WIDTH*2-1+2:0] tmp02_30_9;
	wire [WIDTH*2-1+2:0] tmp02_30_10;
	wire [WIDTH*2-1+2:0] tmp02_30_11;
	wire [WIDTH*2-1+2:0] tmp02_30_12;
	wire [WIDTH*2-1+2:0] tmp02_30_13;
	wire [WIDTH*2-1+2:0] tmp02_30_14;
	wire [WIDTH*2-1+2:0] tmp02_30_15;
	wire [WIDTH*2-1+2:0] tmp02_30_16;
	wire [WIDTH*2-1+2:0] tmp02_30_17;
	wire [WIDTH*2-1+2:0] tmp02_30_18;
	wire [WIDTH*2-1+2:0] tmp02_30_19;
	wire [WIDTH*2-1+2:0] tmp02_30_20;
	wire [WIDTH*2-1+2:0] tmp02_30_21;
	wire [WIDTH*2-1+2:0] tmp02_30_22;
	wire [WIDTH*2-1+2:0] tmp02_30_23;
	wire [WIDTH*2-1+2:0] tmp02_30_24;
	wire [WIDTH*2-1+2:0] tmp02_30_25;
	wire [WIDTH*2-1+2:0] tmp02_30_26;
	wire [WIDTH*2-1+2:0] tmp02_30_27;
	wire [WIDTH*2-1+2:0] tmp02_30_28;
	wire [WIDTH*2-1+2:0] tmp02_30_29;
	wire [WIDTH*2-1+2:0] tmp02_30_30;
	wire [WIDTH*2-1+2:0] tmp02_30_31;
	wire [WIDTH*2-1+2:0] tmp02_30_32;
	wire [WIDTH*2-1+2:0] tmp02_30_33;
	wire [WIDTH*2-1+2:0] tmp02_30_34;
	wire [WIDTH*2-1+2:0] tmp02_30_35;
	wire [WIDTH*2-1+2:0] tmp02_30_36;
	wire [WIDTH*2-1+2:0] tmp02_30_37;
	wire [WIDTH*2-1+2:0] tmp02_30_38;
	wire [WIDTH*2-1+2:0] tmp02_30_39;
	wire [WIDTH*2-1+2:0] tmp02_30_40;
	wire [WIDTH*2-1+2:0] tmp02_30_41;
	wire [WIDTH*2-1+2:0] tmp02_30_42;
	wire [WIDTH*2-1+2:0] tmp02_30_43;
	wire [WIDTH*2-1+2:0] tmp02_30_44;
	wire [WIDTH*2-1+2:0] tmp02_30_45;
	wire [WIDTH*2-1+2:0] tmp02_30_46;
	wire [WIDTH*2-1+2:0] tmp02_30_47;
	wire [WIDTH*2-1+2:0] tmp02_30_48;
	wire [WIDTH*2-1+2:0] tmp02_30_49;
	wire [WIDTH*2-1+2:0] tmp02_30_50;
	wire [WIDTH*2-1+2:0] tmp02_30_51;
	wire [WIDTH*2-1+2:0] tmp02_30_52;
	wire [WIDTH*2-1+2:0] tmp02_30_53;
	wire [WIDTH*2-1+2:0] tmp02_30_54;
	wire [WIDTH*2-1+2:0] tmp02_30_55;
	wire [WIDTH*2-1+2:0] tmp02_30_56;
	wire [WIDTH*2-1+2:0] tmp02_30_57;
	wire [WIDTH*2-1+2:0] tmp02_30_58;
	wire [WIDTH*2-1+2:0] tmp02_30_59;
	wire [WIDTH*2-1+2:0] tmp02_30_60;
	wire [WIDTH*2-1+2:0] tmp02_30_61;
	wire [WIDTH*2-1+2:0] tmp02_30_62;
	wire [WIDTH*2-1+2:0] tmp02_30_63;
	wire [WIDTH*2-1+2:0] tmp02_30_64;
	wire [WIDTH*2-1+2:0] tmp02_30_65;
	wire [WIDTH*2-1+2:0] tmp02_30_66;
	wire [WIDTH*2-1+2:0] tmp02_30_67;
	wire [WIDTH*2-1+2:0] tmp02_30_68;
	wire [WIDTH*2-1+2:0] tmp02_30_69;
	wire [WIDTH*2-1+2:0] tmp02_30_70;
	wire [WIDTH*2-1+2:0] tmp02_30_71;
	wire [WIDTH*2-1+2:0] tmp02_30_72;
	wire [WIDTH*2-1+2:0] tmp02_30_73;
	wire [WIDTH*2-1+2:0] tmp02_30_74;
	wire [WIDTH*2-1+2:0] tmp02_30_75;
	wire [WIDTH*2-1+2:0] tmp02_30_76;
	wire [WIDTH*2-1+2:0] tmp02_30_77;
	wire [WIDTH*2-1+2:0] tmp02_30_78;
	wire [WIDTH*2-1+2:0] tmp02_30_79;
	wire [WIDTH*2-1+2:0] tmp02_30_80;
	wire [WIDTH*2-1+2:0] tmp02_30_81;
	wire [WIDTH*2-1+2:0] tmp02_30_82;
	wire [WIDTH*2-1+2:0] tmp02_30_83;
	wire [WIDTH*2-1+2:0] tmp02_31_0;
	wire [WIDTH*2-1+2:0] tmp02_31_1;
	wire [WIDTH*2-1+2:0] tmp02_31_2;
	wire [WIDTH*2-1+2:0] tmp02_31_3;
	wire [WIDTH*2-1+2:0] tmp02_31_4;
	wire [WIDTH*2-1+2:0] tmp02_31_5;
	wire [WIDTH*2-1+2:0] tmp02_31_6;
	wire [WIDTH*2-1+2:0] tmp02_31_7;
	wire [WIDTH*2-1+2:0] tmp02_31_8;
	wire [WIDTH*2-1+2:0] tmp02_31_9;
	wire [WIDTH*2-1+2:0] tmp02_31_10;
	wire [WIDTH*2-1+2:0] tmp02_31_11;
	wire [WIDTH*2-1+2:0] tmp02_31_12;
	wire [WIDTH*2-1+2:0] tmp02_31_13;
	wire [WIDTH*2-1+2:0] tmp02_31_14;
	wire [WIDTH*2-1+2:0] tmp02_31_15;
	wire [WIDTH*2-1+2:0] tmp02_31_16;
	wire [WIDTH*2-1+2:0] tmp02_31_17;
	wire [WIDTH*2-1+2:0] tmp02_31_18;
	wire [WIDTH*2-1+2:0] tmp02_31_19;
	wire [WIDTH*2-1+2:0] tmp02_31_20;
	wire [WIDTH*2-1+2:0] tmp02_31_21;
	wire [WIDTH*2-1+2:0] tmp02_31_22;
	wire [WIDTH*2-1+2:0] tmp02_31_23;
	wire [WIDTH*2-1+2:0] tmp02_31_24;
	wire [WIDTH*2-1+2:0] tmp02_31_25;
	wire [WIDTH*2-1+2:0] tmp02_31_26;
	wire [WIDTH*2-1+2:0] tmp02_31_27;
	wire [WIDTH*2-1+2:0] tmp02_31_28;
	wire [WIDTH*2-1+2:0] tmp02_31_29;
	wire [WIDTH*2-1+2:0] tmp02_31_30;
	wire [WIDTH*2-1+2:0] tmp02_31_31;
	wire [WIDTH*2-1+2:0] tmp02_31_32;
	wire [WIDTH*2-1+2:0] tmp02_31_33;
	wire [WIDTH*2-1+2:0] tmp02_31_34;
	wire [WIDTH*2-1+2:0] tmp02_31_35;
	wire [WIDTH*2-1+2:0] tmp02_31_36;
	wire [WIDTH*2-1+2:0] tmp02_31_37;
	wire [WIDTH*2-1+2:0] tmp02_31_38;
	wire [WIDTH*2-1+2:0] tmp02_31_39;
	wire [WIDTH*2-1+2:0] tmp02_31_40;
	wire [WIDTH*2-1+2:0] tmp02_31_41;
	wire [WIDTH*2-1+2:0] tmp02_31_42;
	wire [WIDTH*2-1+2:0] tmp02_31_43;
	wire [WIDTH*2-1+2:0] tmp02_31_44;
	wire [WIDTH*2-1+2:0] tmp02_31_45;
	wire [WIDTH*2-1+2:0] tmp02_31_46;
	wire [WIDTH*2-1+2:0] tmp02_31_47;
	wire [WIDTH*2-1+2:0] tmp02_31_48;
	wire [WIDTH*2-1+2:0] tmp02_31_49;
	wire [WIDTH*2-1+2:0] tmp02_31_50;
	wire [WIDTH*2-1+2:0] tmp02_31_51;
	wire [WIDTH*2-1+2:0] tmp02_31_52;
	wire [WIDTH*2-1+2:0] tmp02_31_53;
	wire [WIDTH*2-1+2:0] tmp02_31_54;
	wire [WIDTH*2-1+2:0] tmp02_31_55;
	wire [WIDTH*2-1+2:0] tmp02_31_56;
	wire [WIDTH*2-1+2:0] tmp02_31_57;
	wire [WIDTH*2-1+2:0] tmp02_31_58;
	wire [WIDTH*2-1+2:0] tmp02_31_59;
	wire [WIDTH*2-1+2:0] tmp02_31_60;
	wire [WIDTH*2-1+2:0] tmp02_31_61;
	wire [WIDTH*2-1+2:0] tmp02_31_62;
	wire [WIDTH*2-1+2:0] tmp02_31_63;
	wire [WIDTH*2-1+2:0] tmp02_31_64;
	wire [WIDTH*2-1+2:0] tmp02_31_65;
	wire [WIDTH*2-1+2:0] tmp02_31_66;
	wire [WIDTH*2-1+2:0] tmp02_31_67;
	wire [WIDTH*2-1+2:0] tmp02_31_68;
	wire [WIDTH*2-1+2:0] tmp02_31_69;
	wire [WIDTH*2-1+2:0] tmp02_31_70;
	wire [WIDTH*2-1+2:0] tmp02_31_71;
	wire [WIDTH*2-1+2:0] tmp02_31_72;
	wire [WIDTH*2-1+2:0] tmp02_31_73;
	wire [WIDTH*2-1+2:0] tmp02_31_74;
	wire [WIDTH*2-1+2:0] tmp02_31_75;
	wire [WIDTH*2-1+2:0] tmp02_31_76;
	wire [WIDTH*2-1+2:0] tmp02_31_77;
	wire [WIDTH*2-1+2:0] tmp02_31_78;
	wire [WIDTH*2-1+2:0] tmp02_31_79;
	wire [WIDTH*2-1+2:0] tmp02_31_80;
	wire [WIDTH*2-1+2:0] tmp02_31_81;
	wire [WIDTH*2-1+2:0] tmp02_31_82;
	wire [WIDTH*2-1+2:0] tmp02_31_83;
	wire [WIDTH*2-1+3:0] tmp03_0_0;
	wire [WIDTH*2-1+3:0] tmp03_0_1;
	wire [WIDTH*2-1+3:0] tmp03_0_2;
	wire [WIDTH*2-1+3:0] tmp03_0_3;
	wire [WIDTH*2-1+3:0] tmp03_0_4;
	wire [WIDTH*2-1+3:0] tmp03_0_5;
	wire [WIDTH*2-1+3:0] tmp03_0_6;
	wire [WIDTH*2-1+3:0] tmp03_0_7;
	wire [WIDTH*2-1+3:0] tmp03_0_8;
	wire [WIDTH*2-1+3:0] tmp03_0_9;
	wire [WIDTH*2-1+3:0] tmp03_0_10;
	wire [WIDTH*2-1+3:0] tmp03_0_11;
	wire [WIDTH*2-1+3:0] tmp03_0_12;
	wire [WIDTH*2-1+3:0] tmp03_0_13;
	wire [WIDTH*2-1+3:0] tmp03_0_14;
	wire [WIDTH*2-1+3:0] tmp03_0_15;
	wire [WIDTH*2-1+3:0] tmp03_0_16;
	wire [WIDTH*2-1+3:0] tmp03_0_17;
	wire [WIDTH*2-1+3:0] tmp03_0_18;
	wire [WIDTH*2-1+3:0] tmp03_0_19;
	wire [WIDTH*2-1+3:0] tmp03_0_20;
	wire [WIDTH*2-1+3:0] tmp03_0_21;
	wire [WIDTH*2-1+3:0] tmp03_0_22;
	wire [WIDTH*2-1+3:0] tmp03_0_23;
	wire [WIDTH*2-1+3:0] tmp03_0_24;
	wire [WIDTH*2-1+3:0] tmp03_0_25;
	wire [WIDTH*2-1+3:0] tmp03_0_26;
	wire [WIDTH*2-1+3:0] tmp03_0_27;
	wire [WIDTH*2-1+3:0] tmp03_0_28;
	wire [WIDTH*2-1+3:0] tmp03_0_29;
	wire [WIDTH*2-1+3:0] tmp03_0_30;
	wire [WIDTH*2-1+3:0] tmp03_0_31;
	wire [WIDTH*2-1+3:0] tmp03_0_32;
	wire [WIDTH*2-1+3:0] tmp03_0_33;
	wire [WIDTH*2-1+3:0] tmp03_0_34;
	wire [WIDTH*2-1+3:0] tmp03_0_35;
	wire [WIDTH*2-1+3:0] tmp03_0_36;
	wire [WIDTH*2-1+3:0] tmp03_0_37;
	wire [WIDTH*2-1+3:0] tmp03_0_38;
	wire [WIDTH*2-1+3:0] tmp03_0_39;
	wire [WIDTH*2-1+3:0] tmp03_0_40;
	wire [WIDTH*2-1+3:0] tmp03_0_41;
	wire [WIDTH*2-1+3:0] tmp03_0_42;
	wire [WIDTH*2-1+3:0] tmp03_0_43;
	wire [WIDTH*2-1+3:0] tmp03_0_44;
	wire [WIDTH*2-1+3:0] tmp03_0_45;
	wire [WIDTH*2-1+3:0] tmp03_0_46;
	wire [WIDTH*2-1+3:0] tmp03_0_47;
	wire [WIDTH*2-1+3:0] tmp03_0_48;
	wire [WIDTH*2-1+3:0] tmp03_0_49;
	wire [WIDTH*2-1+3:0] tmp03_0_50;
	wire [WIDTH*2-1+3:0] tmp03_0_51;
	wire [WIDTH*2-1+3:0] tmp03_0_52;
	wire [WIDTH*2-1+3:0] tmp03_0_53;
	wire [WIDTH*2-1+3:0] tmp03_0_54;
	wire [WIDTH*2-1+3:0] tmp03_0_55;
	wire [WIDTH*2-1+3:0] tmp03_0_56;
	wire [WIDTH*2-1+3:0] tmp03_0_57;
	wire [WIDTH*2-1+3:0] tmp03_0_58;
	wire [WIDTH*2-1+3:0] tmp03_0_59;
	wire [WIDTH*2-1+3:0] tmp03_0_60;
	wire [WIDTH*2-1+3:0] tmp03_0_61;
	wire [WIDTH*2-1+3:0] tmp03_0_62;
	wire [WIDTH*2-1+3:0] tmp03_0_63;
	wire [WIDTH*2-1+3:0] tmp03_0_64;
	wire [WIDTH*2-1+3:0] tmp03_0_65;
	wire [WIDTH*2-1+3:0] tmp03_0_66;
	wire [WIDTH*2-1+3:0] tmp03_0_67;
	wire [WIDTH*2-1+3:0] tmp03_0_68;
	wire [WIDTH*2-1+3:0] tmp03_0_69;
	wire [WIDTH*2-1+3:0] tmp03_0_70;
	wire [WIDTH*2-1+3:0] tmp03_0_71;
	wire [WIDTH*2-1+3:0] tmp03_0_72;
	wire [WIDTH*2-1+3:0] tmp03_0_73;
	wire [WIDTH*2-1+3:0] tmp03_0_74;
	wire [WIDTH*2-1+3:0] tmp03_0_75;
	wire [WIDTH*2-1+3:0] tmp03_0_76;
	wire [WIDTH*2-1+3:0] tmp03_0_77;
	wire [WIDTH*2-1+3:0] tmp03_0_78;
	wire [WIDTH*2-1+3:0] tmp03_0_79;
	wire [WIDTH*2-1+3:0] tmp03_0_80;
	wire [WIDTH*2-1+3:0] tmp03_0_81;
	wire [WIDTH*2-1+3:0] tmp03_0_82;
	wire [WIDTH*2-1+3:0] tmp03_0_83;
	wire [WIDTH*2-1+3:0] tmp03_1_0;
	wire [WIDTH*2-1+3:0] tmp03_1_1;
	wire [WIDTH*2-1+3:0] tmp03_1_2;
	wire [WIDTH*2-1+3:0] tmp03_1_3;
	wire [WIDTH*2-1+3:0] tmp03_1_4;
	wire [WIDTH*2-1+3:0] tmp03_1_5;
	wire [WIDTH*2-1+3:0] tmp03_1_6;
	wire [WIDTH*2-1+3:0] tmp03_1_7;
	wire [WIDTH*2-1+3:0] tmp03_1_8;
	wire [WIDTH*2-1+3:0] tmp03_1_9;
	wire [WIDTH*2-1+3:0] tmp03_1_10;
	wire [WIDTH*2-1+3:0] tmp03_1_11;
	wire [WIDTH*2-1+3:0] tmp03_1_12;
	wire [WIDTH*2-1+3:0] tmp03_1_13;
	wire [WIDTH*2-1+3:0] tmp03_1_14;
	wire [WIDTH*2-1+3:0] tmp03_1_15;
	wire [WIDTH*2-1+3:0] tmp03_1_16;
	wire [WIDTH*2-1+3:0] tmp03_1_17;
	wire [WIDTH*2-1+3:0] tmp03_1_18;
	wire [WIDTH*2-1+3:0] tmp03_1_19;
	wire [WIDTH*2-1+3:0] tmp03_1_20;
	wire [WIDTH*2-1+3:0] tmp03_1_21;
	wire [WIDTH*2-1+3:0] tmp03_1_22;
	wire [WIDTH*2-1+3:0] tmp03_1_23;
	wire [WIDTH*2-1+3:0] tmp03_1_24;
	wire [WIDTH*2-1+3:0] tmp03_1_25;
	wire [WIDTH*2-1+3:0] tmp03_1_26;
	wire [WIDTH*2-1+3:0] tmp03_1_27;
	wire [WIDTH*2-1+3:0] tmp03_1_28;
	wire [WIDTH*2-1+3:0] tmp03_1_29;
	wire [WIDTH*2-1+3:0] tmp03_1_30;
	wire [WIDTH*2-1+3:0] tmp03_1_31;
	wire [WIDTH*2-1+3:0] tmp03_1_32;
	wire [WIDTH*2-1+3:0] tmp03_1_33;
	wire [WIDTH*2-1+3:0] tmp03_1_34;
	wire [WIDTH*2-1+3:0] tmp03_1_35;
	wire [WIDTH*2-1+3:0] tmp03_1_36;
	wire [WIDTH*2-1+3:0] tmp03_1_37;
	wire [WIDTH*2-1+3:0] tmp03_1_38;
	wire [WIDTH*2-1+3:0] tmp03_1_39;
	wire [WIDTH*2-1+3:0] tmp03_1_40;
	wire [WIDTH*2-1+3:0] tmp03_1_41;
	wire [WIDTH*2-1+3:0] tmp03_1_42;
	wire [WIDTH*2-1+3:0] tmp03_1_43;
	wire [WIDTH*2-1+3:0] tmp03_1_44;
	wire [WIDTH*2-1+3:0] tmp03_1_45;
	wire [WIDTH*2-1+3:0] tmp03_1_46;
	wire [WIDTH*2-1+3:0] tmp03_1_47;
	wire [WIDTH*2-1+3:0] tmp03_1_48;
	wire [WIDTH*2-1+3:0] tmp03_1_49;
	wire [WIDTH*2-1+3:0] tmp03_1_50;
	wire [WIDTH*2-1+3:0] tmp03_1_51;
	wire [WIDTH*2-1+3:0] tmp03_1_52;
	wire [WIDTH*2-1+3:0] tmp03_1_53;
	wire [WIDTH*2-1+3:0] tmp03_1_54;
	wire [WIDTH*2-1+3:0] tmp03_1_55;
	wire [WIDTH*2-1+3:0] tmp03_1_56;
	wire [WIDTH*2-1+3:0] tmp03_1_57;
	wire [WIDTH*2-1+3:0] tmp03_1_58;
	wire [WIDTH*2-1+3:0] tmp03_1_59;
	wire [WIDTH*2-1+3:0] tmp03_1_60;
	wire [WIDTH*2-1+3:0] tmp03_1_61;
	wire [WIDTH*2-1+3:0] tmp03_1_62;
	wire [WIDTH*2-1+3:0] tmp03_1_63;
	wire [WIDTH*2-1+3:0] tmp03_1_64;
	wire [WIDTH*2-1+3:0] tmp03_1_65;
	wire [WIDTH*2-1+3:0] tmp03_1_66;
	wire [WIDTH*2-1+3:0] tmp03_1_67;
	wire [WIDTH*2-1+3:0] tmp03_1_68;
	wire [WIDTH*2-1+3:0] tmp03_1_69;
	wire [WIDTH*2-1+3:0] tmp03_1_70;
	wire [WIDTH*2-1+3:0] tmp03_1_71;
	wire [WIDTH*2-1+3:0] tmp03_1_72;
	wire [WIDTH*2-1+3:0] tmp03_1_73;
	wire [WIDTH*2-1+3:0] tmp03_1_74;
	wire [WIDTH*2-1+3:0] tmp03_1_75;
	wire [WIDTH*2-1+3:0] tmp03_1_76;
	wire [WIDTH*2-1+3:0] tmp03_1_77;
	wire [WIDTH*2-1+3:0] tmp03_1_78;
	wire [WIDTH*2-1+3:0] tmp03_1_79;
	wire [WIDTH*2-1+3:0] tmp03_1_80;
	wire [WIDTH*2-1+3:0] tmp03_1_81;
	wire [WIDTH*2-1+3:0] tmp03_1_82;
	wire [WIDTH*2-1+3:0] tmp03_1_83;
	wire [WIDTH*2-1+3:0] tmp03_2_0;
	wire [WIDTH*2-1+3:0] tmp03_2_1;
	wire [WIDTH*2-1+3:0] tmp03_2_2;
	wire [WIDTH*2-1+3:0] tmp03_2_3;
	wire [WIDTH*2-1+3:0] tmp03_2_4;
	wire [WIDTH*2-1+3:0] tmp03_2_5;
	wire [WIDTH*2-1+3:0] tmp03_2_6;
	wire [WIDTH*2-1+3:0] tmp03_2_7;
	wire [WIDTH*2-1+3:0] tmp03_2_8;
	wire [WIDTH*2-1+3:0] tmp03_2_9;
	wire [WIDTH*2-1+3:0] tmp03_2_10;
	wire [WIDTH*2-1+3:0] tmp03_2_11;
	wire [WIDTH*2-1+3:0] tmp03_2_12;
	wire [WIDTH*2-1+3:0] tmp03_2_13;
	wire [WIDTH*2-1+3:0] tmp03_2_14;
	wire [WIDTH*2-1+3:0] tmp03_2_15;
	wire [WIDTH*2-1+3:0] tmp03_2_16;
	wire [WIDTH*2-1+3:0] tmp03_2_17;
	wire [WIDTH*2-1+3:0] tmp03_2_18;
	wire [WIDTH*2-1+3:0] tmp03_2_19;
	wire [WIDTH*2-1+3:0] tmp03_2_20;
	wire [WIDTH*2-1+3:0] tmp03_2_21;
	wire [WIDTH*2-1+3:0] tmp03_2_22;
	wire [WIDTH*2-1+3:0] tmp03_2_23;
	wire [WIDTH*2-1+3:0] tmp03_2_24;
	wire [WIDTH*2-1+3:0] tmp03_2_25;
	wire [WIDTH*2-1+3:0] tmp03_2_26;
	wire [WIDTH*2-1+3:0] tmp03_2_27;
	wire [WIDTH*2-1+3:0] tmp03_2_28;
	wire [WIDTH*2-1+3:0] tmp03_2_29;
	wire [WIDTH*2-1+3:0] tmp03_2_30;
	wire [WIDTH*2-1+3:0] tmp03_2_31;
	wire [WIDTH*2-1+3:0] tmp03_2_32;
	wire [WIDTH*2-1+3:0] tmp03_2_33;
	wire [WIDTH*2-1+3:0] tmp03_2_34;
	wire [WIDTH*2-1+3:0] tmp03_2_35;
	wire [WIDTH*2-1+3:0] tmp03_2_36;
	wire [WIDTH*2-1+3:0] tmp03_2_37;
	wire [WIDTH*2-1+3:0] tmp03_2_38;
	wire [WIDTH*2-1+3:0] tmp03_2_39;
	wire [WIDTH*2-1+3:0] tmp03_2_40;
	wire [WIDTH*2-1+3:0] tmp03_2_41;
	wire [WIDTH*2-1+3:0] tmp03_2_42;
	wire [WIDTH*2-1+3:0] tmp03_2_43;
	wire [WIDTH*2-1+3:0] tmp03_2_44;
	wire [WIDTH*2-1+3:0] tmp03_2_45;
	wire [WIDTH*2-1+3:0] tmp03_2_46;
	wire [WIDTH*2-1+3:0] tmp03_2_47;
	wire [WIDTH*2-1+3:0] tmp03_2_48;
	wire [WIDTH*2-1+3:0] tmp03_2_49;
	wire [WIDTH*2-1+3:0] tmp03_2_50;
	wire [WIDTH*2-1+3:0] tmp03_2_51;
	wire [WIDTH*2-1+3:0] tmp03_2_52;
	wire [WIDTH*2-1+3:0] tmp03_2_53;
	wire [WIDTH*2-1+3:0] tmp03_2_54;
	wire [WIDTH*2-1+3:0] tmp03_2_55;
	wire [WIDTH*2-1+3:0] tmp03_2_56;
	wire [WIDTH*2-1+3:0] tmp03_2_57;
	wire [WIDTH*2-1+3:0] tmp03_2_58;
	wire [WIDTH*2-1+3:0] tmp03_2_59;
	wire [WIDTH*2-1+3:0] tmp03_2_60;
	wire [WIDTH*2-1+3:0] tmp03_2_61;
	wire [WIDTH*2-1+3:0] tmp03_2_62;
	wire [WIDTH*2-1+3:0] tmp03_2_63;
	wire [WIDTH*2-1+3:0] tmp03_2_64;
	wire [WIDTH*2-1+3:0] tmp03_2_65;
	wire [WIDTH*2-1+3:0] tmp03_2_66;
	wire [WIDTH*2-1+3:0] tmp03_2_67;
	wire [WIDTH*2-1+3:0] tmp03_2_68;
	wire [WIDTH*2-1+3:0] tmp03_2_69;
	wire [WIDTH*2-1+3:0] tmp03_2_70;
	wire [WIDTH*2-1+3:0] tmp03_2_71;
	wire [WIDTH*2-1+3:0] tmp03_2_72;
	wire [WIDTH*2-1+3:0] tmp03_2_73;
	wire [WIDTH*2-1+3:0] tmp03_2_74;
	wire [WIDTH*2-1+3:0] tmp03_2_75;
	wire [WIDTH*2-1+3:0] tmp03_2_76;
	wire [WIDTH*2-1+3:0] tmp03_2_77;
	wire [WIDTH*2-1+3:0] tmp03_2_78;
	wire [WIDTH*2-1+3:0] tmp03_2_79;
	wire [WIDTH*2-1+3:0] tmp03_2_80;
	wire [WIDTH*2-1+3:0] tmp03_2_81;
	wire [WIDTH*2-1+3:0] tmp03_2_82;
	wire [WIDTH*2-1+3:0] tmp03_2_83;
	wire [WIDTH*2-1+3:0] tmp03_3_0;
	wire [WIDTH*2-1+3:0] tmp03_3_1;
	wire [WIDTH*2-1+3:0] tmp03_3_2;
	wire [WIDTH*2-1+3:0] tmp03_3_3;
	wire [WIDTH*2-1+3:0] tmp03_3_4;
	wire [WIDTH*2-1+3:0] tmp03_3_5;
	wire [WIDTH*2-1+3:0] tmp03_3_6;
	wire [WIDTH*2-1+3:0] tmp03_3_7;
	wire [WIDTH*2-1+3:0] tmp03_3_8;
	wire [WIDTH*2-1+3:0] tmp03_3_9;
	wire [WIDTH*2-1+3:0] tmp03_3_10;
	wire [WIDTH*2-1+3:0] tmp03_3_11;
	wire [WIDTH*2-1+3:0] tmp03_3_12;
	wire [WIDTH*2-1+3:0] tmp03_3_13;
	wire [WIDTH*2-1+3:0] tmp03_3_14;
	wire [WIDTH*2-1+3:0] tmp03_3_15;
	wire [WIDTH*2-1+3:0] tmp03_3_16;
	wire [WIDTH*2-1+3:0] tmp03_3_17;
	wire [WIDTH*2-1+3:0] tmp03_3_18;
	wire [WIDTH*2-1+3:0] tmp03_3_19;
	wire [WIDTH*2-1+3:0] tmp03_3_20;
	wire [WIDTH*2-1+3:0] tmp03_3_21;
	wire [WIDTH*2-1+3:0] tmp03_3_22;
	wire [WIDTH*2-1+3:0] tmp03_3_23;
	wire [WIDTH*2-1+3:0] tmp03_3_24;
	wire [WIDTH*2-1+3:0] tmp03_3_25;
	wire [WIDTH*2-1+3:0] tmp03_3_26;
	wire [WIDTH*2-1+3:0] tmp03_3_27;
	wire [WIDTH*2-1+3:0] tmp03_3_28;
	wire [WIDTH*2-1+3:0] tmp03_3_29;
	wire [WIDTH*2-1+3:0] tmp03_3_30;
	wire [WIDTH*2-1+3:0] tmp03_3_31;
	wire [WIDTH*2-1+3:0] tmp03_3_32;
	wire [WIDTH*2-1+3:0] tmp03_3_33;
	wire [WIDTH*2-1+3:0] tmp03_3_34;
	wire [WIDTH*2-1+3:0] tmp03_3_35;
	wire [WIDTH*2-1+3:0] tmp03_3_36;
	wire [WIDTH*2-1+3:0] tmp03_3_37;
	wire [WIDTH*2-1+3:0] tmp03_3_38;
	wire [WIDTH*2-1+3:0] tmp03_3_39;
	wire [WIDTH*2-1+3:0] tmp03_3_40;
	wire [WIDTH*2-1+3:0] tmp03_3_41;
	wire [WIDTH*2-1+3:0] tmp03_3_42;
	wire [WIDTH*2-1+3:0] tmp03_3_43;
	wire [WIDTH*2-1+3:0] tmp03_3_44;
	wire [WIDTH*2-1+3:0] tmp03_3_45;
	wire [WIDTH*2-1+3:0] tmp03_3_46;
	wire [WIDTH*2-1+3:0] tmp03_3_47;
	wire [WIDTH*2-1+3:0] tmp03_3_48;
	wire [WIDTH*2-1+3:0] tmp03_3_49;
	wire [WIDTH*2-1+3:0] tmp03_3_50;
	wire [WIDTH*2-1+3:0] tmp03_3_51;
	wire [WIDTH*2-1+3:0] tmp03_3_52;
	wire [WIDTH*2-1+3:0] tmp03_3_53;
	wire [WIDTH*2-1+3:0] tmp03_3_54;
	wire [WIDTH*2-1+3:0] tmp03_3_55;
	wire [WIDTH*2-1+3:0] tmp03_3_56;
	wire [WIDTH*2-1+3:0] tmp03_3_57;
	wire [WIDTH*2-1+3:0] tmp03_3_58;
	wire [WIDTH*2-1+3:0] tmp03_3_59;
	wire [WIDTH*2-1+3:0] tmp03_3_60;
	wire [WIDTH*2-1+3:0] tmp03_3_61;
	wire [WIDTH*2-1+3:0] tmp03_3_62;
	wire [WIDTH*2-1+3:0] tmp03_3_63;
	wire [WIDTH*2-1+3:0] tmp03_3_64;
	wire [WIDTH*2-1+3:0] tmp03_3_65;
	wire [WIDTH*2-1+3:0] tmp03_3_66;
	wire [WIDTH*2-1+3:0] tmp03_3_67;
	wire [WIDTH*2-1+3:0] tmp03_3_68;
	wire [WIDTH*2-1+3:0] tmp03_3_69;
	wire [WIDTH*2-1+3:0] tmp03_3_70;
	wire [WIDTH*2-1+3:0] tmp03_3_71;
	wire [WIDTH*2-1+3:0] tmp03_3_72;
	wire [WIDTH*2-1+3:0] tmp03_3_73;
	wire [WIDTH*2-1+3:0] tmp03_3_74;
	wire [WIDTH*2-1+3:0] tmp03_3_75;
	wire [WIDTH*2-1+3:0] tmp03_3_76;
	wire [WIDTH*2-1+3:0] tmp03_3_77;
	wire [WIDTH*2-1+3:0] tmp03_3_78;
	wire [WIDTH*2-1+3:0] tmp03_3_79;
	wire [WIDTH*2-1+3:0] tmp03_3_80;
	wire [WIDTH*2-1+3:0] tmp03_3_81;
	wire [WIDTH*2-1+3:0] tmp03_3_82;
	wire [WIDTH*2-1+3:0] tmp03_3_83;
	wire [WIDTH*2-1+3:0] tmp03_4_0;
	wire [WIDTH*2-1+3:0] tmp03_4_1;
	wire [WIDTH*2-1+3:0] tmp03_4_2;
	wire [WIDTH*2-1+3:0] tmp03_4_3;
	wire [WIDTH*2-1+3:0] tmp03_4_4;
	wire [WIDTH*2-1+3:0] tmp03_4_5;
	wire [WIDTH*2-1+3:0] tmp03_4_6;
	wire [WIDTH*2-1+3:0] tmp03_4_7;
	wire [WIDTH*2-1+3:0] tmp03_4_8;
	wire [WIDTH*2-1+3:0] tmp03_4_9;
	wire [WIDTH*2-1+3:0] tmp03_4_10;
	wire [WIDTH*2-1+3:0] tmp03_4_11;
	wire [WIDTH*2-1+3:0] tmp03_4_12;
	wire [WIDTH*2-1+3:0] tmp03_4_13;
	wire [WIDTH*2-1+3:0] tmp03_4_14;
	wire [WIDTH*2-1+3:0] tmp03_4_15;
	wire [WIDTH*2-1+3:0] tmp03_4_16;
	wire [WIDTH*2-1+3:0] tmp03_4_17;
	wire [WIDTH*2-1+3:0] tmp03_4_18;
	wire [WIDTH*2-1+3:0] tmp03_4_19;
	wire [WIDTH*2-1+3:0] tmp03_4_20;
	wire [WIDTH*2-1+3:0] tmp03_4_21;
	wire [WIDTH*2-1+3:0] tmp03_4_22;
	wire [WIDTH*2-1+3:0] tmp03_4_23;
	wire [WIDTH*2-1+3:0] tmp03_4_24;
	wire [WIDTH*2-1+3:0] tmp03_4_25;
	wire [WIDTH*2-1+3:0] tmp03_4_26;
	wire [WIDTH*2-1+3:0] tmp03_4_27;
	wire [WIDTH*2-1+3:0] tmp03_4_28;
	wire [WIDTH*2-1+3:0] tmp03_4_29;
	wire [WIDTH*2-1+3:0] tmp03_4_30;
	wire [WIDTH*2-1+3:0] tmp03_4_31;
	wire [WIDTH*2-1+3:0] tmp03_4_32;
	wire [WIDTH*2-1+3:0] tmp03_4_33;
	wire [WIDTH*2-1+3:0] tmp03_4_34;
	wire [WIDTH*2-1+3:0] tmp03_4_35;
	wire [WIDTH*2-1+3:0] tmp03_4_36;
	wire [WIDTH*2-1+3:0] tmp03_4_37;
	wire [WIDTH*2-1+3:0] tmp03_4_38;
	wire [WIDTH*2-1+3:0] tmp03_4_39;
	wire [WIDTH*2-1+3:0] tmp03_4_40;
	wire [WIDTH*2-1+3:0] tmp03_4_41;
	wire [WIDTH*2-1+3:0] tmp03_4_42;
	wire [WIDTH*2-1+3:0] tmp03_4_43;
	wire [WIDTH*2-1+3:0] tmp03_4_44;
	wire [WIDTH*2-1+3:0] tmp03_4_45;
	wire [WIDTH*2-1+3:0] tmp03_4_46;
	wire [WIDTH*2-1+3:0] tmp03_4_47;
	wire [WIDTH*2-1+3:0] tmp03_4_48;
	wire [WIDTH*2-1+3:0] tmp03_4_49;
	wire [WIDTH*2-1+3:0] tmp03_4_50;
	wire [WIDTH*2-1+3:0] tmp03_4_51;
	wire [WIDTH*2-1+3:0] tmp03_4_52;
	wire [WIDTH*2-1+3:0] tmp03_4_53;
	wire [WIDTH*2-1+3:0] tmp03_4_54;
	wire [WIDTH*2-1+3:0] tmp03_4_55;
	wire [WIDTH*2-1+3:0] tmp03_4_56;
	wire [WIDTH*2-1+3:0] tmp03_4_57;
	wire [WIDTH*2-1+3:0] tmp03_4_58;
	wire [WIDTH*2-1+3:0] tmp03_4_59;
	wire [WIDTH*2-1+3:0] tmp03_4_60;
	wire [WIDTH*2-1+3:0] tmp03_4_61;
	wire [WIDTH*2-1+3:0] tmp03_4_62;
	wire [WIDTH*2-1+3:0] tmp03_4_63;
	wire [WIDTH*2-1+3:0] tmp03_4_64;
	wire [WIDTH*2-1+3:0] tmp03_4_65;
	wire [WIDTH*2-1+3:0] tmp03_4_66;
	wire [WIDTH*2-1+3:0] tmp03_4_67;
	wire [WIDTH*2-1+3:0] tmp03_4_68;
	wire [WIDTH*2-1+3:0] tmp03_4_69;
	wire [WIDTH*2-1+3:0] tmp03_4_70;
	wire [WIDTH*2-1+3:0] tmp03_4_71;
	wire [WIDTH*2-1+3:0] tmp03_4_72;
	wire [WIDTH*2-1+3:0] tmp03_4_73;
	wire [WIDTH*2-1+3:0] tmp03_4_74;
	wire [WIDTH*2-1+3:0] tmp03_4_75;
	wire [WIDTH*2-1+3:0] tmp03_4_76;
	wire [WIDTH*2-1+3:0] tmp03_4_77;
	wire [WIDTH*2-1+3:0] tmp03_4_78;
	wire [WIDTH*2-1+3:0] tmp03_4_79;
	wire [WIDTH*2-1+3:0] tmp03_4_80;
	wire [WIDTH*2-1+3:0] tmp03_4_81;
	wire [WIDTH*2-1+3:0] tmp03_4_82;
	wire [WIDTH*2-1+3:0] tmp03_4_83;
	wire [WIDTH*2-1+3:0] tmp03_5_0;
	wire [WIDTH*2-1+3:0] tmp03_5_1;
	wire [WIDTH*2-1+3:0] tmp03_5_2;
	wire [WIDTH*2-1+3:0] tmp03_5_3;
	wire [WIDTH*2-1+3:0] tmp03_5_4;
	wire [WIDTH*2-1+3:0] tmp03_5_5;
	wire [WIDTH*2-1+3:0] tmp03_5_6;
	wire [WIDTH*2-1+3:0] tmp03_5_7;
	wire [WIDTH*2-1+3:0] tmp03_5_8;
	wire [WIDTH*2-1+3:0] tmp03_5_9;
	wire [WIDTH*2-1+3:0] tmp03_5_10;
	wire [WIDTH*2-1+3:0] tmp03_5_11;
	wire [WIDTH*2-1+3:0] tmp03_5_12;
	wire [WIDTH*2-1+3:0] tmp03_5_13;
	wire [WIDTH*2-1+3:0] tmp03_5_14;
	wire [WIDTH*2-1+3:0] tmp03_5_15;
	wire [WIDTH*2-1+3:0] tmp03_5_16;
	wire [WIDTH*2-1+3:0] tmp03_5_17;
	wire [WIDTH*2-1+3:0] tmp03_5_18;
	wire [WIDTH*2-1+3:0] tmp03_5_19;
	wire [WIDTH*2-1+3:0] tmp03_5_20;
	wire [WIDTH*2-1+3:0] tmp03_5_21;
	wire [WIDTH*2-1+3:0] tmp03_5_22;
	wire [WIDTH*2-1+3:0] tmp03_5_23;
	wire [WIDTH*2-1+3:0] tmp03_5_24;
	wire [WIDTH*2-1+3:0] tmp03_5_25;
	wire [WIDTH*2-1+3:0] tmp03_5_26;
	wire [WIDTH*2-1+3:0] tmp03_5_27;
	wire [WIDTH*2-1+3:0] tmp03_5_28;
	wire [WIDTH*2-1+3:0] tmp03_5_29;
	wire [WIDTH*2-1+3:0] tmp03_5_30;
	wire [WIDTH*2-1+3:0] tmp03_5_31;
	wire [WIDTH*2-1+3:0] tmp03_5_32;
	wire [WIDTH*2-1+3:0] tmp03_5_33;
	wire [WIDTH*2-1+3:0] tmp03_5_34;
	wire [WIDTH*2-1+3:0] tmp03_5_35;
	wire [WIDTH*2-1+3:0] tmp03_5_36;
	wire [WIDTH*2-1+3:0] tmp03_5_37;
	wire [WIDTH*2-1+3:0] tmp03_5_38;
	wire [WIDTH*2-1+3:0] tmp03_5_39;
	wire [WIDTH*2-1+3:0] tmp03_5_40;
	wire [WIDTH*2-1+3:0] tmp03_5_41;
	wire [WIDTH*2-1+3:0] tmp03_5_42;
	wire [WIDTH*2-1+3:0] tmp03_5_43;
	wire [WIDTH*2-1+3:0] tmp03_5_44;
	wire [WIDTH*2-1+3:0] tmp03_5_45;
	wire [WIDTH*2-1+3:0] tmp03_5_46;
	wire [WIDTH*2-1+3:0] tmp03_5_47;
	wire [WIDTH*2-1+3:0] tmp03_5_48;
	wire [WIDTH*2-1+3:0] tmp03_5_49;
	wire [WIDTH*2-1+3:0] tmp03_5_50;
	wire [WIDTH*2-1+3:0] tmp03_5_51;
	wire [WIDTH*2-1+3:0] tmp03_5_52;
	wire [WIDTH*2-1+3:0] tmp03_5_53;
	wire [WIDTH*2-1+3:0] tmp03_5_54;
	wire [WIDTH*2-1+3:0] tmp03_5_55;
	wire [WIDTH*2-1+3:0] tmp03_5_56;
	wire [WIDTH*2-1+3:0] tmp03_5_57;
	wire [WIDTH*2-1+3:0] tmp03_5_58;
	wire [WIDTH*2-1+3:0] tmp03_5_59;
	wire [WIDTH*2-1+3:0] tmp03_5_60;
	wire [WIDTH*2-1+3:0] tmp03_5_61;
	wire [WIDTH*2-1+3:0] tmp03_5_62;
	wire [WIDTH*2-1+3:0] tmp03_5_63;
	wire [WIDTH*2-1+3:0] tmp03_5_64;
	wire [WIDTH*2-1+3:0] tmp03_5_65;
	wire [WIDTH*2-1+3:0] tmp03_5_66;
	wire [WIDTH*2-1+3:0] tmp03_5_67;
	wire [WIDTH*2-1+3:0] tmp03_5_68;
	wire [WIDTH*2-1+3:0] tmp03_5_69;
	wire [WIDTH*2-1+3:0] tmp03_5_70;
	wire [WIDTH*2-1+3:0] tmp03_5_71;
	wire [WIDTH*2-1+3:0] tmp03_5_72;
	wire [WIDTH*2-1+3:0] tmp03_5_73;
	wire [WIDTH*2-1+3:0] tmp03_5_74;
	wire [WIDTH*2-1+3:0] tmp03_5_75;
	wire [WIDTH*2-1+3:0] tmp03_5_76;
	wire [WIDTH*2-1+3:0] tmp03_5_77;
	wire [WIDTH*2-1+3:0] tmp03_5_78;
	wire [WIDTH*2-1+3:0] tmp03_5_79;
	wire [WIDTH*2-1+3:0] tmp03_5_80;
	wire [WIDTH*2-1+3:0] tmp03_5_81;
	wire [WIDTH*2-1+3:0] tmp03_5_82;
	wire [WIDTH*2-1+3:0] tmp03_5_83;
	wire [WIDTH*2-1+3:0] tmp03_6_0;
	wire [WIDTH*2-1+3:0] tmp03_6_1;
	wire [WIDTH*2-1+3:0] tmp03_6_2;
	wire [WIDTH*2-1+3:0] tmp03_6_3;
	wire [WIDTH*2-1+3:0] tmp03_6_4;
	wire [WIDTH*2-1+3:0] tmp03_6_5;
	wire [WIDTH*2-1+3:0] tmp03_6_6;
	wire [WIDTH*2-1+3:0] tmp03_6_7;
	wire [WIDTH*2-1+3:0] tmp03_6_8;
	wire [WIDTH*2-1+3:0] tmp03_6_9;
	wire [WIDTH*2-1+3:0] tmp03_6_10;
	wire [WIDTH*2-1+3:0] tmp03_6_11;
	wire [WIDTH*2-1+3:0] tmp03_6_12;
	wire [WIDTH*2-1+3:0] tmp03_6_13;
	wire [WIDTH*2-1+3:0] tmp03_6_14;
	wire [WIDTH*2-1+3:0] tmp03_6_15;
	wire [WIDTH*2-1+3:0] tmp03_6_16;
	wire [WIDTH*2-1+3:0] tmp03_6_17;
	wire [WIDTH*2-1+3:0] tmp03_6_18;
	wire [WIDTH*2-1+3:0] tmp03_6_19;
	wire [WIDTH*2-1+3:0] tmp03_6_20;
	wire [WIDTH*2-1+3:0] tmp03_6_21;
	wire [WIDTH*2-1+3:0] tmp03_6_22;
	wire [WIDTH*2-1+3:0] tmp03_6_23;
	wire [WIDTH*2-1+3:0] tmp03_6_24;
	wire [WIDTH*2-1+3:0] tmp03_6_25;
	wire [WIDTH*2-1+3:0] tmp03_6_26;
	wire [WIDTH*2-1+3:0] tmp03_6_27;
	wire [WIDTH*2-1+3:0] tmp03_6_28;
	wire [WIDTH*2-1+3:0] tmp03_6_29;
	wire [WIDTH*2-1+3:0] tmp03_6_30;
	wire [WIDTH*2-1+3:0] tmp03_6_31;
	wire [WIDTH*2-1+3:0] tmp03_6_32;
	wire [WIDTH*2-1+3:0] tmp03_6_33;
	wire [WIDTH*2-1+3:0] tmp03_6_34;
	wire [WIDTH*2-1+3:0] tmp03_6_35;
	wire [WIDTH*2-1+3:0] tmp03_6_36;
	wire [WIDTH*2-1+3:0] tmp03_6_37;
	wire [WIDTH*2-1+3:0] tmp03_6_38;
	wire [WIDTH*2-1+3:0] tmp03_6_39;
	wire [WIDTH*2-1+3:0] tmp03_6_40;
	wire [WIDTH*2-1+3:0] tmp03_6_41;
	wire [WIDTH*2-1+3:0] tmp03_6_42;
	wire [WIDTH*2-1+3:0] tmp03_6_43;
	wire [WIDTH*2-1+3:0] tmp03_6_44;
	wire [WIDTH*2-1+3:0] tmp03_6_45;
	wire [WIDTH*2-1+3:0] tmp03_6_46;
	wire [WIDTH*2-1+3:0] tmp03_6_47;
	wire [WIDTH*2-1+3:0] tmp03_6_48;
	wire [WIDTH*2-1+3:0] tmp03_6_49;
	wire [WIDTH*2-1+3:0] tmp03_6_50;
	wire [WIDTH*2-1+3:0] tmp03_6_51;
	wire [WIDTH*2-1+3:0] tmp03_6_52;
	wire [WIDTH*2-1+3:0] tmp03_6_53;
	wire [WIDTH*2-1+3:0] tmp03_6_54;
	wire [WIDTH*2-1+3:0] tmp03_6_55;
	wire [WIDTH*2-1+3:0] tmp03_6_56;
	wire [WIDTH*2-1+3:0] tmp03_6_57;
	wire [WIDTH*2-1+3:0] tmp03_6_58;
	wire [WIDTH*2-1+3:0] tmp03_6_59;
	wire [WIDTH*2-1+3:0] tmp03_6_60;
	wire [WIDTH*2-1+3:0] tmp03_6_61;
	wire [WIDTH*2-1+3:0] tmp03_6_62;
	wire [WIDTH*2-1+3:0] tmp03_6_63;
	wire [WIDTH*2-1+3:0] tmp03_6_64;
	wire [WIDTH*2-1+3:0] tmp03_6_65;
	wire [WIDTH*2-1+3:0] tmp03_6_66;
	wire [WIDTH*2-1+3:0] tmp03_6_67;
	wire [WIDTH*2-1+3:0] tmp03_6_68;
	wire [WIDTH*2-1+3:0] tmp03_6_69;
	wire [WIDTH*2-1+3:0] tmp03_6_70;
	wire [WIDTH*2-1+3:0] tmp03_6_71;
	wire [WIDTH*2-1+3:0] tmp03_6_72;
	wire [WIDTH*2-1+3:0] tmp03_6_73;
	wire [WIDTH*2-1+3:0] tmp03_6_74;
	wire [WIDTH*2-1+3:0] tmp03_6_75;
	wire [WIDTH*2-1+3:0] tmp03_6_76;
	wire [WIDTH*2-1+3:0] tmp03_6_77;
	wire [WIDTH*2-1+3:0] tmp03_6_78;
	wire [WIDTH*2-1+3:0] tmp03_6_79;
	wire [WIDTH*2-1+3:0] tmp03_6_80;
	wire [WIDTH*2-1+3:0] tmp03_6_81;
	wire [WIDTH*2-1+3:0] tmp03_6_82;
	wire [WIDTH*2-1+3:0] tmp03_6_83;
	wire [WIDTH*2-1+3:0] tmp03_7_0;
	wire [WIDTH*2-1+3:0] tmp03_7_1;
	wire [WIDTH*2-1+3:0] tmp03_7_2;
	wire [WIDTH*2-1+3:0] tmp03_7_3;
	wire [WIDTH*2-1+3:0] tmp03_7_4;
	wire [WIDTH*2-1+3:0] tmp03_7_5;
	wire [WIDTH*2-1+3:0] tmp03_7_6;
	wire [WIDTH*2-1+3:0] tmp03_7_7;
	wire [WIDTH*2-1+3:0] tmp03_7_8;
	wire [WIDTH*2-1+3:0] tmp03_7_9;
	wire [WIDTH*2-1+3:0] tmp03_7_10;
	wire [WIDTH*2-1+3:0] tmp03_7_11;
	wire [WIDTH*2-1+3:0] tmp03_7_12;
	wire [WIDTH*2-1+3:0] tmp03_7_13;
	wire [WIDTH*2-1+3:0] tmp03_7_14;
	wire [WIDTH*2-1+3:0] tmp03_7_15;
	wire [WIDTH*2-1+3:0] tmp03_7_16;
	wire [WIDTH*2-1+3:0] tmp03_7_17;
	wire [WIDTH*2-1+3:0] tmp03_7_18;
	wire [WIDTH*2-1+3:0] tmp03_7_19;
	wire [WIDTH*2-1+3:0] tmp03_7_20;
	wire [WIDTH*2-1+3:0] tmp03_7_21;
	wire [WIDTH*2-1+3:0] tmp03_7_22;
	wire [WIDTH*2-1+3:0] tmp03_7_23;
	wire [WIDTH*2-1+3:0] tmp03_7_24;
	wire [WIDTH*2-1+3:0] tmp03_7_25;
	wire [WIDTH*2-1+3:0] tmp03_7_26;
	wire [WIDTH*2-1+3:0] tmp03_7_27;
	wire [WIDTH*2-1+3:0] tmp03_7_28;
	wire [WIDTH*2-1+3:0] tmp03_7_29;
	wire [WIDTH*2-1+3:0] tmp03_7_30;
	wire [WIDTH*2-1+3:0] tmp03_7_31;
	wire [WIDTH*2-1+3:0] tmp03_7_32;
	wire [WIDTH*2-1+3:0] tmp03_7_33;
	wire [WIDTH*2-1+3:0] tmp03_7_34;
	wire [WIDTH*2-1+3:0] tmp03_7_35;
	wire [WIDTH*2-1+3:0] tmp03_7_36;
	wire [WIDTH*2-1+3:0] tmp03_7_37;
	wire [WIDTH*2-1+3:0] tmp03_7_38;
	wire [WIDTH*2-1+3:0] tmp03_7_39;
	wire [WIDTH*2-1+3:0] tmp03_7_40;
	wire [WIDTH*2-1+3:0] tmp03_7_41;
	wire [WIDTH*2-1+3:0] tmp03_7_42;
	wire [WIDTH*2-1+3:0] tmp03_7_43;
	wire [WIDTH*2-1+3:0] tmp03_7_44;
	wire [WIDTH*2-1+3:0] tmp03_7_45;
	wire [WIDTH*2-1+3:0] tmp03_7_46;
	wire [WIDTH*2-1+3:0] tmp03_7_47;
	wire [WIDTH*2-1+3:0] tmp03_7_48;
	wire [WIDTH*2-1+3:0] tmp03_7_49;
	wire [WIDTH*2-1+3:0] tmp03_7_50;
	wire [WIDTH*2-1+3:0] tmp03_7_51;
	wire [WIDTH*2-1+3:0] tmp03_7_52;
	wire [WIDTH*2-1+3:0] tmp03_7_53;
	wire [WIDTH*2-1+3:0] tmp03_7_54;
	wire [WIDTH*2-1+3:0] tmp03_7_55;
	wire [WIDTH*2-1+3:0] tmp03_7_56;
	wire [WIDTH*2-1+3:0] tmp03_7_57;
	wire [WIDTH*2-1+3:0] tmp03_7_58;
	wire [WIDTH*2-1+3:0] tmp03_7_59;
	wire [WIDTH*2-1+3:0] tmp03_7_60;
	wire [WIDTH*2-1+3:0] tmp03_7_61;
	wire [WIDTH*2-1+3:0] tmp03_7_62;
	wire [WIDTH*2-1+3:0] tmp03_7_63;
	wire [WIDTH*2-1+3:0] tmp03_7_64;
	wire [WIDTH*2-1+3:0] tmp03_7_65;
	wire [WIDTH*2-1+3:0] tmp03_7_66;
	wire [WIDTH*2-1+3:0] tmp03_7_67;
	wire [WIDTH*2-1+3:0] tmp03_7_68;
	wire [WIDTH*2-1+3:0] tmp03_7_69;
	wire [WIDTH*2-1+3:0] tmp03_7_70;
	wire [WIDTH*2-1+3:0] tmp03_7_71;
	wire [WIDTH*2-1+3:0] tmp03_7_72;
	wire [WIDTH*2-1+3:0] tmp03_7_73;
	wire [WIDTH*2-1+3:0] tmp03_7_74;
	wire [WIDTH*2-1+3:0] tmp03_7_75;
	wire [WIDTH*2-1+3:0] tmp03_7_76;
	wire [WIDTH*2-1+3:0] tmp03_7_77;
	wire [WIDTH*2-1+3:0] tmp03_7_78;
	wire [WIDTH*2-1+3:0] tmp03_7_79;
	wire [WIDTH*2-1+3:0] tmp03_7_80;
	wire [WIDTH*2-1+3:0] tmp03_7_81;
	wire [WIDTH*2-1+3:0] tmp03_7_82;
	wire [WIDTH*2-1+3:0] tmp03_7_83;
	wire [WIDTH*2-1+3:0] tmp03_8_0;
	wire [WIDTH*2-1+3:0] tmp03_8_1;
	wire [WIDTH*2-1+3:0] tmp03_8_2;
	wire [WIDTH*2-1+3:0] tmp03_8_3;
	wire [WIDTH*2-1+3:0] tmp03_8_4;
	wire [WIDTH*2-1+3:0] tmp03_8_5;
	wire [WIDTH*2-1+3:0] tmp03_8_6;
	wire [WIDTH*2-1+3:0] tmp03_8_7;
	wire [WIDTH*2-1+3:0] tmp03_8_8;
	wire [WIDTH*2-1+3:0] tmp03_8_9;
	wire [WIDTH*2-1+3:0] tmp03_8_10;
	wire [WIDTH*2-1+3:0] tmp03_8_11;
	wire [WIDTH*2-1+3:0] tmp03_8_12;
	wire [WIDTH*2-1+3:0] tmp03_8_13;
	wire [WIDTH*2-1+3:0] tmp03_8_14;
	wire [WIDTH*2-1+3:0] tmp03_8_15;
	wire [WIDTH*2-1+3:0] tmp03_8_16;
	wire [WIDTH*2-1+3:0] tmp03_8_17;
	wire [WIDTH*2-1+3:0] tmp03_8_18;
	wire [WIDTH*2-1+3:0] tmp03_8_19;
	wire [WIDTH*2-1+3:0] tmp03_8_20;
	wire [WIDTH*2-1+3:0] tmp03_8_21;
	wire [WIDTH*2-1+3:0] tmp03_8_22;
	wire [WIDTH*2-1+3:0] tmp03_8_23;
	wire [WIDTH*2-1+3:0] tmp03_8_24;
	wire [WIDTH*2-1+3:0] tmp03_8_25;
	wire [WIDTH*2-1+3:0] tmp03_8_26;
	wire [WIDTH*2-1+3:0] tmp03_8_27;
	wire [WIDTH*2-1+3:0] tmp03_8_28;
	wire [WIDTH*2-1+3:0] tmp03_8_29;
	wire [WIDTH*2-1+3:0] tmp03_8_30;
	wire [WIDTH*2-1+3:0] tmp03_8_31;
	wire [WIDTH*2-1+3:0] tmp03_8_32;
	wire [WIDTH*2-1+3:0] tmp03_8_33;
	wire [WIDTH*2-1+3:0] tmp03_8_34;
	wire [WIDTH*2-1+3:0] tmp03_8_35;
	wire [WIDTH*2-1+3:0] tmp03_8_36;
	wire [WIDTH*2-1+3:0] tmp03_8_37;
	wire [WIDTH*2-1+3:0] tmp03_8_38;
	wire [WIDTH*2-1+3:0] tmp03_8_39;
	wire [WIDTH*2-1+3:0] tmp03_8_40;
	wire [WIDTH*2-1+3:0] tmp03_8_41;
	wire [WIDTH*2-1+3:0] tmp03_8_42;
	wire [WIDTH*2-1+3:0] tmp03_8_43;
	wire [WIDTH*2-1+3:0] tmp03_8_44;
	wire [WIDTH*2-1+3:0] tmp03_8_45;
	wire [WIDTH*2-1+3:0] tmp03_8_46;
	wire [WIDTH*2-1+3:0] tmp03_8_47;
	wire [WIDTH*2-1+3:0] tmp03_8_48;
	wire [WIDTH*2-1+3:0] tmp03_8_49;
	wire [WIDTH*2-1+3:0] tmp03_8_50;
	wire [WIDTH*2-1+3:0] tmp03_8_51;
	wire [WIDTH*2-1+3:0] tmp03_8_52;
	wire [WIDTH*2-1+3:0] tmp03_8_53;
	wire [WIDTH*2-1+3:0] tmp03_8_54;
	wire [WIDTH*2-1+3:0] tmp03_8_55;
	wire [WIDTH*2-1+3:0] tmp03_8_56;
	wire [WIDTH*2-1+3:0] tmp03_8_57;
	wire [WIDTH*2-1+3:0] tmp03_8_58;
	wire [WIDTH*2-1+3:0] tmp03_8_59;
	wire [WIDTH*2-1+3:0] tmp03_8_60;
	wire [WIDTH*2-1+3:0] tmp03_8_61;
	wire [WIDTH*2-1+3:0] tmp03_8_62;
	wire [WIDTH*2-1+3:0] tmp03_8_63;
	wire [WIDTH*2-1+3:0] tmp03_8_64;
	wire [WIDTH*2-1+3:0] tmp03_8_65;
	wire [WIDTH*2-1+3:0] tmp03_8_66;
	wire [WIDTH*2-1+3:0] tmp03_8_67;
	wire [WIDTH*2-1+3:0] tmp03_8_68;
	wire [WIDTH*2-1+3:0] tmp03_8_69;
	wire [WIDTH*2-1+3:0] tmp03_8_70;
	wire [WIDTH*2-1+3:0] tmp03_8_71;
	wire [WIDTH*2-1+3:0] tmp03_8_72;
	wire [WIDTH*2-1+3:0] tmp03_8_73;
	wire [WIDTH*2-1+3:0] tmp03_8_74;
	wire [WIDTH*2-1+3:0] tmp03_8_75;
	wire [WIDTH*2-1+3:0] tmp03_8_76;
	wire [WIDTH*2-1+3:0] tmp03_8_77;
	wire [WIDTH*2-1+3:0] tmp03_8_78;
	wire [WIDTH*2-1+3:0] tmp03_8_79;
	wire [WIDTH*2-1+3:0] tmp03_8_80;
	wire [WIDTH*2-1+3:0] tmp03_8_81;
	wire [WIDTH*2-1+3:0] tmp03_8_82;
	wire [WIDTH*2-1+3:0] tmp03_8_83;
	wire [WIDTH*2-1+3:0] tmp03_9_0;
	wire [WIDTH*2-1+3:0] tmp03_9_1;
	wire [WIDTH*2-1+3:0] tmp03_9_2;
	wire [WIDTH*2-1+3:0] tmp03_9_3;
	wire [WIDTH*2-1+3:0] tmp03_9_4;
	wire [WIDTH*2-1+3:0] tmp03_9_5;
	wire [WIDTH*2-1+3:0] tmp03_9_6;
	wire [WIDTH*2-1+3:0] tmp03_9_7;
	wire [WIDTH*2-1+3:0] tmp03_9_8;
	wire [WIDTH*2-1+3:0] tmp03_9_9;
	wire [WIDTH*2-1+3:0] tmp03_9_10;
	wire [WIDTH*2-1+3:0] tmp03_9_11;
	wire [WIDTH*2-1+3:0] tmp03_9_12;
	wire [WIDTH*2-1+3:0] tmp03_9_13;
	wire [WIDTH*2-1+3:0] tmp03_9_14;
	wire [WIDTH*2-1+3:0] tmp03_9_15;
	wire [WIDTH*2-1+3:0] tmp03_9_16;
	wire [WIDTH*2-1+3:0] tmp03_9_17;
	wire [WIDTH*2-1+3:0] tmp03_9_18;
	wire [WIDTH*2-1+3:0] tmp03_9_19;
	wire [WIDTH*2-1+3:0] tmp03_9_20;
	wire [WIDTH*2-1+3:0] tmp03_9_21;
	wire [WIDTH*2-1+3:0] tmp03_9_22;
	wire [WIDTH*2-1+3:0] tmp03_9_23;
	wire [WIDTH*2-1+3:0] tmp03_9_24;
	wire [WIDTH*2-1+3:0] tmp03_9_25;
	wire [WIDTH*2-1+3:0] tmp03_9_26;
	wire [WIDTH*2-1+3:0] tmp03_9_27;
	wire [WIDTH*2-1+3:0] tmp03_9_28;
	wire [WIDTH*2-1+3:0] tmp03_9_29;
	wire [WIDTH*2-1+3:0] tmp03_9_30;
	wire [WIDTH*2-1+3:0] tmp03_9_31;
	wire [WIDTH*2-1+3:0] tmp03_9_32;
	wire [WIDTH*2-1+3:0] tmp03_9_33;
	wire [WIDTH*2-1+3:0] tmp03_9_34;
	wire [WIDTH*2-1+3:0] tmp03_9_35;
	wire [WIDTH*2-1+3:0] tmp03_9_36;
	wire [WIDTH*2-1+3:0] tmp03_9_37;
	wire [WIDTH*2-1+3:0] tmp03_9_38;
	wire [WIDTH*2-1+3:0] tmp03_9_39;
	wire [WIDTH*2-1+3:0] tmp03_9_40;
	wire [WIDTH*2-1+3:0] tmp03_9_41;
	wire [WIDTH*2-1+3:0] tmp03_9_42;
	wire [WIDTH*2-1+3:0] tmp03_9_43;
	wire [WIDTH*2-1+3:0] tmp03_9_44;
	wire [WIDTH*2-1+3:0] tmp03_9_45;
	wire [WIDTH*2-1+3:0] tmp03_9_46;
	wire [WIDTH*2-1+3:0] tmp03_9_47;
	wire [WIDTH*2-1+3:0] tmp03_9_48;
	wire [WIDTH*2-1+3:0] tmp03_9_49;
	wire [WIDTH*2-1+3:0] tmp03_9_50;
	wire [WIDTH*2-1+3:0] tmp03_9_51;
	wire [WIDTH*2-1+3:0] tmp03_9_52;
	wire [WIDTH*2-1+3:0] tmp03_9_53;
	wire [WIDTH*2-1+3:0] tmp03_9_54;
	wire [WIDTH*2-1+3:0] tmp03_9_55;
	wire [WIDTH*2-1+3:0] tmp03_9_56;
	wire [WIDTH*2-1+3:0] tmp03_9_57;
	wire [WIDTH*2-1+3:0] tmp03_9_58;
	wire [WIDTH*2-1+3:0] tmp03_9_59;
	wire [WIDTH*2-1+3:0] tmp03_9_60;
	wire [WIDTH*2-1+3:0] tmp03_9_61;
	wire [WIDTH*2-1+3:0] tmp03_9_62;
	wire [WIDTH*2-1+3:0] tmp03_9_63;
	wire [WIDTH*2-1+3:0] tmp03_9_64;
	wire [WIDTH*2-1+3:0] tmp03_9_65;
	wire [WIDTH*2-1+3:0] tmp03_9_66;
	wire [WIDTH*2-1+3:0] tmp03_9_67;
	wire [WIDTH*2-1+3:0] tmp03_9_68;
	wire [WIDTH*2-1+3:0] tmp03_9_69;
	wire [WIDTH*2-1+3:0] tmp03_9_70;
	wire [WIDTH*2-1+3:0] tmp03_9_71;
	wire [WIDTH*2-1+3:0] tmp03_9_72;
	wire [WIDTH*2-1+3:0] tmp03_9_73;
	wire [WIDTH*2-1+3:0] tmp03_9_74;
	wire [WIDTH*2-1+3:0] tmp03_9_75;
	wire [WIDTH*2-1+3:0] tmp03_9_76;
	wire [WIDTH*2-1+3:0] tmp03_9_77;
	wire [WIDTH*2-1+3:0] tmp03_9_78;
	wire [WIDTH*2-1+3:0] tmp03_9_79;
	wire [WIDTH*2-1+3:0] tmp03_9_80;
	wire [WIDTH*2-1+3:0] tmp03_9_81;
	wire [WIDTH*2-1+3:0] tmp03_9_82;
	wire [WIDTH*2-1+3:0] tmp03_9_83;
	wire [WIDTH*2-1+3:0] tmp03_10_0;
	wire [WIDTH*2-1+3:0] tmp03_10_1;
	wire [WIDTH*2-1+3:0] tmp03_10_2;
	wire [WIDTH*2-1+3:0] tmp03_10_3;
	wire [WIDTH*2-1+3:0] tmp03_10_4;
	wire [WIDTH*2-1+3:0] tmp03_10_5;
	wire [WIDTH*2-1+3:0] tmp03_10_6;
	wire [WIDTH*2-1+3:0] tmp03_10_7;
	wire [WIDTH*2-1+3:0] tmp03_10_8;
	wire [WIDTH*2-1+3:0] tmp03_10_9;
	wire [WIDTH*2-1+3:0] tmp03_10_10;
	wire [WIDTH*2-1+3:0] tmp03_10_11;
	wire [WIDTH*2-1+3:0] tmp03_10_12;
	wire [WIDTH*2-1+3:0] tmp03_10_13;
	wire [WIDTH*2-1+3:0] tmp03_10_14;
	wire [WIDTH*2-1+3:0] tmp03_10_15;
	wire [WIDTH*2-1+3:0] tmp03_10_16;
	wire [WIDTH*2-1+3:0] tmp03_10_17;
	wire [WIDTH*2-1+3:0] tmp03_10_18;
	wire [WIDTH*2-1+3:0] tmp03_10_19;
	wire [WIDTH*2-1+3:0] tmp03_10_20;
	wire [WIDTH*2-1+3:0] tmp03_10_21;
	wire [WIDTH*2-1+3:0] tmp03_10_22;
	wire [WIDTH*2-1+3:0] tmp03_10_23;
	wire [WIDTH*2-1+3:0] tmp03_10_24;
	wire [WIDTH*2-1+3:0] tmp03_10_25;
	wire [WIDTH*2-1+3:0] tmp03_10_26;
	wire [WIDTH*2-1+3:0] tmp03_10_27;
	wire [WIDTH*2-1+3:0] tmp03_10_28;
	wire [WIDTH*2-1+3:0] tmp03_10_29;
	wire [WIDTH*2-1+3:0] tmp03_10_30;
	wire [WIDTH*2-1+3:0] tmp03_10_31;
	wire [WIDTH*2-1+3:0] tmp03_10_32;
	wire [WIDTH*2-1+3:0] tmp03_10_33;
	wire [WIDTH*2-1+3:0] tmp03_10_34;
	wire [WIDTH*2-1+3:0] tmp03_10_35;
	wire [WIDTH*2-1+3:0] tmp03_10_36;
	wire [WIDTH*2-1+3:0] tmp03_10_37;
	wire [WIDTH*2-1+3:0] tmp03_10_38;
	wire [WIDTH*2-1+3:0] tmp03_10_39;
	wire [WIDTH*2-1+3:0] tmp03_10_40;
	wire [WIDTH*2-1+3:0] tmp03_10_41;
	wire [WIDTH*2-1+3:0] tmp03_10_42;
	wire [WIDTH*2-1+3:0] tmp03_10_43;
	wire [WIDTH*2-1+3:0] tmp03_10_44;
	wire [WIDTH*2-1+3:0] tmp03_10_45;
	wire [WIDTH*2-1+3:0] tmp03_10_46;
	wire [WIDTH*2-1+3:0] tmp03_10_47;
	wire [WIDTH*2-1+3:0] tmp03_10_48;
	wire [WIDTH*2-1+3:0] tmp03_10_49;
	wire [WIDTH*2-1+3:0] tmp03_10_50;
	wire [WIDTH*2-1+3:0] tmp03_10_51;
	wire [WIDTH*2-1+3:0] tmp03_10_52;
	wire [WIDTH*2-1+3:0] tmp03_10_53;
	wire [WIDTH*2-1+3:0] tmp03_10_54;
	wire [WIDTH*2-1+3:0] tmp03_10_55;
	wire [WIDTH*2-1+3:0] tmp03_10_56;
	wire [WIDTH*2-1+3:0] tmp03_10_57;
	wire [WIDTH*2-1+3:0] tmp03_10_58;
	wire [WIDTH*2-1+3:0] tmp03_10_59;
	wire [WIDTH*2-1+3:0] tmp03_10_60;
	wire [WIDTH*2-1+3:0] tmp03_10_61;
	wire [WIDTH*2-1+3:0] tmp03_10_62;
	wire [WIDTH*2-1+3:0] tmp03_10_63;
	wire [WIDTH*2-1+3:0] tmp03_10_64;
	wire [WIDTH*2-1+3:0] tmp03_10_65;
	wire [WIDTH*2-1+3:0] tmp03_10_66;
	wire [WIDTH*2-1+3:0] tmp03_10_67;
	wire [WIDTH*2-1+3:0] tmp03_10_68;
	wire [WIDTH*2-1+3:0] tmp03_10_69;
	wire [WIDTH*2-1+3:0] tmp03_10_70;
	wire [WIDTH*2-1+3:0] tmp03_10_71;
	wire [WIDTH*2-1+3:0] tmp03_10_72;
	wire [WIDTH*2-1+3:0] tmp03_10_73;
	wire [WIDTH*2-1+3:0] tmp03_10_74;
	wire [WIDTH*2-1+3:0] tmp03_10_75;
	wire [WIDTH*2-1+3:0] tmp03_10_76;
	wire [WIDTH*2-1+3:0] tmp03_10_77;
	wire [WIDTH*2-1+3:0] tmp03_10_78;
	wire [WIDTH*2-1+3:0] tmp03_10_79;
	wire [WIDTH*2-1+3:0] tmp03_10_80;
	wire [WIDTH*2-1+3:0] tmp03_10_81;
	wire [WIDTH*2-1+3:0] tmp03_10_82;
	wire [WIDTH*2-1+3:0] tmp03_10_83;
	wire [WIDTH*2-1+3:0] tmp03_11_0;
	wire [WIDTH*2-1+3:0] tmp03_11_1;
	wire [WIDTH*2-1+3:0] tmp03_11_2;
	wire [WIDTH*2-1+3:0] tmp03_11_3;
	wire [WIDTH*2-1+3:0] tmp03_11_4;
	wire [WIDTH*2-1+3:0] tmp03_11_5;
	wire [WIDTH*2-1+3:0] tmp03_11_6;
	wire [WIDTH*2-1+3:0] tmp03_11_7;
	wire [WIDTH*2-1+3:0] tmp03_11_8;
	wire [WIDTH*2-1+3:0] tmp03_11_9;
	wire [WIDTH*2-1+3:0] tmp03_11_10;
	wire [WIDTH*2-1+3:0] tmp03_11_11;
	wire [WIDTH*2-1+3:0] tmp03_11_12;
	wire [WIDTH*2-1+3:0] tmp03_11_13;
	wire [WIDTH*2-1+3:0] tmp03_11_14;
	wire [WIDTH*2-1+3:0] tmp03_11_15;
	wire [WIDTH*2-1+3:0] tmp03_11_16;
	wire [WIDTH*2-1+3:0] tmp03_11_17;
	wire [WIDTH*2-1+3:0] tmp03_11_18;
	wire [WIDTH*2-1+3:0] tmp03_11_19;
	wire [WIDTH*2-1+3:0] tmp03_11_20;
	wire [WIDTH*2-1+3:0] tmp03_11_21;
	wire [WIDTH*2-1+3:0] tmp03_11_22;
	wire [WIDTH*2-1+3:0] tmp03_11_23;
	wire [WIDTH*2-1+3:0] tmp03_11_24;
	wire [WIDTH*2-1+3:0] tmp03_11_25;
	wire [WIDTH*2-1+3:0] tmp03_11_26;
	wire [WIDTH*2-1+3:0] tmp03_11_27;
	wire [WIDTH*2-1+3:0] tmp03_11_28;
	wire [WIDTH*2-1+3:0] tmp03_11_29;
	wire [WIDTH*2-1+3:0] tmp03_11_30;
	wire [WIDTH*2-1+3:0] tmp03_11_31;
	wire [WIDTH*2-1+3:0] tmp03_11_32;
	wire [WIDTH*2-1+3:0] tmp03_11_33;
	wire [WIDTH*2-1+3:0] tmp03_11_34;
	wire [WIDTH*2-1+3:0] tmp03_11_35;
	wire [WIDTH*2-1+3:0] tmp03_11_36;
	wire [WIDTH*2-1+3:0] tmp03_11_37;
	wire [WIDTH*2-1+3:0] tmp03_11_38;
	wire [WIDTH*2-1+3:0] tmp03_11_39;
	wire [WIDTH*2-1+3:0] tmp03_11_40;
	wire [WIDTH*2-1+3:0] tmp03_11_41;
	wire [WIDTH*2-1+3:0] tmp03_11_42;
	wire [WIDTH*2-1+3:0] tmp03_11_43;
	wire [WIDTH*2-1+3:0] tmp03_11_44;
	wire [WIDTH*2-1+3:0] tmp03_11_45;
	wire [WIDTH*2-1+3:0] tmp03_11_46;
	wire [WIDTH*2-1+3:0] tmp03_11_47;
	wire [WIDTH*2-1+3:0] tmp03_11_48;
	wire [WIDTH*2-1+3:0] tmp03_11_49;
	wire [WIDTH*2-1+3:0] tmp03_11_50;
	wire [WIDTH*2-1+3:0] tmp03_11_51;
	wire [WIDTH*2-1+3:0] tmp03_11_52;
	wire [WIDTH*2-1+3:0] tmp03_11_53;
	wire [WIDTH*2-1+3:0] tmp03_11_54;
	wire [WIDTH*2-1+3:0] tmp03_11_55;
	wire [WIDTH*2-1+3:0] tmp03_11_56;
	wire [WIDTH*2-1+3:0] tmp03_11_57;
	wire [WIDTH*2-1+3:0] tmp03_11_58;
	wire [WIDTH*2-1+3:0] tmp03_11_59;
	wire [WIDTH*2-1+3:0] tmp03_11_60;
	wire [WIDTH*2-1+3:0] tmp03_11_61;
	wire [WIDTH*2-1+3:0] tmp03_11_62;
	wire [WIDTH*2-1+3:0] tmp03_11_63;
	wire [WIDTH*2-1+3:0] tmp03_11_64;
	wire [WIDTH*2-1+3:0] tmp03_11_65;
	wire [WIDTH*2-1+3:0] tmp03_11_66;
	wire [WIDTH*2-1+3:0] tmp03_11_67;
	wire [WIDTH*2-1+3:0] tmp03_11_68;
	wire [WIDTH*2-1+3:0] tmp03_11_69;
	wire [WIDTH*2-1+3:0] tmp03_11_70;
	wire [WIDTH*2-1+3:0] tmp03_11_71;
	wire [WIDTH*2-1+3:0] tmp03_11_72;
	wire [WIDTH*2-1+3:0] tmp03_11_73;
	wire [WIDTH*2-1+3:0] tmp03_11_74;
	wire [WIDTH*2-1+3:0] tmp03_11_75;
	wire [WIDTH*2-1+3:0] tmp03_11_76;
	wire [WIDTH*2-1+3:0] tmp03_11_77;
	wire [WIDTH*2-1+3:0] tmp03_11_78;
	wire [WIDTH*2-1+3:0] tmp03_11_79;
	wire [WIDTH*2-1+3:0] tmp03_11_80;
	wire [WIDTH*2-1+3:0] tmp03_11_81;
	wire [WIDTH*2-1+3:0] tmp03_11_82;
	wire [WIDTH*2-1+3:0] tmp03_11_83;
	wire [WIDTH*2-1+3:0] tmp03_12_0;
	wire [WIDTH*2-1+3:0] tmp03_12_1;
	wire [WIDTH*2-1+3:0] tmp03_12_2;
	wire [WIDTH*2-1+3:0] tmp03_12_3;
	wire [WIDTH*2-1+3:0] tmp03_12_4;
	wire [WIDTH*2-1+3:0] tmp03_12_5;
	wire [WIDTH*2-1+3:0] tmp03_12_6;
	wire [WIDTH*2-1+3:0] tmp03_12_7;
	wire [WIDTH*2-1+3:0] tmp03_12_8;
	wire [WIDTH*2-1+3:0] tmp03_12_9;
	wire [WIDTH*2-1+3:0] tmp03_12_10;
	wire [WIDTH*2-1+3:0] tmp03_12_11;
	wire [WIDTH*2-1+3:0] tmp03_12_12;
	wire [WIDTH*2-1+3:0] tmp03_12_13;
	wire [WIDTH*2-1+3:0] tmp03_12_14;
	wire [WIDTH*2-1+3:0] tmp03_12_15;
	wire [WIDTH*2-1+3:0] tmp03_12_16;
	wire [WIDTH*2-1+3:0] tmp03_12_17;
	wire [WIDTH*2-1+3:0] tmp03_12_18;
	wire [WIDTH*2-1+3:0] tmp03_12_19;
	wire [WIDTH*2-1+3:0] tmp03_12_20;
	wire [WIDTH*2-1+3:0] tmp03_12_21;
	wire [WIDTH*2-1+3:0] tmp03_12_22;
	wire [WIDTH*2-1+3:0] tmp03_12_23;
	wire [WIDTH*2-1+3:0] tmp03_12_24;
	wire [WIDTH*2-1+3:0] tmp03_12_25;
	wire [WIDTH*2-1+3:0] tmp03_12_26;
	wire [WIDTH*2-1+3:0] tmp03_12_27;
	wire [WIDTH*2-1+3:0] tmp03_12_28;
	wire [WIDTH*2-1+3:0] tmp03_12_29;
	wire [WIDTH*2-1+3:0] tmp03_12_30;
	wire [WIDTH*2-1+3:0] tmp03_12_31;
	wire [WIDTH*2-1+3:0] tmp03_12_32;
	wire [WIDTH*2-1+3:0] tmp03_12_33;
	wire [WIDTH*2-1+3:0] tmp03_12_34;
	wire [WIDTH*2-1+3:0] tmp03_12_35;
	wire [WIDTH*2-1+3:0] tmp03_12_36;
	wire [WIDTH*2-1+3:0] tmp03_12_37;
	wire [WIDTH*2-1+3:0] tmp03_12_38;
	wire [WIDTH*2-1+3:0] tmp03_12_39;
	wire [WIDTH*2-1+3:0] tmp03_12_40;
	wire [WIDTH*2-1+3:0] tmp03_12_41;
	wire [WIDTH*2-1+3:0] tmp03_12_42;
	wire [WIDTH*2-1+3:0] tmp03_12_43;
	wire [WIDTH*2-1+3:0] tmp03_12_44;
	wire [WIDTH*2-1+3:0] tmp03_12_45;
	wire [WIDTH*2-1+3:0] tmp03_12_46;
	wire [WIDTH*2-1+3:0] tmp03_12_47;
	wire [WIDTH*2-1+3:0] tmp03_12_48;
	wire [WIDTH*2-1+3:0] tmp03_12_49;
	wire [WIDTH*2-1+3:0] tmp03_12_50;
	wire [WIDTH*2-1+3:0] tmp03_12_51;
	wire [WIDTH*2-1+3:0] tmp03_12_52;
	wire [WIDTH*2-1+3:0] tmp03_12_53;
	wire [WIDTH*2-1+3:0] tmp03_12_54;
	wire [WIDTH*2-1+3:0] tmp03_12_55;
	wire [WIDTH*2-1+3:0] tmp03_12_56;
	wire [WIDTH*2-1+3:0] tmp03_12_57;
	wire [WIDTH*2-1+3:0] tmp03_12_58;
	wire [WIDTH*2-1+3:0] tmp03_12_59;
	wire [WIDTH*2-1+3:0] tmp03_12_60;
	wire [WIDTH*2-1+3:0] tmp03_12_61;
	wire [WIDTH*2-1+3:0] tmp03_12_62;
	wire [WIDTH*2-1+3:0] tmp03_12_63;
	wire [WIDTH*2-1+3:0] tmp03_12_64;
	wire [WIDTH*2-1+3:0] tmp03_12_65;
	wire [WIDTH*2-1+3:0] tmp03_12_66;
	wire [WIDTH*2-1+3:0] tmp03_12_67;
	wire [WIDTH*2-1+3:0] tmp03_12_68;
	wire [WIDTH*2-1+3:0] tmp03_12_69;
	wire [WIDTH*2-1+3:0] tmp03_12_70;
	wire [WIDTH*2-1+3:0] tmp03_12_71;
	wire [WIDTH*2-1+3:0] tmp03_12_72;
	wire [WIDTH*2-1+3:0] tmp03_12_73;
	wire [WIDTH*2-1+3:0] tmp03_12_74;
	wire [WIDTH*2-1+3:0] tmp03_12_75;
	wire [WIDTH*2-1+3:0] tmp03_12_76;
	wire [WIDTH*2-1+3:0] tmp03_12_77;
	wire [WIDTH*2-1+3:0] tmp03_12_78;
	wire [WIDTH*2-1+3:0] tmp03_12_79;
	wire [WIDTH*2-1+3:0] tmp03_12_80;
	wire [WIDTH*2-1+3:0] tmp03_12_81;
	wire [WIDTH*2-1+3:0] tmp03_12_82;
	wire [WIDTH*2-1+3:0] tmp03_12_83;
	wire [WIDTH*2-1+3:0] tmp03_13_0;
	wire [WIDTH*2-1+3:0] tmp03_13_1;
	wire [WIDTH*2-1+3:0] tmp03_13_2;
	wire [WIDTH*2-1+3:0] tmp03_13_3;
	wire [WIDTH*2-1+3:0] tmp03_13_4;
	wire [WIDTH*2-1+3:0] tmp03_13_5;
	wire [WIDTH*2-1+3:0] tmp03_13_6;
	wire [WIDTH*2-1+3:0] tmp03_13_7;
	wire [WIDTH*2-1+3:0] tmp03_13_8;
	wire [WIDTH*2-1+3:0] tmp03_13_9;
	wire [WIDTH*2-1+3:0] tmp03_13_10;
	wire [WIDTH*2-1+3:0] tmp03_13_11;
	wire [WIDTH*2-1+3:0] tmp03_13_12;
	wire [WIDTH*2-1+3:0] tmp03_13_13;
	wire [WIDTH*2-1+3:0] tmp03_13_14;
	wire [WIDTH*2-1+3:0] tmp03_13_15;
	wire [WIDTH*2-1+3:0] tmp03_13_16;
	wire [WIDTH*2-1+3:0] tmp03_13_17;
	wire [WIDTH*2-1+3:0] tmp03_13_18;
	wire [WIDTH*2-1+3:0] tmp03_13_19;
	wire [WIDTH*2-1+3:0] tmp03_13_20;
	wire [WIDTH*2-1+3:0] tmp03_13_21;
	wire [WIDTH*2-1+3:0] tmp03_13_22;
	wire [WIDTH*2-1+3:0] tmp03_13_23;
	wire [WIDTH*2-1+3:0] tmp03_13_24;
	wire [WIDTH*2-1+3:0] tmp03_13_25;
	wire [WIDTH*2-1+3:0] tmp03_13_26;
	wire [WIDTH*2-1+3:0] tmp03_13_27;
	wire [WIDTH*2-1+3:0] tmp03_13_28;
	wire [WIDTH*2-1+3:0] tmp03_13_29;
	wire [WIDTH*2-1+3:0] tmp03_13_30;
	wire [WIDTH*2-1+3:0] tmp03_13_31;
	wire [WIDTH*2-1+3:0] tmp03_13_32;
	wire [WIDTH*2-1+3:0] tmp03_13_33;
	wire [WIDTH*2-1+3:0] tmp03_13_34;
	wire [WIDTH*2-1+3:0] tmp03_13_35;
	wire [WIDTH*2-1+3:0] tmp03_13_36;
	wire [WIDTH*2-1+3:0] tmp03_13_37;
	wire [WIDTH*2-1+3:0] tmp03_13_38;
	wire [WIDTH*2-1+3:0] tmp03_13_39;
	wire [WIDTH*2-1+3:0] tmp03_13_40;
	wire [WIDTH*2-1+3:0] tmp03_13_41;
	wire [WIDTH*2-1+3:0] tmp03_13_42;
	wire [WIDTH*2-1+3:0] tmp03_13_43;
	wire [WIDTH*2-1+3:0] tmp03_13_44;
	wire [WIDTH*2-1+3:0] tmp03_13_45;
	wire [WIDTH*2-1+3:0] tmp03_13_46;
	wire [WIDTH*2-1+3:0] tmp03_13_47;
	wire [WIDTH*2-1+3:0] tmp03_13_48;
	wire [WIDTH*2-1+3:0] tmp03_13_49;
	wire [WIDTH*2-1+3:0] tmp03_13_50;
	wire [WIDTH*2-1+3:0] tmp03_13_51;
	wire [WIDTH*2-1+3:0] tmp03_13_52;
	wire [WIDTH*2-1+3:0] tmp03_13_53;
	wire [WIDTH*2-1+3:0] tmp03_13_54;
	wire [WIDTH*2-1+3:0] tmp03_13_55;
	wire [WIDTH*2-1+3:0] tmp03_13_56;
	wire [WIDTH*2-1+3:0] tmp03_13_57;
	wire [WIDTH*2-1+3:0] tmp03_13_58;
	wire [WIDTH*2-1+3:0] tmp03_13_59;
	wire [WIDTH*2-1+3:0] tmp03_13_60;
	wire [WIDTH*2-1+3:0] tmp03_13_61;
	wire [WIDTH*2-1+3:0] tmp03_13_62;
	wire [WIDTH*2-1+3:0] tmp03_13_63;
	wire [WIDTH*2-1+3:0] tmp03_13_64;
	wire [WIDTH*2-1+3:0] tmp03_13_65;
	wire [WIDTH*2-1+3:0] tmp03_13_66;
	wire [WIDTH*2-1+3:0] tmp03_13_67;
	wire [WIDTH*2-1+3:0] tmp03_13_68;
	wire [WIDTH*2-1+3:0] tmp03_13_69;
	wire [WIDTH*2-1+3:0] tmp03_13_70;
	wire [WIDTH*2-1+3:0] tmp03_13_71;
	wire [WIDTH*2-1+3:0] tmp03_13_72;
	wire [WIDTH*2-1+3:0] tmp03_13_73;
	wire [WIDTH*2-1+3:0] tmp03_13_74;
	wire [WIDTH*2-1+3:0] tmp03_13_75;
	wire [WIDTH*2-1+3:0] tmp03_13_76;
	wire [WIDTH*2-1+3:0] tmp03_13_77;
	wire [WIDTH*2-1+3:0] tmp03_13_78;
	wire [WIDTH*2-1+3:0] tmp03_13_79;
	wire [WIDTH*2-1+3:0] tmp03_13_80;
	wire [WIDTH*2-1+3:0] tmp03_13_81;
	wire [WIDTH*2-1+3:0] tmp03_13_82;
	wire [WIDTH*2-1+3:0] tmp03_13_83;
	wire [WIDTH*2-1+3:0] tmp03_14_0;
	wire [WIDTH*2-1+3:0] tmp03_14_1;
	wire [WIDTH*2-1+3:0] tmp03_14_2;
	wire [WIDTH*2-1+3:0] tmp03_14_3;
	wire [WIDTH*2-1+3:0] tmp03_14_4;
	wire [WIDTH*2-1+3:0] tmp03_14_5;
	wire [WIDTH*2-1+3:0] tmp03_14_6;
	wire [WIDTH*2-1+3:0] tmp03_14_7;
	wire [WIDTH*2-1+3:0] tmp03_14_8;
	wire [WIDTH*2-1+3:0] tmp03_14_9;
	wire [WIDTH*2-1+3:0] tmp03_14_10;
	wire [WIDTH*2-1+3:0] tmp03_14_11;
	wire [WIDTH*2-1+3:0] tmp03_14_12;
	wire [WIDTH*2-1+3:0] tmp03_14_13;
	wire [WIDTH*2-1+3:0] tmp03_14_14;
	wire [WIDTH*2-1+3:0] tmp03_14_15;
	wire [WIDTH*2-1+3:0] tmp03_14_16;
	wire [WIDTH*2-1+3:0] tmp03_14_17;
	wire [WIDTH*2-1+3:0] tmp03_14_18;
	wire [WIDTH*2-1+3:0] tmp03_14_19;
	wire [WIDTH*2-1+3:0] tmp03_14_20;
	wire [WIDTH*2-1+3:0] tmp03_14_21;
	wire [WIDTH*2-1+3:0] tmp03_14_22;
	wire [WIDTH*2-1+3:0] tmp03_14_23;
	wire [WIDTH*2-1+3:0] tmp03_14_24;
	wire [WIDTH*2-1+3:0] tmp03_14_25;
	wire [WIDTH*2-1+3:0] tmp03_14_26;
	wire [WIDTH*2-1+3:0] tmp03_14_27;
	wire [WIDTH*2-1+3:0] tmp03_14_28;
	wire [WIDTH*2-1+3:0] tmp03_14_29;
	wire [WIDTH*2-1+3:0] tmp03_14_30;
	wire [WIDTH*2-1+3:0] tmp03_14_31;
	wire [WIDTH*2-1+3:0] tmp03_14_32;
	wire [WIDTH*2-1+3:0] tmp03_14_33;
	wire [WIDTH*2-1+3:0] tmp03_14_34;
	wire [WIDTH*2-1+3:0] tmp03_14_35;
	wire [WIDTH*2-1+3:0] tmp03_14_36;
	wire [WIDTH*2-1+3:0] tmp03_14_37;
	wire [WIDTH*2-1+3:0] tmp03_14_38;
	wire [WIDTH*2-1+3:0] tmp03_14_39;
	wire [WIDTH*2-1+3:0] tmp03_14_40;
	wire [WIDTH*2-1+3:0] tmp03_14_41;
	wire [WIDTH*2-1+3:0] tmp03_14_42;
	wire [WIDTH*2-1+3:0] tmp03_14_43;
	wire [WIDTH*2-1+3:0] tmp03_14_44;
	wire [WIDTH*2-1+3:0] tmp03_14_45;
	wire [WIDTH*2-1+3:0] tmp03_14_46;
	wire [WIDTH*2-1+3:0] tmp03_14_47;
	wire [WIDTH*2-1+3:0] tmp03_14_48;
	wire [WIDTH*2-1+3:0] tmp03_14_49;
	wire [WIDTH*2-1+3:0] tmp03_14_50;
	wire [WIDTH*2-1+3:0] tmp03_14_51;
	wire [WIDTH*2-1+3:0] tmp03_14_52;
	wire [WIDTH*2-1+3:0] tmp03_14_53;
	wire [WIDTH*2-1+3:0] tmp03_14_54;
	wire [WIDTH*2-1+3:0] tmp03_14_55;
	wire [WIDTH*2-1+3:0] tmp03_14_56;
	wire [WIDTH*2-1+3:0] tmp03_14_57;
	wire [WIDTH*2-1+3:0] tmp03_14_58;
	wire [WIDTH*2-1+3:0] tmp03_14_59;
	wire [WIDTH*2-1+3:0] tmp03_14_60;
	wire [WIDTH*2-1+3:0] tmp03_14_61;
	wire [WIDTH*2-1+3:0] tmp03_14_62;
	wire [WIDTH*2-1+3:0] tmp03_14_63;
	wire [WIDTH*2-1+3:0] tmp03_14_64;
	wire [WIDTH*2-1+3:0] tmp03_14_65;
	wire [WIDTH*2-1+3:0] tmp03_14_66;
	wire [WIDTH*2-1+3:0] tmp03_14_67;
	wire [WIDTH*2-1+3:0] tmp03_14_68;
	wire [WIDTH*2-1+3:0] tmp03_14_69;
	wire [WIDTH*2-1+3:0] tmp03_14_70;
	wire [WIDTH*2-1+3:0] tmp03_14_71;
	wire [WIDTH*2-1+3:0] tmp03_14_72;
	wire [WIDTH*2-1+3:0] tmp03_14_73;
	wire [WIDTH*2-1+3:0] tmp03_14_74;
	wire [WIDTH*2-1+3:0] tmp03_14_75;
	wire [WIDTH*2-1+3:0] tmp03_14_76;
	wire [WIDTH*2-1+3:0] tmp03_14_77;
	wire [WIDTH*2-1+3:0] tmp03_14_78;
	wire [WIDTH*2-1+3:0] tmp03_14_79;
	wire [WIDTH*2-1+3:0] tmp03_14_80;
	wire [WIDTH*2-1+3:0] tmp03_14_81;
	wire [WIDTH*2-1+3:0] tmp03_14_82;
	wire [WIDTH*2-1+3:0] tmp03_14_83;
	wire [WIDTH*2-1+3:0] tmp03_15_0;
	wire [WIDTH*2-1+3:0] tmp03_15_1;
	wire [WIDTH*2-1+3:0] tmp03_15_2;
	wire [WIDTH*2-1+3:0] tmp03_15_3;
	wire [WIDTH*2-1+3:0] tmp03_15_4;
	wire [WIDTH*2-1+3:0] tmp03_15_5;
	wire [WIDTH*2-1+3:0] tmp03_15_6;
	wire [WIDTH*2-1+3:0] tmp03_15_7;
	wire [WIDTH*2-1+3:0] tmp03_15_8;
	wire [WIDTH*2-1+3:0] tmp03_15_9;
	wire [WIDTH*2-1+3:0] tmp03_15_10;
	wire [WIDTH*2-1+3:0] tmp03_15_11;
	wire [WIDTH*2-1+3:0] tmp03_15_12;
	wire [WIDTH*2-1+3:0] tmp03_15_13;
	wire [WIDTH*2-1+3:0] tmp03_15_14;
	wire [WIDTH*2-1+3:0] tmp03_15_15;
	wire [WIDTH*2-1+3:0] tmp03_15_16;
	wire [WIDTH*2-1+3:0] tmp03_15_17;
	wire [WIDTH*2-1+3:0] tmp03_15_18;
	wire [WIDTH*2-1+3:0] tmp03_15_19;
	wire [WIDTH*2-1+3:0] tmp03_15_20;
	wire [WIDTH*2-1+3:0] tmp03_15_21;
	wire [WIDTH*2-1+3:0] tmp03_15_22;
	wire [WIDTH*2-1+3:0] tmp03_15_23;
	wire [WIDTH*2-1+3:0] tmp03_15_24;
	wire [WIDTH*2-1+3:0] tmp03_15_25;
	wire [WIDTH*2-1+3:0] tmp03_15_26;
	wire [WIDTH*2-1+3:0] tmp03_15_27;
	wire [WIDTH*2-1+3:0] tmp03_15_28;
	wire [WIDTH*2-1+3:0] tmp03_15_29;
	wire [WIDTH*2-1+3:0] tmp03_15_30;
	wire [WIDTH*2-1+3:0] tmp03_15_31;
	wire [WIDTH*2-1+3:0] tmp03_15_32;
	wire [WIDTH*2-1+3:0] tmp03_15_33;
	wire [WIDTH*2-1+3:0] tmp03_15_34;
	wire [WIDTH*2-1+3:0] tmp03_15_35;
	wire [WIDTH*2-1+3:0] tmp03_15_36;
	wire [WIDTH*2-1+3:0] tmp03_15_37;
	wire [WIDTH*2-1+3:0] tmp03_15_38;
	wire [WIDTH*2-1+3:0] tmp03_15_39;
	wire [WIDTH*2-1+3:0] tmp03_15_40;
	wire [WIDTH*2-1+3:0] tmp03_15_41;
	wire [WIDTH*2-1+3:0] tmp03_15_42;
	wire [WIDTH*2-1+3:0] tmp03_15_43;
	wire [WIDTH*2-1+3:0] tmp03_15_44;
	wire [WIDTH*2-1+3:0] tmp03_15_45;
	wire [WIDTH*2-1+3:0] tmp03_15_46;
	wire [WIDTH*2-1+3:0] tmp03_15_47;
	wire [WIDTH*2-1+3:0] tmp03_15_48;
	wire [WIDTH*2-1+3:0] tmp03_15_49;
	wire [WIDTH*2-1+3:0] tmp03_15_50;
	wire [WIDTH*2-1+3:0] tmp03_15_51;
	wire [WIDTH*2-1+3:0] tmp03_15_52;
	wire [WIDTH*2-1+3:0] tmp03_15_53;
	wire [WIDTH*2-1+3:0] tmp03_15_54;
	wire [WIDTH*2-1+3:0] tmp03_15_55;
	wire [WIDTH*2-1+3:0] tmp03_15_56;
	wire [WIDTH*2-1+3:0] tmp03_15_57;
	wire [WIDTH*2-1+3:0] tmp03_15_58;
	wire [WIDTH*2-1+3:0] tmp03_15_59;
	wire [WIDTH*2-1+3:0] tmp03_15_60;
	wire [WIDTH*2-1+3:0] tmp03_15_61;
	wire [WIDTH*2-1+3:0] tmp03_15_62;
	wire [WIDTH*2-1+3:0] tmp03_15_63;
	wire [WIDTH*2-1+3:0] tmp03_15_64;
	wire [WIDTH*2-1+3:0] tmp03_15_65;
	wire [WIDTH*2-1+3:0] tmp03_15_66;
	wire [WIDTH*2-1+3:0] tmp03_15_67;
	wire [WIDTH*2-1+3:0] tmp03_15_68;
	wire [WIDTH*2-1+3:0] tmp03_15_69;
	wire [WIDTH*2-1+3:0] tmp03_15_70;
	wire [WIDTH*2-1+3:0] tmp03_15_71;
	wire [WIDTH*2-1+3:0] tmp03_15_72;
	wire [WIDTH*2-1+3:0] tmp03_15_73;
	wire [WIDTH*2-1+3:0] tmp03_15_74;
	wire [WIDTH*2-1+3:0] tmp03_15_75;
	wire [WIDTH*2-1+3:0] tmp03_15_76;
	wire [WIDTH*2-1+3:0] tmp03_15_77;
	wire [WIDTH*2-1+3:0] tmp03_15_78;
	wire [WIDTH*2-1+3:0] tmp03_15_79;
	wire [WIDTH*2-1+3:0] tmp03_15_80;
	wire [WIDTH*2-1+3:0] tmp03_15_81;
	wire [WIDTH*2-1+3:0] tmp03_15_82;
	wire [WIDTH*2-1+3:0] tmp03_15_83;
	wire [WIDTH*2-1+4:0] tmp04_0_0;
	wire [WIDTH*2-1+4:0] tmp04_0_1;
	wire [WIDTH*2-1+4:0] tmp04_0_2;
	wire [WIDTH*2-1+4:0] tmp04_0_3;
	wire [WIDTH*2-1+4:0] tmp04_0_4;
	wire [WIDTH*2-1+4:0] tmp04_0_5;
	wire [WIDTH*2-1+4:0] tmp04_0_6;
	wire [WIDTH*2-1+4:0] tmp04_0_7;
	wire [WIDTH*2-1+4:0] tmp04_0_8;
	wire [WIDTH*2-1+4:0] tmp04_0_9;
	wire [WIDTH*2-1+4:0] tmp04_0_10;
	wire [WIDTH*2-1+4:0] tmp04_0_11;
	wire [WIDTH*2-1+4:0] tmp04_0_12;
	wire [WIDTH*2-1+4:0] tmp04_0_13;
	wire [WIDTH*2-1+4:0] tmp04_0_14;
	wire [WIDTH*2-1+4:0] tmp04_0_15;
	wire [WIDTH*2-1+4:0] tmp04_0_16;
	wire [WIDTH*2-1+4:0] tmp04_0_17;
	wire [WIDTH*2-1+4:0] tmp04_0_18;
	wire [WIDTH*2-1+4:0] tmp04_0_19;
	wire [WIDTH*2-1+4:0] tmp04_0_20;
	wire [WIDTH*2-1+4:0] tmp04_0_21;
	wire [WIDTH*2-1+4:0] tmp04_0_22;
	wire [WIDTH*2-1+4:0] tmp04_0_23;
	wire [WIDTH*2-1+4:0] tmp04_0_24;
	wire [WIDTH*2-1+4:0] tmp04_0_25;
	wire [WIDTH*2-1+4:0] tmp04_0_26;
	wire [WIDTH*2-1+4:0] tmp04_0_27;
	wire [WIDTH*2-1+4:0] tmp04_0_28;
	wire [WIDTH*2-1+4:0] tmp04_0_29;
	wire [WIDTH*2-1+4:0] tmp04_0_30;
	wire [WIDTH*2-1+4:0] tmp04_0_31;
	wire [WIDTH*2-1+4:0] tmp04_0_32;
	wire [WIDTH*2-1+4:0] tmp04_0_33;
	wire [WIDTH*2-1+4:0] tmp04_0_34;
	wire [WIDTH*2-1+4:0] tmp04_0_35;
	wire [WIDTH*2-1+4:0] tmp04_0_36;
	wire [WIDTH*2-1+4:0] tmp04_0_37;
	wire [WIDTH*2-1+4:0] tmp04_0_38;
	wire [WIDTH*2-1+4:0] tmp04_0_39;
	wire [WIDTH*2-1+4:0] tmp04_0_40;
	wire [WIDTH*2-1+4:0] tmp04_0_41;
	wire [WIDTH*2-1+4:0] tmp04_0_42;
	wire [WIDTH*2-1+4:0] tmp04_0_43;
	wire [WIDTH*2-1+4:0] tmp04_0_44;
	wire [WIDTH*2-1+4:0] tmp04_0_45;
	wire [WIDTH*2-1+4:0] tmp04_0_46;
	wire [WIDTH*2-1+4:0] tmp04_0_47;
	wire [WIDTH*2-1+4:0] tmp04_0_48;
	wire [WIDTH*2-1+4:0] tmp04_0_49;
	wire [WIDTH*2-1+4:0] tmp04_0_50;
	wire [WIDTH*2-1+4:0] tmp04_0_51;
	wire [WIDTH*2-1+4:0] tmp04_0_52;
	wire [WIDTH*2-1+4:0] tmp04_0_53;
	wire [WIDTH*2-1+4:0] tmp04_0_54;
	wire [WIDTH*2-1+4:0] tmp04_0_55;
	wire [WIDTH*2-1+4:0] tmp04_0_56;
	wire [WIDTH*2-1+4:0] tmp04_0_57;
	wire [WIDTH*2-1+4:0] tmp04_0_58;
	wire [WIDTH*2-1+4:0] tmp04_0_59;
	wire [WIDTH*2-1+4:0] tmp04_0_60;
	wire [WIDTH*2-1+4:0] tmp04_0_61;
	wire [WIDTH*2-1+4:0] tmp04_0_62;
	wire [WIDTH*2-1+4:0] tmp04_0_63;
	wire [WIDTH*2-1+4:0] tmp04_0_64;
	wire [WIDTH*2-1+4:0] tmp04_0_65;
	wire [WIDTH*2-1+4:0] tmp04_0_66;
	wire [WIDTH*2-1+4:0] tmp04_0_67;
	wire [WIDTH*2-1+4:0] tmp04_0_68;
	wire [WIDTH*2-1+4:0] tmp04_0_69;
	wire [WIDTH*2-1+4:0] tmp04_0_70;
	wire [WIDTH*2-1+4:0] tmp04_0_71;
	wire [WIDTH*2-1+4:0] tmp04_0_72;
	wire [WIDTH*2-1+4:0] tmp04_0_73;
	wire [WIDTH*2-1+4:0] tmp04_0_74;
	wire [WIDTH*2-1+4:0] tmp04_0_75;
	wire [WIDTH*2-1+4:0] tmp04_0_76;
	wire [WIDTH*2-1+4:0] tmp04_0_77;
	wire [WIDTH*2-1+4:0] tmp04_0_78;
	wire [WIDTH*2-1+4:0] tmp04_0_79;
	wire [WIDTH*2-1+4:0] tmp04_0_80;
	wire [WIDTH*2-1+4:0] tmp04_0_81;
	wire [WIDTH*2-1+4:0] tmp04_0_82;
	wire [WIDTH*2-1+4:0] tmp04_0_83;
	wire [WIDTH*2-1+4:0] tmp04_1_0;
	wire [WIDTH*2-1+4:0] tmp04_1_1;
	wire [WIDTH*2-1+4:0] tmp04_1_2;
	wire [WIDTH*2-1+4:0] tmp04_1_3;
	wire [WIDTH*2-1+4:0] tmp04_1_4;
	wire [WIDTH*2-1+4:0] tmp04_1_5;
	wire [WIDTH*2-1+4:0] tmp04_1_6;
	wire [WIDTH*2-1+4:0] tmp04_1_7;
	wire [WIDTH*2-1+4:0] tmp04_1_8;
	wire [WIDTH*2-1+4:0] tmp04_1_9;
	wire [WIDTH*2-1+4:0] tmp04_1_10;
	wire [WIDTH*2-1+4:0] tmp04_1_11;
	wire [WIDTH*2-1+4:0] tmp04_1_12;
	wire [WIDTH*2-1+4:0] tmp04_1_13;
	wire [WIDTH*2-1+4:0] tmp04_1_14;
	wire [WIDTH*2-1+4:0] tmp04_1_15;
	wire [WIDTH*2-1+4:0] tmp04_1_16;
	wire [WIDTH*2-1+4:0] tmp04_1_17;
	wire [WIDTH*2-1+4:0] tmp04_1_18;
	wire [WIDTH*2-1+4:0] tmp04_1_19;
	wire [WIDTH*2-1+4:0] tmp04_1_20;
	wire [WIDTH*2-1+4:0] tmp04_1_21;
	wire [WIDTH*2-1+4:0] tmp04_1_22;
	wire [WIDTH*2-1+4:0] tmp04_1_23;
	wire [WIDTH*2-1+4:0] tmp04_1_24;
	wire [WIDTH*2-1+4:0] tmp04_1_25;
	wire [WIDTH*2-1+4:0] tmp04_1_26;
	wire [WIDTH*2-1+4:0] tmp04_1_27;
	wire [WIDTH*2-1+4:0] tmp04_1_28;
	wire [WIDTH*2-1+4:0] tmp04_1_29;
	wire [WIDTH*2-1+4:0] tmp04_1_30;
	wire [WIDTH*2-1+4:0] tmp04_1_31;
	wire [WIDTH*2-1+4:0] tmp04_1_32;
	wire [WIDTH*2-1+4:0] tmp04_1_33;
	wire [WIDTH*2-1+4:0] tmp04_1_34;
	wire [WIDTH*2-1+4:0] tmp04_1_35;
	wire [WIDTH*2-1+4:0] tmp04_1_36;
	wire [WIDTH*2-1+4:0] tmp04_1_37;
	wire [WIDTH*2-1+4:0] tmp04_1_38;
	wire [WIDTH*2-1+4:0] tmp04_1_39;
	wire [WIDTH*2-1+4:0] tmp04_1_40;
	wire [WIDTH*2-1+4:0] tmp04_1_41;
	wire [WIDTH*2-1+4:0] tmp04_1_42;
	wire [WIDTH*2-1+4:0] tmp04_1_43;
	wire [WIDTH*2-1+4:0] tmp04_1_44;
	wire [WIDTH*2-1+4:0] tmp04_1_45;
	wire [WIDTH*2-1+4:0] tmp04_1_46;
	wire [WIDTH*2-1+4:0] tmp04_1_47;
	wire [WIDTH*2-1+4:0] tmp04_1_48;
	wire [WIDTH*2-1+4:0] tmp04_1_49;
	wire [WIDTH*2-1+4:0] tmp04_1_50;
	wire [WIDTH*2-1+4:0] tmp04_1_51;
	wire [WIDTH*2-1+4:0] tmp04_1_52;
	wire [WIDTH*2-1+4:0] tmp04_1_53;
	wire [WIDTH*2-1+4:0] tmp04_1_54;
	wire [WIDTH*2-1+4:0] tmp04_1_55;
	wire [WIDTH*2-1+4:0] tmp04_1_56;
	wire [WIDTH*2-1+4:0] tmp04_1_57;
	wire [WIDTH*2-1+4:0] tmp04_1_58;
	wire [WIDTH*2-1+4:0] tmp04_1_59;
	wire [WIDTH*2-1+4:0] tmp04_1_60;
	wire [WIDTH*2-1+4:0] tmp04_1_61;
	wire [WIDTH*2-1+4:0] tmp04_1_62;
	wire [WIDTH*2-1+4:0] tmp04_1_63;
	wire [WIDTH*2-1+4:0] tmp04_1_64;
	wire [WIDTH*2-1+4:0] tmp04_1_65;
	wire [WIDTH*2-1+4:0] tmp04_1_66;
	wire [WIDTH*2-1+4:0] tmp04_1_67;
	wire [WIDTH*2-1+4:0] tmp04_1_68;
	wire [WIDTH*2-1+4:0] tmp04_1_69;
	wire [WIDTH*2-1+4:0] tmp04_1_70;
	wire [WIDTH*2-1+4:0] tmp04_1_71;
	wire [WIDTH*2-1+4:0] tmp04_1_72;
	wire [WIDTH*2-1+4:0] tmp04_1_73;
	wire [WIDTH*2-1+4:0] tmp04_1_74;
	wire [WIDTH*2-1+4:0] tmp04_1_75;
	wire [WIDTH*2-1+4:0] tmp04_1_76;
	wire [WIDTH*2-1+4:0] tmp04_1_77;
	wire [WIDTH*2-1+4:0] tmp04_1_78;
	wire [WIDTH*2-1+4:0] tmp04_1_79;
	wire [WIDTH*2-1+4:0] tmp04_1_80;
	wire [WIDTH*2-1+4:0] tmp04_1_81;
	wire [WIDTH*2-1+4:0] tmp04_1_82;
	wire [WIDTH*2-1+4:0] tmp04_1_83;
	wire [WIDTH*2-1+4:0] tmp04_2_0;
	wire [WIDTH*2-1+4:0] tmp04_2_1;
	wire [WIDTH*2-1+4:0] tmp04_2_2;
	wire [WIDTH*2-1+4:0] tmp04_2_3;
	wire [WIDTH*2-1+4:0] tmp04_2_4;
	wire [WIDTH*2-1+4:0] tmp04_2_5;
	wire [WIDTH*2-1+4:0] tmp04_2_6;
	wire [WIDTH*2-1+4:0] tmp04_2_7;
	wire [WIDTH*2-1+4:0] tmp04_2_8;
	wire [WIDTH*2-1+4:0] tmp04_2_9;
	wire [WIDTH*2-1+4:0] tmp04_2_10;
	wire [WIDTH*2-1+4:0] tmp04_2_11;
	wire [WIDTH*2-1+4:0] tmp04_2_12;
	wire [WIDTH*2-1+4:0] tmp04_2_13;
	wire [WIDTH*2-1+4:0] tmp04_2_14;
	wire [WIDTH*2-1+4:0] tmp04_2_15;
	wire [WIDTH*2-1+4:0] tmp04_2_16;
	wire [WIDTH*2-1+4:0] tmp04_2_17;
	wire [WIDTH*2-1+4:0] tmp04_2_18;
	wire [WIDTH*2-1+4:0] tmp04_2_19;
	wire [WIDTH*2-1+4:0] tmp04_2_20;
	wire [WIDTH*2-1+4:0] tmp04_2_21;
	wire [WIDTH*2-1+4:0] tmp04_2_22;
	wire [WIDTH*2-1+4:0] tmp04_2_23;
	wire [WIDTH*2-1+4:0] tmp04_2_24;
	wire [WIDTH*2-1+4:0] tmp04_2_25;
	wire [WIDTH*2-1+4:0] tmp04_2_26;
	wire [WIDTH*2-1+4:0] tmp04_2_27;
	wire [WIDTH*2-1+4:0] tmp04_2_28;
	wire [WIDTH*2-1+4:0] tmp04_2_29;
	wire [WIDTH*2-1+4:0] tmp04_2_30;
	wire [WIDTH*2-1+4:0] tmp04_2_31;
	wire [WIDTH*2-1+4:0] tmp04_2_32;
	wire [WIDTH*2-1+4:0] tmp04_2_33;
	wire [WIDTH*2-1+4:0] tmp04_2_34;
	wire [WIDTH*2-1+4:0] tmp04_2_35;
	wire [WIDTH*2-1+4:0] tmp04_2_36;
	wire [WIDTH*2-1+4:0] tmp04_2_37;
	wire [WIDTH*2-1+4:0] tmp04_2_38;
	wire [WIDTH*2-1+4:0] tmp04_2_39;
	wire [WIDTH*2-1+4:0] tmp04_2_40;
	wire [WIDTH*2-1+4:0] tmp04_2_41;
	wire [WIDTH*2-1+4:0] tmp04_2_42;
	wire [WIDTH*2-1+4:0] tmp04_2_43;
	wire [WIDTH*2-1+4:0] tmp04_2_44;
	wire [WIDTH*2-1+4:0] tmp04_2_45;
	wire [WIDTH*2-1+4:0] tmp04_2_46;
	wire [WIDTH*2-1+4:0] tmp04_2_47;
	wire [WIDTH*2-1+4:0] tmp04_2_48;
	wire [WIDTH*2-1+4:0] tmp04_2_49;
	wire [WIDTH*2-1+4:0] tmp04_2_50;
	wire [WIDTH*2-1+4:0] tmp04_2_51;
	wire [WIDTH*2-1+4:0] tmp04_2_52;
	wire [WIDTH*2-1+4:0] tmp04_2_53;
	wire [WIDTH*2-1+4:0] tmp04_2_54;
	wire [WIDTH*2-1+4:0] tmp04_2_55;
	wire [WIDTH*2-1+4:0] tmp04_2_56;
	wire [WIDTH*2-1+4:0] tmp04_2_57;
	wire [WIDTH*2-1+4:0] tmp04_2_58;
	wire [WIDTH*2-1+4:0] tmp04_2_59;
	wire [WIDTH*2-1+4:0] tmp04_2_60;
	wire [WIDTH*2-1+4:0] tmp04_2_61;
	wire [WIDTH*2-1+4:0] tmp04_2_62;
	wire [WIDTH*2-1+4:0] tmp04_2_63;
	wire [WIDTH*2-1+4:0] tmp04_2_64;
	wire [WIDTH*2-1+4:0] tmp04_2_65;
	wire [WIDTH*2-1+4:0] tmp04_2_66;
	wire [WIDTH*2-1+4:0] tmp04_2_67;
	wire [WIDTH*2-1+4:0] tmp04_2_68;
	wire [WIDTH*2-1+4:0] tmp04_2_69;
	wire [WIDTH*2-1+4:0] tmp04_2_70;
	wire [WIDTH*2-1+4:0] tmp04_2_71;
	wire [WIDTH*2-1+4:0] tmp04_2_72;
	wire [WIDTH*2-1+4:0] tmp04_2_73;
	wire [WIDTH*2-1+4:0] tmp04_2_74;
	wire [WIDTH*2-1+4:0] tmp04_2_75;
	wire [WIDTH*2-1+4:0] tmp04_2_76;
	wire [WIDTH*2-1+4:0] tmp04_2_77;
	wire [WIDTH*2-1+4:0] tmp04_2_78;
	wire [WIDTH*2-1+4:0] tmp04_2_79;
	wire [WIDTH*2-1+4:0] tmp04_2_80;
	wire [WIDTH*2-1+4:0] tmp04_2_81;
	wire [WIDTH*2-1+4:0] tmp04_2_82;
	wire [WIDTH*2-1+4:0] tmp04_2_83;
	wire [WIDTH*2-1+4:0] tmp04_3_0;
	wire [WIDTH*2-1+4:0] tmp04_3_1;
	wire [WIDTH*2-1+4:0] tmp04_3_2;
	wire [WIDTH*2-1+4:0] tmp04_3_3;
	wire [WIDTH*2-1+4:0] tmp04_3_4;
	wire [WIDTH*2-1+4:0] tmp04_3_5;
	wire [WIDTH*2-1+4:0] tmp04_3_6;
	wire [WIDTH*2-1+4:0] tmp04_3_7;
	wire [WIDTH*2-1+4:0] tmp04_3_8;
	wire [WIDTH*2-1+4:0] tmp04_3_9;
	wire [WIDTH*2-1+4:0] tmp04_3_10;
	wire [WIDTH*2-1+4:0] tmp04_3_11;
	wire [WIDTH*2-1+4:0] tmp04_3_12;
	wire [WIDTH*2-1+4:0] tmp04_3_13;
	wire [WIDTH*2-1+4:0] tmp04_3_14;
	wire [WIDTH*2-1+4:0] tmp04_3_15;
	wire [WIDTH*2-1+4:0] tmp04_3_16;
	wire [WIDTH*2-1+4:0] tmp04_3_17;
	wire [WIDTH*2-1+4:0] tmp04_3_18;
	wire [WIDTH*2-1+4:0] tmp04_3_19;
	wire [WIDTH*2-1+4:0] tmp04_3_20;
	wire [WIDTH*2-1+4:0] tmp04_3_21;
	wire [WIDTH*2-1+4:0] tmp04_3_22;
	wire [WIDTH*2-1+4:0] tmp04_3_23;
	wire [WIDTH*2-1+4:0] tmp04_3_24;
	wire [WIDTH*2-1+4:0] tmp04_3_25;
	wire [WIDTH*2-1+4:0] tmp04_3_26;
	wire [WIDTH*2-1+4:0] tmp04_3_27;
	wire [WIDTH*2-1+4:0] tmp04_3_28;
	wire [WIDTH*2-1+4:0] tmp04_3_29;
	wire [WIDTH*2-1+4:0] tmp04_3_30;
	wire [WIDTH*2-1+4:0] tmp04_3_31;
	wire [WIDTH*2-1+4:0] tmp04_3_32;
	wire [WIDTH*2-1+4:0] tmp04_3_33;
	wire [WIDTH*2-1+4:0] tmp04_3_34;
	wire [WIDTH*2-1+4:0] tmp04_3_35;
	wire [WIDTH*2-1+4:0] tmp04_3_36;
	wire [WIDTH*2-1+4:0] tmp04_3_37;
	wire [WIDTH*2-1+4:0] tmp04_3_38;
	wire [WIDTH*2-1+4:0] tmp04_3_39;
	wire [WIDTH*2-1+4:0] tmp04_3_40;
	wire [WIDTH*2-1+4:0] tmp04_3_41;
	wire [WIDTH*2-1+4:0] tmp04_3_42;
	wire [WIDTH*2-1+4:0] tmp04_3_43;
	wire [WIDTH*2-1+4:0] tmp04_3_44;
	wire [WIDTH*2-1+4:0] tmp04_3_45;
	wire [WIDTH*2-1+4:0] tmp04_3_46;
	wire [WIDTH*2-1+4:0] tmp04_3_47;
	wire [WIDTH*2-1+4:0] tmp04_3_48;
	wire [WIDTH*2-1+4:0] tmp04_3_49;
	wire [WIDTH*2-1+4:0] tmp04_3_50;
	wire [WIDTH*2-1+4:0] tmp04_3_51;
	wire [WIDTH*2-1+4:0] tmp04_3_52;
	wire [WIDTH*2-1+4:0] tmp04_3_53;
	wire [WIDTH*2-1+4:0] tmp04_3_54;
	wire [WIDTH*2-1+4:0] tmp04_3_55;
	wire [WIDTH*2-1+4:0] tmp04_3_56;
	wire [WIDTH*2-1+4:0] tmp04_3_57;
	wire [WIDTH*2-1+4:0] tmp04_3_58;
	wire [WIDTH*2-1+4:0] tmp04_3_59;
	wire [WIDTH*2-1+4:0] tmp04_3_60;
	wire [WIDTH*2-1+4:0] tmp04_3_61;
	wire [WIDTH*2-1+4:0] tmp04_3_62;
	wire [WIDTH*2-1+4:0] tmp04_3_63;
	wire [WIDTH*2-1+4:0] tmp04_3_64;
	wire [WIDTH*2-1+4:0] tmp04_3_65;
	wire [WIDTH*2-1+4:0] tmp04_3_66;
	wire [WIDTH*2-1+4:0] tmp04_3_67;
	wire [WIDTH*2-1+4:0] tmp04_3_68;
	wire [WIDTH*2-1+4:0] tmp04_3_69;
	wire [WIDTH*2-1+4:0] tmp04_3_70;
	wire [WIDTH*2-1+4:0] tmp04_3_71;
	wire [WIDTH*2-1+4:0] tmp04_3_72;
	wire [WIDTH*2-1+4:0] tmp04_3_73;
	wire [WIDTH*2-1+4:0] tmp04_3_74;
	wire [WIDTH*2-1+4:0] tmp04_3_75;
	wire [WIDTH*2-1+4:0] tmp04_3_76;
	wire [WIDTH*2-1+4:0] tmp04_3_77;
	wire [WIDTH*2-1+4:0] tmp04_3_78;
	wire [WIDTH*2-1+4:0] tmp04_3_79;
	wire [WIDTH*2-1+4:0] tmp04_3_80;
	wire [WIDTH*2-1+4:0] tmp04_3_81;
	wire [WIDTH*2-1+4:0] tmp04_3_82;
	wire [WIDTH*2-1+4:0] tmp04_3_83;
	wire [WIDTH*2-1+4:0] tmp04_4_0;
	wire [WIDTH*2-1+4:0] tmp04_4_1;
	wire [WIDTH*2-1+4:0] tmp04_4_2;
	wire [WIDTH*2-1+4:0] tmp04_4_3;
	wire [WIDTH*2-1+4:0] tmp04_4_4;
	wire [WIDTH*2-1+4:0] tmp04_4_5;
	wire [WIDTH*2-1+4:0] tmp04_4_6;
	wire [WIDTH*2-1+4:0] tmp04_4_7;
	wire [WIDTH*2-1+4:0] tmp04_4_8;
	wire [WIDTH*2-1+4:0] tmp04_4_9;
	wire [WIDTH*2-1+4:0] tmp04_4_10;
	wire [WIDTH*2-1+4:0] tmp04_4_11;
	wire [WIDTH*2-1+4:0] tmp04_4_12;
	wire [WIDTH*2-1+4:0] tmp04_4_13;
	wire [WIDTH*2-1+4:0] tmp04_4_14;
	wire [WIDTH*2-1+4:0] tmp04_4_15;
	wire [WIDTH*2-1+4:0] tmp04_4_16;
	wire [WIDTH*2-1+4:0] tmp04_4_17;
	wire [WIDTH*2-1+4:0] tmp04_4_18;
	wire [WIDTH*2-1+4:0] tmp04_4_19;
	wire [WIDTH*2-1+4:0] tmp04_4_20;
	wire [WIDTH*2-1+4:0] tmp04_4_21;
	wire [WIDTH*2-1+4:0] tmp04_4_22;
	wire [WIDTH*2-1+4:0] tmp04_4_23;
	wire [WIDTH*2-1+4:0] tmp04_4_24;
	wire [WIDTH*2-1+4:0] tmp04_4_25;
	wire [WIDTH*2-1+4:0] tmp04_4_26;
	wire [WIDTH*2-1+4:0] tmp04_4_27;
	wire [WIDTH*2-1+4:0] tmp04_4_28;
	wire [WIDTH*2-1+4:0] tmp04_4_29;
	wire [WIDTH*2-1+4:0] tmp04_4_30;
	wire [WIDTH*2-1+4:0] tmp04_4_31;
	wire [WIDTH*2-1+4:0] tmp04_4_32;
	wire [WIDTH*2-1+4:0] tmp04_4_33;
	wire [WIDTH*2-1+4:0] tmp04_4_34;
	wire [WIDTH*2-1+4:0] tmp04_4_35;
	wire [WIDTH*2-1+4:0] tmp04_4_36;
	wire [WIDTH*2-1+4:0] tmp04_4_37;
	wire [WIDTH*2-1+4:0] tmp04_4_38;
	wire [WIDTH*2-1+4:0] tmp04_4_39;
	wire [WIDTH*2-1+4:0] tmp04_4_40;
	wire [WIDTH*2-1+4:0] tmp04_4_41;
	wire [WIDTH*2-1+4:0] tmp04_4_42;
	wire [WIDTH*2-1+4:0] tmp04_4_43;
	wire [WIDTH*2-1+4:0] tmp04_4_44;
	wire [WIDTH*2-1+4:0] tmp04_4_45;
	wire [WIDTH*2-1+4:0] tmp04_4_46;
	wire [WIDTH*2-1+4:0] tmp04_4_47;
	wire [WIDTH*2-1+4:0] tmp04_4_48;
	wire [WIDTH*2-1+4:0] tmp04_4_49;
	wire [WIDTH*2-1+4:0] tmp04_4_50;
	wire [WIDTH*2-1+4:0] tmp04_4_51;
	wire [WIDTH*2-1+4:0] tmp04_4_52;
	wire [WIDTH*2-1+4:0] tmp04_4_53;
	wire [WIDTH*2-1+4:0] tmp04_4_54;
	wire [WIDTH*2-1+4:0] tmp04_4_55;
	wire [WIDTH*2-1+4:0] tmp04_4_56;
	wire [WIDTH*2-1+4:0] tmp04_4_57;
	wire [WIDTH*2-1+4:0] tmp04_4_58;
	wire [WIDTH*2-1+4:0] tmp04_4_59;
	wire [WIDTH*2-1+4:0] tmp04_4_60;
	wire [WIDTH*2-1+4:0] tmp04_4_61;
	wire [WIDTH*2-1+4:0] tmp04_4_62;
	wire [WIDTH*2-1+4:0] tmp04_4_63;
	wire [WIDTH*2-1+4:0] tmp04_4_64;
	wire [WIDTH*2-1+4:0] tmp04_4_65;
	wire [WIDTH*2-1+4:0] tmp04_4_66;
	wire [WIDTH*2-1+4:0] tmp04_4_67;
	wire [WIDTH*2-1+4:0] tmp04_4_68;
	wire [WIDTH*2-1+4:0] tmp04_4_69;
	wire [WIDTH*2-1+4:0] tmp04_4_70;
	wire [WIDTH*2-1+4:0] tmp04_4_71;
	wire [WIDTH*2-1+4:0] tmp04_4_72;
	wire [WIDTH*2-1+4:0] tmp04_4_73;
	wire [WIDTH*2-1+4:0] tmp04_4_74;
	wire [WIDTH*2-1+4:0] tmp04_4_75;
	wire [WIDTH*2-1+4:0] tmp04_4_76;
	wire [WIDTH*2-1+4:0] tmp04_4_77;
	wire [WIDTH*2-1+4:0] tmp04_4_78;
	wire [WIDTH*2-1+4:0] tmp04_4_79;
	wire [WIDTH*2-1+4:0] tmp04_4_80;
	wire [WIDTH*2-1+4:0] tmp04_4_81;
	wire [WIDTH*2-1+4:0] tmp04_4_82;
	wire [WIDTH*2-1+4:0] tmp04_4_83;
	wire [WIDTH*2-1+4:0] tmp04_5_0;
	wire [WIDTH*2-1+4:0] tmp04_5_1;
	wire [WIDTH*2-1+4:0] tmp04_5_2;
	wire [WIDTH*2-1+4:0] tmp04_5_3;
	wire [WIDTH*2-1+4:0] tmp04_5_4;
	wire [WIDTH*2-1+4:0] tmp04_5_5;
	wire [WIDTH*2-1+4:0] tmp04_5_6;
	wire [WIDTH*2-1+4:0] tmp04_5_7;
	wire [WIDTH*2-1+4:0] tmp04_5_8;
	wire [WIDTH*2-1+4:0] tmp04_5_9;
	wire [WIDTH*2-1+4:0] tmp04_5_10;
	wire [WIDTH*2-1+4:0] tmp04_5_11;
	wire [WIDTH*2-1+4:0] tmp04_5_12;
	wire [WIDTH*2-1+4:0] tmp04_5_13;
	wire [WIDTH*2-1+4:0] tmp04_5_14;
	wire [WIDTH*2-1+4:0] tmp04_5_15;
	wire [WIDTH*2-1+4:0] tmp04_5_16;
	wire [WIDTH*2-1+4:0] tmp04_5_17;
	wire [WIDTH*2-1+4:0] tmp04_5_18;
	wire [WIDTH*2-1+4:0] tmp04_5_19;
	wire [WIDTH*2-1+4:0] tmp04_5_20;
	wire [WIDTH*2-1+4:0] tmp04_5_21;
	wire [WIDTH*2-1+4:0] tmp04_5_22;
	wire [WIDTH*2-1+4:0] tmp04_5_23;
	wire [WIDTH*2-1+4:0] tmp04_5_24;
	wire [WIDTH*2-1+4:0] tmp04_5_25;
	wire [WIDTH*2-1+4:0] tmp04_5_26;
	wire [WIDTH*2-1+4:0] tmp04_5_27;
	wire [WIDTH*2-1+4:0] tmp04_5_28;
	wire [WIDTH*2-1+4:0] tmp04_5_29;
	wire [WIDTH*2-1+4:0] tmp04_5_30;
	wire [WIDTH*2-1+4:0] tmp04_5_31;
	wire [WIDTH*2-1+4:0] tmp04_5_32;
	wire [WIDTH*2-1+4:0] tmp04_5_33;
	wire [WIDTH*2-1+4:0] tmp04_5_34;
	wire [WIDTH*2-1+4:0] tmp04_5_35;
	wire [WIDTH*2-1+4:0] tmp04_5_36;
	wire [WIDTH*2-1+4:0] tmp04_5_37;
	wire [WIDTH*2-1+4:0] tmp04_5_38;
	wire [WIDTH*2-1+4:0] tmp04_5_39;
	wire [WIDTH*2-1+4:0] tmp04_5_40;
	wire [WIDTH*2-1+4:0] tmp04_5_41;
	wire [WIDTH*2-1+4:0] tmp04_5_42;
	wire [WIDTH*2-1+4:0] tmp04_5_43;
	wire [WIDTH*2-1+4:0] tmp04_5_44;
	wire [WIDTH*2-1+4:0] tmp04_5_45;
	wire [WIDTH*2-1+4:0] tmp04_5_46;
	wire [WIDTH*2-1+4:0] tmp04_5_47;
	wire [WIDTH*2-1+4:0] tmp04_5_48;
	wire [WIDTH*2-1+4:0] tmp04_5_49;
	wire [WIDTH*2-1+4:0] tmp04_5_50;
	wire [WIDTH*2-1+4:0] tmp04_5_51;
	wire [WIDTH*2-1+4:0] tmp04_5_52;
	wire [WIDTH*2-1+4:0] tmp04_5_53;
	wire [WIDTH*2-1+4:0] tmp04_5_54;
	wire [WIDTH*2-1+4:0] tmp04_5_55;
	wire [WIDTH*2-1+4:0] tmp04_5_56;
	wire [WIDTH*2-1+4:0] tmp04_5_57;
	wire [WIDTH*2-1+4:0] tmp04_5_58;
	wire [WIDTH*2-1+4:0] tmp04_5_59;
	wire [WIDTH*2-1+4:0] tmp04_5_60;
	wire [WIDTH*2-1+4:0] tmp04_5_61;
	wire [WIDTH*2-1+4:0] tmp04_5_62;
	wire [WIDTH*2-1+4:0] tmp04_5_63;
	wire [WIDTH*2-1+4:0] tmp04_5_64;
	wire [WIDTH*2-1+4:0] tmp04_5_65;
	wire [WIDTH*2-1+4:0] tmp04_5_66;
	wire [WIDTH*2-1+4:0] tmp04_5_67;
	wire [WIDTH*2-1+4:0] tmp04_5_68;
	wire [WIDTH*2-1+4:0] tmp04_5_69;
	wire [WIDTH*2-1+4:0] tmp04_5_70;
	wire [WIDTH*2-1+4:0] tmp04_5_71;
	wire [WIDTH*2-1+4:0] tmp04_5_72;
	wire [WIDTH*2-1+4:0] tmp04_5_73;
	wire [WIDTH*2-1+4:0] tmp04_5_74;
	wire [WIDTH*2-1+4:0] tmp04_5_75;
	wire [WIDTH*2-1+4:0] tmp04_5_76;
	wire [WIDTH*2-1+4:0] tmp04_5_77;
	wire [WIDTH*2-1+4:0] tmp04_5_78;
	wire [WIDTH*2-1+4:0] tmp04_5_79;
	wire [WIDTH*2-1+4:0] tmp04_5_80;
	wire [WIDTH*2-1+4:0] tmp04_5_81;
	wire [WIDTH*2-1+4:0] tmp04_5_82;
	wire [WIDTH*2-1+4:0] tmp04_5_83;
	wire [WIDTH*2-1+4:0] tmp04_6_0;
	wire [WIDTH*2-1+4:0] tmp04_6_1;
	wire [WIDTH*2-1+4:0] tmp04_6_2;
	wire [WIDTH*2-1+4:0] tmp04_6_3;
	wire [WIDTH*2-1+4:0] tmp04_6_4;
	wire [WIDTH*2-1+4:0] tmp04_6_5;
	wire [WIDTH*2-1+4:0] tmp04_6_6;
	wire [WIDTH*2-1+4:0] tmp04_6_7;
	wire [WIDTH*2-1+4:0] tmp04_6_8;
	wire [WIDTH*2-1+4:0] tmp04_6_9;
	wire [WIDTH*2-1+4:0] tmp04_6_10;
	wire [WIDTH*2-1+4:0] tmp04_6_11;
	wire [WIDTH*2-1+4:0] tmp04_6_12;
	wire [WIDTH*2-1+4:0] tmp04_6_13;
	wire [WIDTH*2-1+4:0] tmp04_6_14;
	wire [WIDTH*2-1+4:0] tmp04_6_15;
	wire [WIDTH*2-1+4:0] tmp04_6_16;
	wire [WIDTH*2-1+4:0] tmp04_6_17;
	wire [WIDTH*2-1+4:0] tmp04_6_18;
	wire [WIDTH*2-1+4:0] tmp04_6_19;
	wire [WIDTH*2-1+4:0] tmp04_6_20;
	wire [WIDTH*2-1+4:0] tmp04_6_21;
	wire [WIDTH*2-1+4:0] tmp04_6_22;
	wire [WIDTH*2-1+4:0] tmp04_6_23;
	wire [WIDTH*2-1+4:0] tmp04_6_24;
	wire [WIDTH*2-1+4:0] tmp04_6_25;
	wire [WIDTH*2-1+4:0] tmp04_6_26;
	wire [WIDTH*2-1+4:0] tmp04_6_27;
	wire [WIDTH*2-1+4:0] tmp04_6_28;
	wire [WIDTH*2-1+4:0] tmp04_6_29;
	wire [WIDTH*2-1+4:0] tmp04_6_30;
	wire [WIDTH*2-1+4:0] tmp04_6_31;
	wire [WIDTH*2-1+4:0] tmp04_6_32;
	wire [WIDTH*2-1+4:0] tmp04_6_33;
	wire [WIDTH*2-1+4:0] tmp04_6_34;
	wire [WIDTH*2-1+4:0] tmp04_6_35;
	wire [WIDTH*2-1+4:0] tmp04_6_36;
	wire [WIDTH*2-1+4:0] tmp04_6_37;
	wire [WIDTH*2-1+4:0] tmp04_6_38;
	wire [WIDTH*2-1+4:0] tmp04_6_39;
	wire [WIDTH*2-1+4:0] tmp04_6_40;
	wire [WIDTH*2-1+4:0] tmp04_6_41;
	wire [WIDTH*2-1+4:0] tmp04_6_42;
	wire [WIDTH*2-1+4:0] tmp04_6_43;
	wire [WIDTH*2-1+4:0] tmp04_6_44;
	wire [WIDTH*2-1+4:0] tmp04_6_45;
	wire [WIDTH*2-1+4:0] tmp04_6_46;
	wire [WIDTH*2-1+4:0] tmp04_6_47;
	wire [WIDTH*2-1+4:0] tmp04_6_48;
	wire [WIDTH*2-1+4:0] tmp04_6_49;
	wire [WIDTH*2-1+4:0] tmp04_6_50;
	wire [WIDTH*2-1+4:0] tmp04_6_51;
	wire [WIDTH*2-1+4:0] tmp04_6_52;
	wire [WIDTH*2-1+4:0] tmp04_6_53;
	wire [WIDTH*2-1+4:0] tmp04_6_54;
	wire [WIDTH*2-1+4:0] tmp04_6_55;
	wire [WIDTH*2-1+4:0] tmp04_6_56;
	wire [WIDTH*2-1+4:0] tmp04_6_57;
	wire [WIDTH*2-1+4:0] tmp04_6_58;
	wire [WIDTH*2-1+4:0] tmp04_6_59;
	wire [WIDTH*2-1+4:0] tmp04_6_60;
	wire [WIDTH*2-1+4:0] tmp04_6_61;
	wire [WIDTH*2-1+4:0] tmp04_6_62;
	wire [WIDTH*2-1+4:0] tmp04_6_63;
	wire [WIDTH*2-1+4:0] tmp04_6_64;
	wire [WIDTH*2-1+4:0] tmp04_6_65;
	wire [WIDTH*2-1+4:0] tmp04_6_66;
	wire [WIDTH*2-1+4:0] tmp04_6_67;
	wire [WIDTH*2-1+4:0] tmp04_6_68;
	wire [WIDTH*2-1+4:0] tmp04_6_69;
	wire [WIDTH*2-1+4:0] tmp04_6_70;
	wire [WIDTH*2-1+4:0] tmp04_6_71;
	wire [WIDTH*2-1+4:0] tmp04_6_72;
	wire [WIDTH*2-1+4:0] tmp04_6_73;
	wire [WIDTH*2-1+4:0] tmp04_6_74;
	wire [WIDTH*2-1+4:0] tmp04_6_75;
	wire [WIDTH*2-1+4:0] tmp04_6_76;
	wire [WIDTH*2-1+4:0] tmp04_6_77;
	wire [WIDTH*2-1+4:0] tmp04_6_78;
	wire [WIDTH*2-1+4:0] tmp04_6_79;
	wire [WIDTH*2-1+4:0] tmp04_6_80;
	wire [WIDTH*2-1+4:0] tmp04_6_81;
	wire [WIDTH*2-1+4:0] tmp04_6_82;
	wire [WIDTH*2-1+4:0] tmp04_6_83;
	wire [WIDTH*2-1+4:0] tmp04_7_0;
	wire [WIDTH*2-1+4:0] tmp04_7_1;
	wire [WIDTH*2-1+4:0] tmp04_7_2;
	wire [WIDTH*2-1+4:0] tmp04_7_3;
	wire [WIDTH*2-1+4:0] tmp04_7_4;
	wire [WIDTH*2-1+4:0] tmp04_7_5;
	wire [WIDTH*2-1+4:0] tmp04_7_6;
	wire [WIDTH*2-1+4:0] tmp04_7_7;
	wire [WIDTH*2-1+4:0] tmp04_7_8;
	wire [WIDTH*2-1+4:0] tmp04_7_9;
	wire [WIDTH*2-1+4:0] tmp04_7_10;
	wire [WIDTH*2-1+4:0] tmp04_7_11;
	wire [WIDTH*2-1+4:0] tmp04_7_12;
	wire [WIDTH*2-1+4:0] tmp04_7_13;
	wire [WIDTH*2-1+4:0] tmp04_7_14;
	wire [WIDTH*2-1+4:0] tmp04_7_15;
	wire [WIDTH*2-1+4:0] tmp04_7_16;
	wire [WIDTH*2-1+4:0] tmp04_7_17;
	wire [WIDTH*2-1+4:0] tmp04_7_18;
	wire [WIDTH*2-1+4:0] tmp04_7_19;
	wire [WIDTH*2-1+4:0] tmp04_7_20;
	wire [WIDTH*2-1+4:0] tmp04_7_21;
	wire [WIDTH*2-1+4:0] tmp04_7_22;
	wire [WIDTH*2-1+4:0] tmp04_7_23;
	wire [WIDTH*2-1+4:0] tmp04_7_24;
	wire [WIDTH*2-1+4:0] tmp04_7_25;
	wire [WIDTH*2-1+4:0] tmp04_7_26;
	wire [WIDTH*2-1+4:0] tmp04_7_27;
	wire [WIDTH*2-1+4:0] tmp04_7_28;
	wire [WIDTH*2-1+4:0] tmp04_7_29;
	wire [WIDTH*2-1+4:0] tmp04_7_30;
	wire [WIDTH*2-1+4:0] tmp04_7_31;
	wire [WIDTH*2-1+4:0] tmp04_7_32;
	wire [WIDTH*2-1+4:0] tmp04_7_33;
	wire [WIDTH*2-1+4:0] tmp04_7_34;
	wire [WIDTH*2-1+4:0] tmp04_7_35;
	wire [WIDTH*2-1+4:0] tmp04_7_36;
	wire [WIDTH*2-1+4:0] tmp04_7_37;
	wire [WIDTH*2-1+4:0] tmp04_7_38;
	wire [WIDTH*2-1+4:0] tmp04_7_39;
	wire [WIDTH*2-1+4:0] tmp04_7_40;
	wire [WIDTH*2-1+4:0] tmp04_7_41;
	wire [WIDTH*2-1+4:0] tmp04_7_42;
	wire [WIDTH*2-1+4:0] tmp04_7_43;
	wire [WIDTH*2-1+4:0] tmp04_7_44;
	wire [WIDTH*2-1+4:0] tmp04_7_45;
	wire [WIDTH*2-1+4:0] tmp04_7_46;
	wire [WIDTH*2-1+4:0] tmp04_7_47;
	wire [WIDTH*2-1+4:0] tmp04_7_48;
	wire [WIDTH*2-1+4:0] tmp04_7_49;
	wire [WIDTH*2-1+4:0] tmp04_7_50;
	wire [WIDTH*2-1+4:0] tmp04_7_51;
	wire [WIDTH*2-1+4:0] tmp04_7_52;
	wire [WIDTH*2-1+4:0] tmp04_7_53;
	wire [WIDTH*2-1+4:0] tmp04_7_54;
	wire [WIDTH*2-1+4:0] tmp04_7_55;
	wire [WIDTH*2-1+4:0] tmp04_7_56;
	wire [WIDTH*2-1+4:0] tmp04_7_57;
	wire [WIDTH*2-1+4:0] tmp04_7_58;
	wire [WIDTH*2-1+4:0] tmp04_7_59;
	wire [WIDTH*2-1+4:0] tmp04_7_60;
	wire [WIDTH*2-1+4:0] tmp04_7_61;
	wire [WIDTH*2-1+4:0] tmp04_7_62;
	wire [WIDTH*2-1+4:0] tmp04_7_63;
	wire [WIDTH*2-1+4:0] tmp04_7_64;
	wire [WIDTH*2-1+4:0] tmp04_7_65;
	wire [WIDTH*2-1+4:0] tmp04_7_66;
	wire [WIDTH*2-1+4:0] tmp04_7_67;
	wire [WIDTH*2-1+4:0] tmp04_7_68;
	wire [WIDTH*2-1+4:0] tmp04_7_69;
	wire [WIDTH*2-1+4:0] tmp04_7_70;
	wire [WIDTH*2-1+4:0] tmp04_7_71;
	wire [WIDTH*2-1+4:0] tmp04_7_72;
	wire [WIDTH*2-1+4:0] tmp04_7_73;
	wire [WIDTH*2-1+4:0] tmp04_7_74;
	wire [WIDTH*2-1+4:0] tmp04_7_75;
	wire [WIDTH*2-1+4:0] tmp04_7_76;
	wire [WIDTH*2-1+4:0] tmp04_7_77;
	wire [WIDTH*2-1+4:0] tmp04_7_78;
	wire [WIDTH*2-1+4:0] tmp04_7_79;
	wire [WIDTH*2-1+4:0] tmp04_7_80;
	wire [WIDTH*2-1+4:0] tmp04_7_81;
	wire [WIDTH*2-1+4:0] tmp04_7_82;
	wire [WIDTH*2-1+4:0] tmp04_7_83;
	wire [WIDTH*2-1+5:0] tmp05_0_0;
	wire [WIDTH*2-1+5:0] tmp05_0_1;
	wire [WIDTH*2-1+5:0] tmp05_0_2;
	wire [WIDTH*2-1+5:0] tmp05_0_3;
	wire [WIDTH*2-1+5:0] tmp05_0_4;
	wire [WIDTH*2-1+5:0] tmp05_0_5;
	wire [WIDTH*2-1+5:0] tmp05_0_6;
	wire [WIDTH*2-1+5:0] tmp05_0_7;
	wire [WIDTH*2-1+5:0] tmp05_0_8;
	wire [WIDTH*2-1+5:0] tmp05_0_9;
	wire [WIDTH*2-1+5:0] tmp05_0_10;
	wire [WIDTH*2-1+5:0] tmp05_0_11;
	wire [WIDTH*2-1+5:0] tmp05_0_12;
	wire [WIDTH*2-1+5:0] tmp05_0_13;
	wire [WIDTH*2-1+5:0] tmp05_0_14;
	wire [WIDTH*2-1+5:0] tmp05_0_15;
	wire [WIDTH*2-1+5:0] tmp05_0_16;
	wire [WIDTH*2-1+5:0] tmp05_0_17;
	wire [WIDTH*2-1+5:0] tmp05_0_18;
	wire [WIDTH*2-1+5:0] tmp05_0_19;
	wire [WIDTH*2-1+5:0] tmp05_0_20;
	wire [WIDTH*2-1+5:0] tmp05_0_21;
	wire [WIDTH*2-1+5:0] tmp05_0_22;
	wire [WIDTH*2-1+5:0] tmp05_0_23;
	wire [WIDTH*2-1+5:0] tmp05_0_24;
	wire [WIDTH*2-1+5:0] tmp05_0_25;
	wire [WIDTH*2-1+5:0] tmp05_0_26;
	wire [WIDTH*2-1+5:0] tmp05_0_27;
	wire [WIDTH*2-1+5:0] tmp05_0_28;
	wire [WIDTH*2-1+5:0] tmp05_0_29;
	wire [WIDTH*2-1+5:0] tmp05_0_30;
	wire [WIDTH*2-1+5:0] tmp05_0_31;
	wire [WIDTH*2-1+5:0] tmp05_0_32;
	wire [WIDTH*2-1+5:0] tmp05_0_33;
	wire [WIDTH*2-1+5:0] tmp05_0_34;
	wire [WIDTH*2-1+5:0] tmp05_0_35;
	wire [WIDTH*2-1+5:0] tmp05_0_36;
	wire [WIDTH*2-1+5:0] tmp05_0_37;
	wire [WIDTH*2-1+5:0] tmp05_0_38;
	wire [WIDTH*2-1+5:0] tmp05_0_39;
	wire [WIDTH*2-1+5:0] tmp05_0_40;
	wire [WIDTH*2-1+5:0] tmp05_0_41;
	wire [WIDTH*2-1+5:0] tmp05_0_42;
	wire [WIDTH*2-1+5:0] tmp05_0_43;
	wire [WIDTH*2-1+5:0] tmp05_0_44;
	wire [WIDTH*2-1+5:0] tmp05_0_45;
	wire [WIDTH*2-1+5:0] tmp05_0_46;
	wire [WIDTH*2-1+5:0] tmp05_0_47;
	wire [WIDTH*2-1+5:0] tmp05_0_48;
	wire [WIDTH*2-1+5:0] tmp05_0_49;
	wire [WIDTH*2-1+5:0] tmp05_0_50;
	wire [WIDTH*2-1+5:0] tmp05_0_51;
	wire [WIDTH*2-1+5:0] tmp05_0_52;
	wire [WIDTH*2-1+5:0] tmp05_0_53;
	wire [WIDTH*2-1+5:0] tmp05_0_54;
	wire [WIDTH*2-1+5:0] tmp05_0_55;
	wire [WIDTH*2-1+5:0] tmp05_0_56;
	wire [WIDTH*2-1+5:0] tmp05_0_57;
	wire [WIDTH*2-1+5:0] tmp05_0_58;
	wire [WIDTH*2-1+5:0] tmp05_0_59;
	wire [WIDTH*2-1+5:0] tmp05_0_60;
	wire [WIDTH*2-1+5:0] tmp05_0_61;
	wire [WIDTH*2-1+5:0] tmp05_0_62;
	wire [WIDTH*2-1+5:0] tmp05_0_63;
	wire [WIDTH*2-1+5:0] tmp05_0_64;
	wire [WIDTH*2-1+5:0] tmp05_0_65;
	wire [WIDTH*2-1+5:0] tmp05_0_66;
	wire [WIDTH*2-1+5:0] tmp05_0_67;
	wire [WIDTH*2-1+5:0] tmp05_0_68;
	wire [WIDTH*2-1+5:0] tmp05_0_69;
	wire [WIDTH*2-1+5:0] tmp05_0_70;
	wire [WIDTH*2-1+5:0] tmp05_0_71;
	wire [WIDTH*2-1+5:0] tmp05_0_72;
	wire [WIDTH*2-1+5:0] tmp05_0_73;
	wire [WIDTH*2-1+5:0] tmp05_0_74;
	wire [WIDTH*2-1+5:0] tmp05_0_75;
	wire [WIDTH*2-1+5:0] tmp05_0_76;
	wire [WIDTH*2-1+5:0] tmp05_0_77;
	wire [WIDTH*2-1+5:0] tmp05_0_78;
	wire [WIDTH*2-1+5:0] tmp05_0_79;
	wire [WIDTH*2-1+5:0] tmp05_0_80;
	wire [WIDTH*2-1+5:0] tmp05_0_81;
	wire [WIDTH*2-1+5:0] tmp05_0_82;
	wire [WIDTH*2-1+5:0] tmp05_0_83;
	wire [WIDTH*2-1+5:0] tmp05_1_0;
	wire [WIDTH*2-1+5:0] tmp05_1_1;
	wire [WIDTH*2-1+5:0] tmp05_1_2;
	wire [WIDTH*2-1+5:0] tmp05_1_3;
	wire [WIDTH*2-1+5:0] tmp05_1_4;
	wire [WIDTH*2-1+5:0] tmp05_1_5;
	wire [WIDTH*2-1+5:0] tmp05_1_6;
	wire [WIDTH*2-1+5:0] tmp05_1_7;
	wire [WIDTH*2-1+5:0] tmp05_1_8;
	wire [WIDTH*2-1+5:0] tmp05_1_9;
	wire [WIDTH*2-1+5:0] tmp05_1_10;
	wire [WIDTH*2-1+5:0] tmp05_1_11;
	wire [WIDTH*2-1+5:0] tmp05_1_12;
	wire [WIDTH*2-1+5:0] tmp05_1_13;
	wire [WIDTH*2-1+5:0] tmp05_1_14;
	wire [WIDTH*2-1+5:0] tmp05_1_15;
	wire [WIDTH*2-1+5:0] tmp05_1_16;
	wire [WIDTH*2-1+5:0] tmp05_1_17;
	wire [WIDTH*2-1+5:0] tmp05_1_18;
	wire [WIDTH*2-1+5:0] tmp05_1_19;
	wire [WIDTH*2-1+5:0] tmp05_1_20;
	wire [WIDTH*2-1+5:0] tmp05_1_21;
	wire [WIDTH*2-1+5:0] tmp05_1_22;
	wire [WIDTH*2-1+5:0] tmp05_1_23;
	wire [WIDTH*2-1+5:0] tmp05_1_24;
	wire [WIDTH*2-1+5:0] tmp05_1_25;
	wire [WIDTH*2-1+5:0] tmp05_1_26;
	wire [WIDTH*2-1+5:0] tmp05_1_27;
	wire [WIDTH*2-1+5:0] tmp05_1_28;
	wire [WIDTH*2-1+5:0] tmp05_1_29;
	wire [WIDTH*2-1+5:0] tmp05_1_30;
	wire [WIDTH*2-1+5:0] tmp05_1_31;
	wire [WIDTH*2-1+5:0] tmp05_1_32;
	wire [WIDTH*2-1+5:0] tmp05_1_33;
	wire [WIDTH*2-1+5:0] tmp05_1_34;
	wire [WIDTH*2-1+5:0] tmp05_1_35;
	wire [WIDTH*2-1+5:0] tmp05_1_36;
	wire [WIDTH*2-1+5:0] tmp05_1_37;
	wire [WIDTH*2-1+5:0] tmp05_1_38;
	wire [WIDTH*2-1+5:0] tmp05_1_39;
	wire [WIDTH*2-1+5:0] tmp05_1_40;
	wire [WIDTH*2-1+5:0] tmp05_1_41;
	wire [WIDTH*2-1+5:0] tmp05_1_42;
	wire [WIDTH*2-1+5:0] tmp05_1_43;
	wire [WIDTH*2-1+5:0] tmp05_1_44;
	wire [WIDTH*2-1+5:0] tmp05_1_45;
	wire [WIDTH*2-1+5:0] tmp05_1_46;
	wire [WIDTH*2-1+5:0] tmp05_1_47;
	wire [WIDTH*2-1+5:0] tmp05_1_48;
	wire [WIDTH*2-1+5:0] tmp05_1_49;
	wire [WIDTH*2-1+5:0] tmp05_1_50;
	wire [WIDTH*2-1+5:0] tmp05_1_51;
	wire [WIDTH*2-1+5:0] tmp05_1_52;
	wire [WIDTH*2-1+5:0] tmp05_1_53;
	wire [WIDTH*2-1+5:0] tmp05_1_54;
	wire [WIDTH*2-1+5:0] tmp05_1_55;
	wire [WIDTH*2-1+5:0] tmp05_1_56;
	wire [WIDTH*2-1+5:0] tmp05_1_57;
	wire [WIDTH*2-1+5:0] tmp05_1_58;
	wire [WIDTH*2-1+5:0] tmp05_1_59;
	wire [WIDTH*2-1+5:0] tmp05_1_60;
	wire [WIDTH*2-1+5:0] tmp05_1_61;
	wire [WIDTH*2-1+5:0] tmp05_1_62;
	wire [WIDTH*2-1+5:0] tmp05_1_63;
	wire [WIDTH*2-1+5:0] tmp05_1_64;
	wire [WIDTH*2-1+5:0] tmp05_1_65;
	wire [WIDTH*2-1+5:0] tmp05_1_66;
	wire [WIDTH*2-1+5:0] tmp05_1_67;
	wire [WIDTH*2-1+5:0] tmp05_1_68;
	wire [WIDTH*2-1+5:0] tmp05_1_69;
	wire [WIDTH*2-1+5:0] tmp05_1_70;
	wire [WIDTH*2-1+5:0] tmp05_1_71;
	wire [WIDTH*2-1+5:0] tmp05_1_72;
	wire [WIDTH*2-1+5:0] tmp05_1_73;
	wire [WIDTH*2-1+5:0] tmp05_1_74;
	wire [WIDTH*2-1+5:0] tmp05_1_75;
	wire [WIDTH*2-1+5:0] tmp05_1_76;
	wire [WIDTH*2-1+5:0] tmp05_1_77;
	wire [WIDTH*2-1+5:0] tmp05_1_78;
	wire [WIDTH*2-1+5:0] tmp05_1_79;
	wire [WIDTH*2-1+5:0] tmp05_1_80;
	wire [WIDTH*2-1+5:0] tmp05_1_81;
	wire [WIDTH*2-1+5:0] tmp05_1_82;
	wire [WIDTH*2-1+5:0] tmp05_1_83;
	wire [WIDTH*2-1+5:0] tmp05_2_0;
	wire [WIDTH*2-1+5:0] tmp05_2_1;
	wire [WIDTH*2-1+5:0] tmp05_2_2;
	wire [WIDTH*2-1+5:0] tmp05_2_3;
	wire [WIDTH*2-1+5:0] tmp05_2_4;
	wire [WIDTH*2-1+5:0] tmp05_2_5;
	wire [WIDTH*2-1+5:0] tmp05_2_6;
	wire [WIDTH*2-1+5:0] tmp05_2_7;
	wire [WIDTH*2-1+5:0] tmp05_2_8;
	wire [WIDTH*2-1+5:0] tmp05_2_9;
	wire [WIDTH*2-1+5:0] tmp05_2_10;
	wire [WIDTH*2-1+5:0] tmp05_2_11;
	wire [WIDTH*2-1+5:0] tmp05_2_12;
	wire [WIDTH*2-1+5:0] tmp05_2_13;
	wire [WIDTH*2-1+5:0] tmp05_2_14;
	wire [WIDTH*2-1+5:0] tmp05_2_15;
	wire [WIDTH*2-1+5:0] tmp05_2_16;
	wire [WIDTH*2-1+5:0] tmp05_2_17;
	wire [WIDTH*2-1+5:0] tmp05_2_18;
	wire [WIDTH*2-1+5:0] tmp05_2_19;
	wire [WIDTH*2-1+5:0] tmp05_2_20;
	wire [WIDTH*2-1+5:0] tmp05_2_21;
	wire [WIDTH*2-1+5:0] tmp05_2_22;
	wire [WIDTH*2-1+5:0] tmp05_2_23;
	wire [WIDTH*2-1+5:0] tmp05_2_24;
	wire [WIDTH*2-1+5:0] tmp05_2_25;
	wire [WIDTH*2-1+5:0] tmp05_2_26;
	wire [WIDTH*2-1+5:0] tmp05_2_27;
	wire [WIDTH*2-1+5:0] tmp05_2_28;
	wire [WIDTH*2-1+5:0] tmp05_2_29;
	wire [WIDTH*2-1+5:0] tmp05_2_30;
	wire [WIDTH*2-1+5:0] tmp05_2_31;
	wire [WIDTH*2-1+5:0] tmp05_2_32;
	wire [WIDTH*2-1+5:0] tmp05_2_33;
	wire [WIDTH*2-1+5:0] tmp05_2_34;
	wire [WIDTH*2-1+5:0] tmp05_2_35;
	wire [WIDTH*2-1+5:0] tmp05_2_36;
	wire [WIDTH*2-1+5:0] tmp05_2_37;
	wire [WIDTH*2-1+5:0] tmp05_2_38;
	wire [WIDTH*2-1+5:0] tmp05_2_39;
	wire [WIDTH*2-1+5:0] tmp05_2_40;
	wire [WIDTH*2-1+5:0] tmp05_2_41;
	wire [WIDTH*2-1+5:0] tmp05_2_42;
	wire [WIDTH*2-1+5:0] tmp05_2_43;
	wire [WIDTH*2-1+5:0] tmp05_2_44;
	wire [WIDTH*2-1+5:0] tmp05_2_45;
	wire [WIDTH*2-1+5:0] tmp05_2_46;
	wire [WIDTH*2-1+5:0] tmp05_2_47;
	wire [WIDTH*2-1+5:0] tmp05_2_48;
	wire [WIDTH*2-1+5:0] tmp05_2_49;
	wire [WIDTH*2-1+5:0] tmp05_2_50;
	wire [WIDTH*2-1+5:0] tmp05_2_51;
	wire [WIDTH*2-1+5:0] tmp05_2_52;
	wire [WIDTH*2-1+5:0] tmp05_2_53;
	wire [WIDTH*2-1+5:0] tmp05_2_54;
	wire [WIDTH*2-1+5:0] tmp05_2_55;
	wire [WIDTH*2-1+5:0] tmp05_2_56;
	wire [WIDTH*2-1+5:0] tmp05_2_57;
	wire [WIDTH*2-1+5:0] tmp05_2_58;
	wire [WIDTH*2-1+5:0] tmp05_2_59;
	wire [WIDTH*2-1+5:0] tmp05_2_60;
	wire [WIDTH*2-1+5:0] tmp05_2_61;
	wire [WIDTH*2-1+5:0] tmp05_2_62;
	wire [WIDTH*2-1+5:0] tmp05_2_63;
	wire [WIDTH*2-1+5:0] tmp05_2_64;
	wire [WIDTH*2-1+5:0] tmp05_2_65;
	wire [WIDTH*2-1+5:0] tmp05_2_66;
	wire [WIDTH*2-1+5:0] tmp05_2_67;
	wire [WIDTH*2-1+5:0] tmp05_2_68;
	wire [WIDTH*2-1+5:0] tmp05_2_69;
	wire [WIDTH*2-1+5:0] tmp05_2_70;
	wire [WIDTH*2-1+5:0] tmp05_2_71;
	wire [WIDTH*2-1+5:0] tmp05_2_72;
	wire [WIDTH*2-1+5:0] tmp05_2_73;
	wire [WIDTH*2-1+5:0] tmp05_2_74;
	wire [WIDTH*2-1+5:0] tmp05_2_75;
	wire [WIDTH*2-1+5:0] tmp05_2_76;
	wire [WIDTH*2-1+5:0] tmp05_2_77;
	wire [WIDTH*2-1+5:0] tmp05_2_78;
	wire [WIDTH*2-1+5:0] tmp05_2_79;
	wire [WIDTH*2-1+5:0] tmp05_2_80;
	wire [WIDTH*2-1+5:0] tmp05_2_81;
	wire [WIDTH*2-1+5:0] tmp05_2_82;
	wire [WIDTH*2-1+5:0] tmp05_2_83;
	wire [WIDTH*2-1+5:0] tmp05_3_0;
	wire [WIDTH*2-1+5:0] tmp05_3_1;
	wire [WIDTH*2-1+5:0] tmp05_3_2;
	wire [WIDTH*2-1+5:0] tmp05_3_3;
	wire [WIDTH*2-1+5:0] tmp05_3_4;
	wire [WIDTH*2-1+5:0] tmp05_3_5;
	wire [WIDTH*2-1+5:0] tmp05_3_6;
	wire [WIDTH*2-1+5:0] tmp05_3_7;
	wire [WIDTH*2-1+5:0] tmp05_3_8;
	wire [WIDTH*2-1+5:0] tmp05_3_9;
	wire [WIDTH*2-1+5:0] tmp05_3_10;
	wire [WIDTH*2-1+5:0] tmp05_3_11;
	wire [WIDTH*2-1+5:0] tmp05_3_12;
	wire [WIDTH*2-1+5:0] tmp05_3_13;
	wire [WIDTH*2-1+5:0] tmp05_3_14;
	wire [WIDTH*2-1+5:0] tmp05_3_15;
	wire [WIDTH*2-1+5:0] tmp05_3_16;
	wire [WIDTH*2-1+5:0] tmp05_3_17;
	wire [WIDTH*2-1+5:0] tmp05_3_18;
	wire [WIDTH*2-1+5:0] tmp05_3_19;
	wire [WIDTH*2-1+5:0] tmp05_3_20;
	wire [WIDTH*2-1+5:0] tmp05_3_21;
	wire [WIDTH*2-1+5:0] tmp05_3_22;
	wire [WIDTH*2-1+5:0] tmp05_3_23;
	wire [WIDTH*2-1+5:0] tmp05_3_24;
	wire [WIDTH*2-1+5:0] tmp05_3_25;
	wire [WIDTH*2-1+5:0] tmp05_3_26;
	wire [WIDTH*2-1+5:0] tmp05_3_27;
	wire [WIDTH*2-1+5:0] tmp05_3_28;
	wire [WIDTH*2-1+5:0] tmp05_3_29;
	wire [WIDTH*2-1+5:0] tmp05_3_30;
	wire [WIDTH*2-1+5:0] tmp05_3_31;
	wire [WIDTH*2-1+5:0] tmp05_3_32;
	wire [WIDTH*2-1+5:0] tmp05_3_33;
	wire [WIDTH*2-1+5:0] tmp05_3_34;
	wire [WIDTH*2-1+5:0] tmp05_3_35;
	wire [WIDTH*2-1+5:0] tmp05_3_36;
	wire [WIDTH*2-1+5:0] tmp05_3_37;
	wire [WIDTH*2-1+5:0] tmp05_3_38;
	wire [WIDTH*2-1+5:0] tmp05_3_39;
	wire [WIDTH*2-1+5:0] tmp05_3_40;
	wire [WIDTH*2-1+5:0] tmp05_3_41;
	wire [WIDTH*2-1+5:0] tmp05_3_42;
	wire [WIDTH*2-1+5:0] tmp05_3_43;
	wire [WIDTH*2-1+5:0] tmp05_3_44;
	wire [WIDTH*2-1+5:0] tmp05_3_45;
	wire [WIDTH*2-1+5:0] tmp05_3_46;
	wire [WIDTH*2-1+5:0] tmp05_3_47;
	wire [WIDTH*2-1+5:0] tmp05_3_48;
	wire [WIDTH*2-1+5:0] tmp05_3_49;
	wire [WIDTH*2-1+5:0] tmp05_3_50;
	wire [WIDTH*2-1+5:0] tmp05_3_51;
	wire [WIDTH*2-1+5:0] tmp05_3_52;
	wire [WIDTH*2-1+5:0] tmp05_3_53;
	wire [WIDTH*2-1+5:0] tmp05_3_54;
	wire [WIDTH*2-1+5:0] tmp05_3_55;
	wire [WIDTH*2-1+5:0] tmp05_3_56;
	wire [WIDTH*2-1+5:0] tmp05_3_57;
	wire [WIDTH*2-1+5:0] tmp05_3_58;
	wire [WIDTH*2-1+5:0] tmp05_3_59;
	wire [WIDTH*2-1+5:0] tmp05_3_60;
	wire [WIDTH*2-1+5:0] tmp05_3_61;
	wire [WIDTH*2-1+5:0] tmp05_3_62;
	wire [WIDTH*2-1+5:0] tmp05_3_63;
	wire [WIDTH*2-1+5:0] tmp05_3_64;
	wire [WIDTH*2-1+5:0] tmp05_3_65;
	wire [WIDTH*2-1+5:0] tmp05_3_66;
	wire [WIDTH*2-1+5:0] tmp05_3_67;
	wire [WIDTH*2-1+5:0] tmp05_3_68;
	wire [WIDTH*2-1+5:0] tmp05_3_69;
	wire [WIDTH*2-1+5:0] tmp05_3_70;
	wire [WIDTH*2-1+5:0] tmp05_3_71;
	wire [WIDTH*2-1+5:0] tmp05_3_72;
	wire [WIDTH*2-1+5:0] tmp05_3_73;
	wire [WIDTH*2-1+5:0] tmp05_3_74;
	wire [WIDTH*2-1+5:0] tmp05_3_75;
	wire [WIDTH*2-1+5:0] tmp05_3_76;
	wire [WIDTH*2-1+5:0] tmp05_3_77;
	wire [WIDTH*2-1+5:0] tmp05_3_78;
	wire [WIDTH*2-1+5:0] tmp05_3_79;
	wire [WIDTH*2-1+5:0] tmp05_3_80;
	wire [WIDTH*2-1+5:0] tmp05_3_81;
	wire [WIDTH*2-1+5:0] tmp05_3_82;
	wire [WIDTH*2-1+5:0] tmp05_3_83;
	wire [WIDTH*2-1+6:0] tmp06_0_0;
	wire [WIDTH*2-1+6:0] tmp06_0_1;
	wire [WIDTH*2-1+6:0] tmp06_0_2;
	wire [WIDTH*2-1+6:0] tmp06_0_3;
	wire [WIDTH*2-1+6:0] tmp06_0_4;
	wire [WIDTH*2-1+6:0] tmp06_0_5;
	wire [WIDTH*2-1+6:0] tmp06_0_6;
	wire [WIDTH*2-1+6:0] tmp06_0_7;
	wire [WIDTH*2-1+6:0] tmp06_0_8;
	wire [WIDTH*2-1+6:0] tmp06_0_9;
	wire [WIDTH*2-1+6:0] tmp06_0_10;
	wire [WIDTH*2-1+6:0] tmp06_0_11;
	wire [WIDTH*2-1+6:0] tmp06_0_12;
	wire [WIDTH*2-1+6:0] tmp06_0_13;
	wire [WIDTH*2-1+6:0] tmp06_0_14;
	wire [WIDTH*2-1+6:0] tmp06_0_15;
	wire [WIDTH*2-1+6:0] tmp06_0_16;
	wire [WIDTH*2-1+6:0] tmp06_0_17;
	wire [WIDTH*2-1+6:0] tmp06_0_18;
	wire [WIDTH*2-1+6:0] tmp06_0_19;
	wire [WIDTH*2-1+6:0] tmp06_0_20;
	wire [WIDTH*2-1+6:0] tmp06_0_21;
	wire [WIDTH*2-1+6:0] tmp06_0_22;
	wire [WIDTH*2-1+6:0] tmp06_0_23;
	wire [WIDTH*2-1+6:0] tmp06_0_24;
	wire [WIDTH*2-1+6:0] tmp06_0_25;
	wire [WIDTH*2-1+6:0] tmp06_0_26;
	wire [WIDTH*2-1+6:0] tmp06_0_27;
	wire [WIDTH*2-1+6:0] tmp06_0_28;
	wire [WIDTH*2-1+6:0] tmp06_0_29;
	wire [WIDTH*2-1+6:0] tmp06_0_30;
	wire [WIDTH*2-1+6:0] tmp06_0_31;
	wire [WIDTH*2-1+6:0] tmp06_0_32;
	wire [WIDTH*2-1+6:0] tmp06_0_33;
	wire [WIDTH*2-1+6:0] tmp06_0_34;
	wire [WIDTH*2-1+6:0] tmp06_0_35;
	wire [WIDTH*2-1+6:0] tmp06_0_36;
	wire [WIDTH*2-1+6:0] tmp06_0_37;
	wire [WIDTH*2-1+6:0] tmp06_0_38;
	wire [WIDTH*2-1+6:0] tmp06_0_39;
	wire [WIDTH*2-1+6:0] tmp06_0_40;
	wire [WIDTH*2-1+6:0] tmp06_0_41;
	wire [WIDTH*2-1+6:0] tmp06_0_42;
	wire [WIDTH*2-1+6:0] tmp06_0_43;
	wire [WIDTH*2-1+6:0] tmp06_0_44;
	wire [WIDTH*2-1+6:0] tmp06_0_45;
	wire [WIDTH*2-1+6:0] tmp06_0_46;
	wire [WIDTH*2-1+6:0] tmp06_0_47;
	wire [WIDTH*2-1+6:0] tmp06_0_48;
	wire [WIDTH*2-1+6:0] tmp06_0_49;
	wire [WIDTH*2-1+6:0] tmp06_0_50;
	wire [WIDTH*2-1+6:0] tmp06_0_51;
	wire [WIDTH*2-1+6:0] tmp06_0_52;
	wire [WIDTH*2-1+6:0] tmp06_0_53;
	wire [WIDTH*2-1+6:0] tmp06_0_54;
	wire [WIDTH*2-1+6:0] tmp06_0_55;
	wire [WIDTH*2-1+6:0] tmp06_0_56;
	wire [WIDTH*2-1+6:0] tmp06_0_57;
	wire [WIDTH*2-1+6:0] tmp06_0_58;
	wire [WIDTH*2-1+6:0] tmp06_0_59;
	wire [WIDTH*2-1+6:0] tmp06_0_60;
	wire [WIDTH*2-1+6:0] tmp06_0_61;
	wire [WIDTH*2-1+6:0] tmp06_0_62;
	wire [WIDTH*2-1+6:0] tmp06_0_63;
	wire [WIDTH*2-1+6:0] tmp06_0_64;
	wire [WIDTH*2-1+6:0] tmp06_0_65;
	wire [WIDTH*2-1+6:0] tmp06_0_66;
	wire [WIDTH*2-1+6:0] tmp06_0_67;
	wire [WIDTH*2-1+6:0] tmp06_0_68;
	wire [WIDTH*2-1+6:0] tmp06_0_69;
	wire [WIDTH*2-1+6:0] tmp06_0_70;
	wire [WIDTH*2-1+6:0] tmp06_0_71;
	wire [WIDTH*2-1+6:0] tmp06_0_72;
	wire [WIDTH*2-1+6:0] tmp06_0_73;
	wire [WIDTH*2-1+6:0] tmp06_0_74;
	wire [WIDTH*2-1+6:0] tmp06_0_75;
	wire [WIDTH*2-1+6:0] tmp06_0_76;
	wire [WIDTH*2-1+6:0] tmp06_0_77;
	wire [WIDTH*2-1+6:0] tmp06_0_78;
	wire [WIDTH*2-1+6:0] tmp06_0_79;
	wire [WIDTH*2-1+6:0] tmp06_0_80;
	wire [WIDTH*2-1+6:0] tmp06_0_81;
	wire [WIDTH*2-1+6:0] tmp06_0_82;
	wire [WIDTH*2-1+6:0] tmp06_0_83;
	wire [WIDTH*2-1+6:0] tmp06_1_0;
	wire [WIDTH*2-1+6:0] tmp06_1_1;
	wire [WIDTH*2-1+6:0] tmp06_1_2;
	wire [WIDTH*2-1+6:0] tmp06_1_3;
	wire [WIDTH*2-1+6:0] tmp06_1_4;
	wire [WIDTH*2-1+6:0] tmp06_1_5;
	wire [WIDTH*2-1+6:0] tmp06_1_6;
	wire [WIDTH*2-1+6:0] tmp06_1_7;
	wire [WIDTH*2-1+6:0] tmp06_1_8;
	wire [WIDTH*2-1+6:0] tmp06_1_9;
	wire [WIDTH*2-1+6:0] tmp06_1_10;
	wire [WIDTH*2-1+6:0] tmp06_1_11;
	wire [WIDTH*2-1+6:0] tmp06_1_12;
	wire [WIDTH*2-1+6:0] tmp06_1_13;
	wire [WIDTH*2-1+6:0] tmp06_1_14;
	wire [WIDTH*2-1+6:0] tmp06_1_15;
	wire [WIDTH*2-1+6:0] tmp06_1_16;
	wire [WIDTH*2-1+6:0] tmp06_1_17;
	wire [WIDTH*2-1+6:0] tmp06_1_18;
	wire [WIDTH*2-1+6:0] tmp06_1_19;
	wire [WIDTH*2-1+6:0] tmp06_1_20;
	wire [WIDTH*2-1+6:0] tmp06_1_21;
	wire [WIDTH*2-1+6:0] tmp06_1_22;
	wire [WIDTH*2-1+6:0] tmp06_1_23;
	wire [WIDTH*2-1+6:0] tmp06_1_24;
	wire [WIDTH*2-1+6:0] tmp06_1_25;
	wire [WIDTH*2-1+6:0] tmp06_1_26;
	wire [WIDTH*2-1+6:0] tmp06_1_27;
	wire [WIDTH*2-1+6:0] tmp06_1_28;
	wire [WIDTH*2-1+6:0] tmp06_1_29;
	wire [WIDTH*2-1+6:0] tmp06_1_30;
	wire [WIDTH*2-1+6:0] tmp06_1_31;
	wire [WIDTH*2-1+6:0] tmp06_1_32;
	wire [WIDTH*2-1+6:0] tmp06_1_33;
	wire [WIDTH*2-1+6:0] tmp06_1_34;
	wire [WIDTH*2-1+6:0] tmp06_1_35;
	wire [WIDTH*2-1+6:0] tmp06_1_36;
	wire [WIDTH*2-1+6:0] tmp06_1_37;
	wire [WIDTH*2-1+6:0] tmp06_1_38;
	wire [WIDTH*2-1+6:0] tmp06_1_39;
	wire [WIDTH*2-1+6:0] tmp06_1_40;
	wire [WIDTH*2-1+6:0] tmp06_1_41;
	wire [WIDTH*2-1+6:0] tmp06_1_42;
	wire [WIDTH*2-1+6:0] tmp06_1_43;
	wire [WIDTH*2-1+6:0] tmp06_1_44;
	wire [WIDTH*2-1+6:0] tmp06_1_45;
	wire [WIDTH*2-1+6:0] tmp06_1_46;
	wire [WIDTH*2-1+6:0] tmp06_1_47;
	wire [WIDTH*2-1+6:0] tmp06_1_48;
	wire [WIDTH*2-1+6:0] tmp06_1_49;
	wire [WIDTH*2-1+6:0] tmp06_1_50;
	wire [WIDTH*2-1+6:0] tmp06_1_51;
	wire [WIDTH*2-1+6:0] tmp06_1_52;
	wire [WIDTH*2-1+6:0] tmp06_1_53;
	wire [WIDTH*2-1+6:0] tmp06_1_54;
	wire [WIDTH*2-1+6:0] tmp06_1_55;
	wire [WIDTH*2-1+6:0] tmp06_1_56;
	wire [WIDTH*2-1+6:0] tmp06_1_57;
	wire [WIDTH*2-1+6:0] tmp06_1_58;
	wire [WIDTH*2-1+6:0] tmp06_1_59;
	wire [WIDTH*2-1+6:0] tmp06_1_60;
	wire [WIDTH*2-1+6:0] tmp06_1_61;
	wire [WIDTH*2-1+6:0] tmp06_1_62;
	wire [WIDTH*2-1+6:0] tmp06_1_63;
	wire [WIDTH*2-1+6:0] tmp06_1_64;
	wire [WIDTH*2-1+6:0] tmp06_1_65;
	wire [WIDTH*2-1+6:0] tmp06_1_66;
	wire [WIDTH*2-1+6:0] tmp06_1_67;
	wire [WIDTH*2-1+6:0] tmp06_1_68;
	wire [WIDTH*2-1+6:0] tmp06_1_69;
	wire [WIDTH*2-1+6:0] tmp06_1_70;
	wire [WIDTH*2-1+6:0] tmp06_1_71;
	wire [WIDTH*2-1+6:0] tmp06_1_72;
	wire [WIDTH*2-1+6:0] tmp06_1_73;
	wire [WIDTH*2-1+6:0] tmp06_1_74;
	wire [WIDTH*2-1+6:0] tmp06_1_75;
	wire [WIDTH*2-1+6:0] tmp06_1_76;
	wire [WIDTH*2-1+6:0] tmp06_1_77;
	wire [WIDTH*2-1+6:0] tmp06_1_78;
	wire [WIDTH*2-1+6:0] tmp06_1_79;
	wire [WIDTH*2-1+6:0] tmp06_1_80;
	wire [WIDTH*2-1+6:0] tmp06_1_81;
	wire [WIDTH*2-1+6:0] tmp06_1_82;
	wire [WIDTH*2-1+6:0] tmp06_1_83;
	wire [WIDTH*2-1+7:0] tmp07_0_0;
	wire [WIDTH*2-1+7:0] tmp07_0_1;
	wire [WIDTH*2-1+7:0] tmp07_0_2;
	wire [WIDTH*2-1+7:0] tmp07_0_3;
	wire [WIDTH*2-1+7:0] tmp07_0_4;
	wire [WIDTH*2-1+7:0] tmp07_0_5;
	wire [WIDTH*2-1+7:0] tmp07_0_6;
	wire [WIDTH*2-1+7:0] tmp07_0_7;
	wire [WIDTH*2-1+7:0] tmp07_0_8;
	wire [WIDTH*2-1+7:0] tmp07_0_9;
	wire [WIDTH*2-1+7:0] tmp07_0_10;
	wire [WIDTH*2-1+7:0] tmp07_0_11;
	wire [WIDTH*2-1+7:0] tmp07_0_12;
	wire [WIDTH*2-1+7:0] tmp07_0_13;
	wire [WIDTH*2-1+7:0] tmp07_0_14;
	wire [WIDTH*2-1+7:0] tmp07_0_15;
	wire [WIDTH*2-1+7:0] tmp07_0_16;
	wire [WIDTH*2-1+7:0] tmp07_0_17;
	wire [WIDTH*2-1+7:0] tmp07_0_18;
	wire [WIDTH*2-1+7:0] tmp07_0_19;
	wire [WIDTH*2-1+7:0] tmp07_0_20;
	wire [WIDTH*2-1+7:0] tmp07_0_21;
	wire [WIDTH*2-1+7:0] tmp07_0_22;
	wire [WIDTH*2-1+7:0] tmp07_0_23;
	wire [WIDTH*2-1+7:0] tmp07_0_24;
	wire [WIDTH*2-1+7:0] tmp07_0_25;
	wire [WIDTH*2-1+7:0] tmp07_0_26;
	wire [WIDTH*2-1+7:0] tmp07_0_27;
	wire [WIDTH*2-1+7:0] tmp07_0_28;
	wire [WIDTH*2-1+7:0] tmp07_0_29;
	wire [WIDTH*2-1+7:0] tmp07_0_30;
	wire [WIDTH*2-1+7:0] tmp07_0_31;
	wire [WIDTH*2-1+7:0] tmp07_0_32;
	wire [WIDTH*2-1+7:0] tmp07_0_33;
	wire [WIDTH*2-1+7:0] tmp07_0_34;
	wire [WIDTH*2-1+7:0] tmp07_0_35;
	wire [WIDTH*2-1+7:0] tmp07_0_36;
	wire [WIDTH*2-1+7:0] tmp07_0_37;
	wire [WIDTH*2-1+7:0] tmp07_0_38;
	wire [WIDTH*2-1+7:0] tmp07_0_39;
	wire [WIDTH*2-1+7:0] tmp07_0_40;
	wire [WIDTH*2-1+7:0] tmp07_0_41;
	wire [WIDTH*2-1+7:0] tmp07_0_42;
	wire [WIDTH*2-1+7:0] tmp07_0_43;
	wire [WIDTH*2-1+7:0] tmp07_0_44;
	wire [WIDTH*2-1+7:0] tmp07_0_45;
	wire [WIDTH*2-1+7:0] tmp07_0_46;
	wire [WIDTH*2-1+7:0] tmp07_0_47;
	wire [WIDTH*2-1+7:0] tmp07_0_48;
	wire [WIDTH*2-1+7:0] tmp07_0_49;
	wire [WIDTH*2-1+7:0] tmp07_0_50;
	wire [WIDTH*2-1+7:0] tmp07_0_51;
	wire [WIDTH*2-1+7:0] tmp07_0_52;
	wire [WIDTH*2-1+7:0] tmp07_0_53;
	wire [WIDTH*2-1+7:0] tmp07_0_54;
	wire [WIDTH*2-1+7:0] tmp07_0_55;
	wire [WIDTH*2-1+7:0] tmp07_0_56;
	wire [WIDTH*2-1+7:0] tmp07_0_57;
	wire [WIDTH*2-1+7:0] tmp07_0_58;
	wire [WIDTH*2-1+7:0] tmp07_0_59;
	wire [WIDTH*2-1+7:0] tmp07_0_60;
	wire [WIDTH*2-1+7:0] tmp07_0_61;
	wire [WIDTH*2-1+7:0] tmp07_0_62;
	wire [WIDTH*2-1+7:0] tmp07_0_63;
	wire [WIDTH*2-1+7:0] tmp07_0_64;
	wire [WIDTH*2-1+7:0] tmp07_0_65;
	wire [WIDTH*2-1+7:0] tmp07_0_66;
	wire [WIDTH*2-1+7:0] tmp07_0_67;
	wire [WIDTH*2-1+7:0] tmp07_0_68;
	wire [WIDTH*2-1+7:0] tmp07_0_69;
	wire [WIDTH*2-1+7:0] tmp07_0_70;
	wire [WIDTH*2-1+7:0] tmp07_0_71;
	wire [WIDTH*2-1+7:0] tmp07_0_72;
	wire [WIDTH*2-1+7:0] tmp07_0_73;
	wire [WIDTH*2-1+7:0] tmp07_0_74;
	wire [WIDTH*2-1+7:0] tmp07_0_75;
	wire [WIDTH*2-1+7:0] tmp07_0_76;
	wire [WIDTH*2-1+7:0] tmp07_0_77;
	wire [WIDTH*2-1+7:0] tmp07_0_78;
	wire [WIDTH*2-1+7:0] tmp07_0_79;
	wire [WIDTH*2-1+7:0] tmp07_0_80;
	wire [WIDTH*2-1+7:0] tmp07_0_81;
	wire [WIDTH*2-1+7:0] tmp07_0_82;
	wire [WIDTH*2-1+7:0] tmp07_0_83;

	booth_0002 #(.WIDTH(WIDTH)) mul00000000(.x(x_0), .z(tmp00_0_0));
	booth_0010 #(.WIDTH(WIDTH)) mul00000001(.x(x_1), .z(tmp00_1_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000002(.x(x_2), .z(tmp00_2_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000003(.x(x_3), .z(tmp00_3_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000004(.x(x_4), .z(tmp00_4_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000005(.x(x_5), .z(tmp00_5_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000006(.x(x_6), .z(tmp00_6_0));
	booth_0012 #(.WIDTH(WIDTH)) mul00000007(.x(x_7), .z(tmp00_7_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000008(.x(x_8), .z(tmp00_8_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000009(.x(x_9), .z(tmp00_9_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000010(.x(x_10), .z(tmp00_10_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000011(.x(x_11), .z(tmp00_11_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000012(.x(x_12), .z(tmp00_12_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000013(.x(x_13), .z(tmp00_13_0));
	booth_0002 #(.WIDTH(WIDTH)) mul00000014(.x(x_14), .z(tmp00_14_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000015(.x(x_15), .z(tmp00_15_0));
	booth__006 #(.WIDTH(WIDTH)) mul00000016(.x(x_16), .z(tmp00_16_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000017(.x(x_17), .z(tmp00_17_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000018(.x(x_18), .z(tmp00_18_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000019(.x(x_19), .z(tmp00_19_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000020(.x(x_20), .z(tmp00_20_0));
	booth__010 #(.WIDTH(WIDTH)) mul00000021(.x(x_21), .z(tmp00_21_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000022(.x(x_22), .z(tmp00_22_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000023(.x(x_23), .z(tmp00_23_0));
	booth__002 #(.WIDTH(WIDTH)) mul00000024(.x(x_24), .z(tmp00_24_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000025(.x(x_25), .z(tmp00_25_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000026(.x(x_26), .z(tmp00_26_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000027(.x(x_27), .z(tmp00_27_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000028(.x(x_28), .z(tmp00_28_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000029(.x(x_29), .z(tmp00_29_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000030(.x(x_30), .z(tmp00_30_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000031(.x(x_31), .z(tmp00_31_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000032(.x(x_32), .z(tmp00_32_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000033(.x(x_33), .z(tmp00_33_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000034(.x(x_34), .z(tmp00_34_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000035(.x(x_35), .z(tmp00_35_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000036(.x(x_36), .z(tmp00_36_0));
	booth_0002 #(.WIDTH(WIDTH)) mul00000037(.x(x_37), .z(tmp00_37_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000038(.x(x_38), .z(tmp00_38_0));
	booth__010 #(.WIDTH(WIDTH)) mul00000039(.x(x_39), .z(tmp00_39_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000040(.x(x_40), .z(tmp00_40_0));
	booth__006 #(.WIDTH(WIDTH)) mul00000041(.x(x_41), .z(tmp00_41_0));
	booth_0012 #(.WIDTH(WIDTH)) mul00000042(.x(x_42), .z(tmp00_42_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000043(.x(x_43), .z(tmp00_43_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000044(.x(x_44), .z(tmp00_44_0));
	booth_0010 #(.WIDTH(WIDTH)) mul00000045(.x(x_45), .z(tmp00_45_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000046(.x(x_46), .z(tmp00_46_0));
	booth_0016 #(.WIDTH(WIDTH)) mul00000047(.x(x_47), .z(tmp00_47_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000048(.x(x_48), .z(tmp00_48_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000049(.x(x_49), .z(tmp00_49_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000050(.x(x_50), .z(tmp00_50_0));
	booth_0002 #(.WIDTH(WIDTH)) mul00000051(.x(x_51), .z(tmp00_51_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000052(.x(x_52), .z(tmp00_52_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000053(.x(x_53), .z(tmp00_53_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000054(.x(x_54), .z(tmp00_54_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000055(.x(x_55), .z(tmp00_55_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000056(.x(x_56), .z(tmp00_56_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000057(.x(x_57), .z(tmp00_57_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000058(.x(x_58), .z(tmp00_58_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000059(.x(x_59), .z(tmp00_59_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000060(.x(x_60), .z(tmp00_60_0));
	booth_0010 #(.WIDTH(WIDTH)) mul00000061(.x(x_61), .z(tmp00_61_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000062(.x(x_62), .z(tmp00_62_0));
	booth__010 #(.WIDTH(WIDTH)) mul00000063(.x(x_63), .z(tmp00_63_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000064(.x(x_64), .z(tmp00_64_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000065(.x(x_65), .z(tmp00_65_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000066(.x(x_66), .z(tmp00_66_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000067(.x(x_67), .z(tmp00_67_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000068(.x(x_68), .z(tmp00_68_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000069(.x(x_69), .z(tmp00_69_0));
	booth__006 #(.WIDTH(WIDTH)) mul00000070(.x(x_70), .z(tmp00_70_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000071(.x(x_71), .z(tmp00_71_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000072(.x(x_72), .z(tmp00_72_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000073(.x(x_73), .z(tmp00_73_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000074(.x(x_74), .z(tmp00_74_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000075(.x(x_75), .z(tmp00_75_0));
	booth_0010 #(.WIDTH(WIDTH)) mul00000076(.x(x_76), .z(tmp00_76_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000077(.x(x_77), .z(tmp00_77_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000078(.x(x_78), .z(tmp00_78_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000079(.x(x_79), .z(tmp00_79_0));
	booth_0012 #(.WIDTH(WIDTH)) mul00000080(.x(x_80), .z(tmp00_80_0));
	booth_0002 #(.WIDTH(WIDTH)) mul00000081(.x(x_81), .z(tmp00_81_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000082(.x(x_82), .z(tmp00_82_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000083(.x(x_83), .z(tmp00_83_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000084(.x(x_84), .z(tmp00_84_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000085(.x(x_85), .z(tmp00_85_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000086(.x(x_86), .z(tmp00_86_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000087(.x(x_87), .z(tmp00_87_0));
	booth__010 #(.WIDTH(WIDTH)) mul00000088(.x(x_88), .z(tmp00_88_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000089(.x(x_89), .z(tmp00_89_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000090(.x(x_90), .z(tmp00_90_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000091(.x(x_91), .z(tmp00_91_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000092(.x(x_92), .z(tmp00_92_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000093(.x(x_93), .z(tmp00_93_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000094(.x(x_94), .z(tmp00_94_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000095(.x(x_95), .z(tmp00_95_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000096(.x(x_96), .z(tmp00_96_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000097(.x(x_97), .z(tmp00_97_0));
	booth_0012 #(.WIDTH(WIDTH)) mul00000098(.x(x_98), .z(tmp00_98_0));
	booth__006 #(.WIDTH(WIDTH)) mul00000099(.x(x_99), .z(tmp00_99_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000100(.x(x_100), .z(tmp00_100_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000101(.x(x_101), .z(tmp00_101_0));
	booth_0002 #(.WIDTH(WIDTH)) mul00000102(.x(x_102), .z(tmp00_102_0));
	booth__002 #(.WIDTH(WIDTH)) mul00000103(.x(x_103), .z(tmp00_103_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000104(.x(x_104), .z(tmp00_104_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000105(.x(x_105), .z(tmp00_105_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000106(.x(x_106), .z(tmp00_106_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000107(.x(x_107), .z(tmp00_107_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000108(.x(x_108), .z(tmp00_108_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000109(.x(x_109), .z(tmp00_109_0));
	booth__002 #(.WIDTH(WIDTH)) mul00000110(.x(x_110), .z(tmp00_110_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000111(.x(x_111), .z(tmp00_111_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000112(.x(x_112), .z(tmp00_112_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000113(.x(x_113), .z(tmp00_113_0));
	booth_0010 #(.WIDTH(WIDTH)) mul00000114(.x(x_114), .z(tmp00_114_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000115(.x(x_115), .z(tmp00_115_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000116(.x(x_116), .z(tmp00_116_0));
	booth__002 #(.WIDTH(WIDTH)) mul00000117(.x(x_117), .z(tmp00_117_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000118(.x(x_118), .z(tmp00_118_0));
	booth_0016 #(.WIDTH(WIDTH)) mul00000119(.x(x_119), .z(tmp00_119_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000120(.x(x_120), .z(tmp00_120_0));
	booth_0012 #(.WIDTH(WIDTH)) mul00000121(.x(x_121), .z(tmp00_121_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000122(.x(x_122), .z(tmp00_122_0));
	booth__010 #(.WIDTH(WIDTH)) mul00000123(.x(x_123), .z(tmp00_123_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000124(.x(x_124), .z(tmp00_124_0));
	booth__002 #(.WIDTH(WIDTH)) mul00000125(.x(x_125), .z(tmp00_125_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000126(.x(x_126), .z(tmp00_126_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000127(.x(x_127), .z(tmp00_127_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00010000(.x(x_0), .z(tmp00_0_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010001(.x(x_1), .z(tmp00_1_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010002(.x(x_2), .z(tmp00_2_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010003(.x(x_3), .z(tmp00_3_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010004(.x(x_4), .z(tmp00_4_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010005(.x(x_5), .z(tmp00_5_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010006(.x(x_6), .z(tmp00_6_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010007(.x(x_7), .z(tmp00_7_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010008(.x(x_8), .z(tmp00_8_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010009(.x(x_9), .z(tmp00_9_1));
	booth__010 #(.WIDTH(WIDTH)) mul00010010(.x(x_10), .z(tmp00_10_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010011(.x(x_11), .z(tmp00_11_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010012(.x(x_12), .z(tmp00_12_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010013(.x(x_13), .z(tmp00_13_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010014(.x(x_14), .z(tmp00_14_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010015(.x(x_15), .z(tmp00_15_1));
	booth__010 #(.WIDTH(WIDTH)) mul00010016(.x(x_16), .z(tmp00_16_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010017(.x(x_17), .z(tmp00_17_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010018(.x(x_18), .z(tmp00_18_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010019(.x(x_19), .z(tmp00_19_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010020(.x(x_20), .z(tmp00_20_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010021(.x(x_21), .z(tmp00_21_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010022(.x(x_22), .z(tmp00_22_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010023(.x(x_23), .z(tmp00_23_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010024(.x(x_24), .z(tmp00_24_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010025(.x(x_25), .z(tmp00_25_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010026(.x(x_26), .z(tmp00_26_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010027(.x(x_27), .z(tmp00_27_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010028(.x(x_28), .z(tmp00_28_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010029(.x(x_29), .z(tmp00_29_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010030(.x(x_30), .z(tmp00_30_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010031(.x(x_31), .z(tmp00_31_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010032(.x(x_32), .z(tmp00_32_1));
	booth__002 #(.WIDTH(WIDTH)) mul00010033(.x(x_33), .z(tmp00_33_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010034(.x(x_34), .z(tmp00_34_1));
	booth_0012 #(.WIDTH(WIDTH)) mul00010035(.x(x_35), .z(tmp00_35_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010036(.x(x_36), .z(tmp00_36_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010037(.x(x_37), .z(tmp00_37_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010038(.x(x_38), .z(tmp00_38_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010039(.x(x_39), .z(tmp00_39_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010040(.x(x_40), .z(tmp00_40_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010041(.x(x_41), .z(tmp00_41_1));
	booth_0012 #(.WIDTH(WIDTH)) mul00010042(.x(x_42), .z(tmp00_42_1));
	booth__010 #(.WIDTH(WIDTH)) mul00010043(.x(x_43), .z(tmp00_43_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010044(.x(x_44), .z(tmp00_44_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010045(.x(x_45), .z(tmp00_45_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010046(.x(x_46), .z(tmp00_46_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010047(.x(x_47), .z(tmp00_47_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010048(.x(x_48), .z(tmp00_48_1));
	booth_0016 #(.WIDTH(WIDTH)) mul00010049(.x(x_49), .z(tmp00_49_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010050(.x(x_50), .z(tmp00_50_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010051(.x(x_51), .z(tmp00_51_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010052(.x(x_52), .z(tmp00_52_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010053(.x(x_53), .z(tmp00_53_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010054(.x(x_54), .z(tmp00_54_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010055(.x(x_55), .z(tmp00_55_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010056(.x(x_56), .z(tmp00_56_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010057(.x(x_57), .z(tmp00_57_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010058(.x(x_58), .z(tmp00_58_1));
	booth__002 #(.WIDTH(WIDTH)) mul00010059(.x(x_59), .z(tmp00_59_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010060(.x(x_60), .z(tmp00_60_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010061(.x(x_61), .z(tmp00_61_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010062(.x(x_62), .z(tmp00_62_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010063(.x(x_63), .z(tmp00_63_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010064(.x(x_64), .z(tmp00_64_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010065(.x(x_65), .z(tmp00_65_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010066(.x(x_66), .z(tmp00_66_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010067(.x(x_67), .z(tmp00_67_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010068(.x(x_68), .z(tmp00_68_1));
	booth__010 #(.WIDTH(WIDTH)) mul00010069(.x(x_69), .z(tmp00_69_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010070(.x(x_70), .z(tmp00_70_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010071(.x(x_71), .z(tmp00_71_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010072(.x(x_72), .z(tmp00_72_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010073(.x(x_73), .z(tmp00_73_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010074(.x(x_74), .z(tmp00_74_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010075(.x(x_75), .z(tmp00_75_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010076(.x(x_76), .z(tmp00_76_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010077(.x(x_77), .z(tmp00_77_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010078(.x(x_78), .z(tmp00_78_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010079(.x(x_79), .z(tmp00_79_1));
	booth_0012 #(.WIDTH(WIDTH)) mul00010080(.x(x_80), .z(tmp00_80_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010081(.x(x_81), .z(tmp00_81_1));
	booth__012 #(.WIDTH(WIDTH)) mul00010082(.x(x_82), .z(tmp00_82_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010083(.x(x_83), .z(tmp00_83_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010084(.x(x_84), .z(tmp00_84_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010085(.x(x_85), .z(tmp00_85_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010086(.x(x_86), .z(tmp00_86_1));
	booth_0012 #(.WIDTH(WIDTH)) mul00010087(.x(x_87), .z(tmp00_87_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010088(.x(x_88), .z(tmp00_88_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010089(.x(x_89), .z(tmp00_89_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010090(.x(x_90), .z(tmp00_90_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010091(.x(x_91), .z(tmp00_91_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010092(.x(x_92), .z(tmp00_92_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010093(.x(x_93), .z(tmp00_93_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010094(.x(x_94), .z(tmp00_94_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010095(.x(x_95), .z(tmp00_95_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010096(.x(x_96), .z(tmp00_96_1));
	booth__010 #(.WIDTH(WIDTH)) mul00010097(.x(x_97), .z(tmp00_97_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010098(.x(x_98), .z(tmp00_98_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010099(.x(x_99), .z(tmp00_99_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010100(.x(x_100), .z(tmp00_100_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010101(.x(x_101), .z(tmp00_101_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010102(.x(x_102), .z(tmp00_102_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010103(.x(x_103), .z(tmp00_103_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010104(.x(x_104), .z(tmp00_104_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010105(.x(x_105), .z(tmp00_105_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010106(.x(x_106), .z(tmp00_106_1));
	booth__002 #(.WIDTH(WIDTH)) mul00010107(.x(x_107), .z(tmp00_107_1));
	booth__012 #(.WIDTH(WIDTH)) mul00010108(.x(x_108), .z(tmp00_108_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010109(.x(x_109), .z(tmp00_109_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010110(.x(x_110), .z(tmp00_110_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010111(.x(x_111), .z(tmp00_111_1));
	booth__012 #(.WIDTH(WIDTH)) mul00010112(.x(x_112), .z(tmp00_112_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010113(.x(x_113), .z(tmp00_113_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010114(.x(x_114), .z(tmp00_114_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010115(.x(x_115), .z(tmp00_115_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010116(.x(x_116), .z(tmp00_116_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010117(.x(x_117), .z(tmp00_117_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010118(.x(x_118), .z(tmp00_118_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010119(.x(x_119), .z(tmp00_119_1));
	booth__012 #(.WIDTH(WIDTH)) mul00010120(.x(x_120), .z(tmp00_120_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010121(.x(x_121), .z(tmp00_121_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010122(.x(x_122), .z(tmp00_122_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010123(.x(x_123), .z(tmp00_123_1));
	booth_0010 #(.WIDTH(WIDTH)) mul00010124(.x(x_124), .z(tmp00_124_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010125(.x(x_125), .z(tmp00_125_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010126(.x(x_126), .z(tmp00_126_1));
	booth_0012 #(.WIDTH(WIDTH)) mul00010127(.x(x_127), .z(tmp00_127_1));
	booth__008 #(.WIDTH(WIDTH)) mul00020000(.x(x_0), .z(tmp00_0_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020001(.x(x_1), .z(tmp00_1_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020002(.x(x_2), .z(tmp00_2_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020003(.x(x_3), .z(tmp00_3_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020004(.x(x_4), .z(tmp00_4_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020005(.x(x_5), .z(tmp00_5_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020006(.x(x_6), .z(tmp00_6_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020007(.x(x_7), .z(tmp00_7_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020008(.x(x_8), .z(tmp00_8_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020009(.x(x_9), .z(tmp00_9_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020010(.x(x_10), .z(tmp00_10_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020011(.x(x_11), .z(tmp00_11_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020012(.x(x_12), .z(tmp00_12_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020013(.x(x_13), .z(tmp00_13_2));
	booth_0010 #(.WIDTH(WIDTH)) mul00020014(.x(x_14), .z(tmp00_14_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020015(.x(x_15), .z(tmp00_15_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020016(.x(x_16), .z(tmp00_16_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020017(.x(x_17), .z(tmp00_17_2));
	booth_0012 #(.WIDTH(WIDTH)) mul00020018(.x(x_18), .z(tmp00_18_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020019(.x(x_19), .z(tmp00_19_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020020(.x(x_20), .z(tmp00_20_2));
	booth__006 #(.WIDTH(WIDTH)) mul00020021(.x(x_21), .z(tmp00_21_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020022(.x(x_22), .z(tmp00_22_2));
	booth_0014 #(.WIDTH(WIDTH)) mul00020023(.x(x_23), .z(tmp00_23_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020024(.x(x_24), .z(tmp00_24_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020025(.x(x_25), .z(tmp00_25_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020026(.x(x_26), .z(tmp00_26_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020027(.x(x_27), .z(tmp00_27_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020028(.x(x_28), .z(tmp00_28_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020029(.x(x_29), .z(tmp00_29_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020030(.x(x_30), .z(tmp00_30_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020031(.x(x_31), .z(tmp00_31_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020032(.x(x_32), .z(tmp00_32_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020033(.x(x_33), .z(tmp00_33_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020034(.x(x_34), .z(tmp00_34_2));
	booth_0010 #(.WIDTH(WIDTH)) mul00020035(.x(x_35), .z(tmp00_35_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020036(.x(x_36), .z(tmp00_36_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020037(.x(x_37), .z(tmp00_37_2));
	booth__014 #(.WIDTH(WIDTH)) mul00020038(.x(x_38), .z(tmp00_38_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020039(.x(x_39), .z(tmp00_39_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020040(.x(x_40), .z(tmp00_40_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020041(.x(x_41), .z(tmp00_41_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020042(.x(x_42), .z(tmp00_42_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020043(.x(x_43), .z(tmp00_43_2));
	booth_0010 #(.WIDTH(WIDTH)) mul00020044(.x(x_44), .z(tmp00_44_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020045(.x(x_45), .z(tmp00_45_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020046(.x(x_46), .z(tmp00_46_2));
	booth_0010 #(.WIDTH(WIDTH)) mul00020047(.x(x_47), .z(tmp00_47_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020048(.x(x_48), .z(tmp00_48_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020049(.x(x_49), .z(tmp00_49_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020050(.x(x_50), .z(tmp00_50_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020051(.x(x_51), .z(tmp00_51_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020052(.x(x_52), .z(tmp00_52_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020053(.x(x_53), .z(tmp00_53_2));
	booth_0012 #(.WIDTH(WIDTH)) mul00020054(.x(x_54), .z(tmp00_54_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020055(.x(x_55), .z(tmp00_55_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020056(.x(x_56), .z(tmp00_56_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020057(.x(x_57), .z(tmp00_57_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020058(.x(x_58), .z(tmp00_58_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020059(.x(x_59), .z(tmp00_59_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020060(.x(x_60), .z(tmp00_60_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020061(.x(x_61), .z(tmp00_61_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020062(.x(x_62), .z(tmp00_62_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020063(.x(x_63), .z(tmp00_63_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020064(.x(x_64), .z(tmp00_64_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020065(.x(x_65), .z(tmp00_65_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020066(.x(x_66), .z(tmp00_66_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020067(.x(x_67), .z(tmp00_67_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020068(.x(x_68), .z(tmp00_68_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020069(.x(x_69), .z(tmp00_69_2));
	booth_0002 #(.WIDTH(WIDTH)) mul00020070(.x(x_70), .z(tmp00_70_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020071(.x(x_71), .z(tmp00_71_2));
	booth_0012 #(.WIDTH(WIDTH)) mul00020072(.x(x_72), .z(tmp00_72_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020073(.x(x_73), .z(tmp00_73_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020074(.x(x_74), .z(tmp00_74_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020075(.x(x_75), .z(tmp00_75_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020076(.x(x_76), .z(tmp00_76_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020077(.x(x_77), .z(tmp00_77_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020078(.x(x_78), .z(tmp00_78_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020079(.x(x_79), .z(tmp00_79_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020080(.x(x_80), .z(tmp00_80_2));
	booth__012 #(.WIDTH(WIDTH)) mul00020081(.x(x_81), .z(tmp00_81_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020082(.x(x_82), .z(tmp00_82_2));
	booth__010 #(.WIDTH(WIDTH)) mul00020083(.x(x_83), .z(tmp00_83_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020084(.x(x_84), .z(tmp00_84_2));
	booth__012 #(.WIDTH(WIDTH)) mul00020085(.x(x_85), .z(tmp00_85_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020086(.x(x_86), .z(tmp00_86_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020087(.x(x_87), .z(tmp00_87_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020088(.x(x_88), .z(tmp00_88_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020089(.x(x_89), .z(tmp00_89_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020090(.x(x_90), .z(tmp00_90_2));
	booth__012 #(.WIDTH(WIDTH)) mul00020091(.x(x_91), .z(tmp00_91_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020092(.x(x_92), .z(tmp00_92_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020093(.x(x_93), .z(tmp00_93_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020094(.x(x_94), .z(tmp00_94_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020095(.x(x_95), .z(tmp00_95_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020096(.x(x_96), .z(tmp00_96_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020097(.x(x_97), .z(tmp00_97_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020098(.x(x_98), .z(tmp00_98_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020099(.x(x_99), .z(tmp00_99_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020100(.x(x_100), .z(tmp00_100_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020101(.x(x_101), .z(tmp00_101_2));
	booth__010 #(.WIDTH(WIDTH)) mul00020102(.x(x_102), .z(tmp00_102_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020103(.x(x_103), .z(tmp00_103_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020104(.x(x_104), .z(tmp00_104_2));
	booth__006 #(.WIDTH(WIDTH)) mul00020105(.x(x_105), .z(tmp00_105_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020106(.x(x_106), .z(tmp00_106_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020107(.x(x_107), .z(tmp00_107_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020108(.x(x_108), .z(tmp00_108_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020109(.x(x_109), .z(tmp00_109_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020110(.x(x_110), .z(tmp00_110_2));
	booth_0010 #(.WIDTH(WIDTH)) mul00020111(.x(x_111), .z(tmp00_111_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020112(.x(x_112), .z(tmp00_112_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020113(.x(x_113), .z(tmp00_113_2));
	booth_0016 #(.WIDTH(WIDTH)) mul00020114(.x(x_114), .z(tmp00_114_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020115(.x(x_115), .z(tmp00_115_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020116(.x(x_116), .z(tmp00_116_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020117(.x(x_117), .z(tmp00_117_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020118(.x(x_118), .z(tmp00_118_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020119(.x(x_119), .z(tmp00_119_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020120(.x(x_120), .z(tmp00_120_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020121(.x(x_121), .z(tmp00_121_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020122(.x(x_122), .z(tmp00_122_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020123(.x(x_123), .z(tmp00_123_2));
	booth_0002 #(.WIDTH(WIDTH)) mul00020124(.x(x_124), .z(tmp00_124_2));
	booth__010 #(.WIDTH(WIDTH)) mul00020125(.x(x_125), .z(tmp00_125_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020126(.x(x_126), .z(tmp00_126_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020127(.x(x_127), .z(tmp00_127_2));
	booth__010 #(.WIDTH(WIDTH)) mul00030000(.x(x_0), .z(tmp00_0_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030001(.x(x_1), .z(tmp00_1_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030002(.x(x_2), .z(tmp00_2_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030003(.x(x_3), .z(tmp00_3_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030004(.x(x_4), .z(tmp00_4_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030005(.x(x_5), .z(tmp00_5_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030006(.x(x_6), .z(tmp00_6_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030007(.x(x_7), .z(tmp00_7_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030008(.x(x_8), .z(tmp00_8_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030009(.x(x_9), .z(tmp00_9_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030010(.x(x_10), .z(tmp00_10_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030011(.x(x_11), .z(tmp00_11_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030012(.x(x_12), .z(tmp00_12_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030013(.x(x_13), .z(tmp00_13_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030014(.x(x_14), .z(tmp00_14_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030015(.x(x_15), .z(tmp00_15_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030016(.x(x_16), .z(tmp00_16_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030017(.x(x_17), .z(tmp00_17_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030018(.x(x_18), .z(tmp00_18_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030019(.x(x_19), .z(tmp00_19_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030020(.x(x_20), .z(tmp00_20_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030021(.x(x_21), .z(tmp00_21_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030022(.x(x_22), .z(tmp00_22_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030023(.x(x_23), .z(tmp00_23_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030024(.x(x_24), .z(tmp00_24_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030025(.x(x_25), .z(tmp00_25_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030026(.x(x_26), .z(tmp00_26_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030027(.x(x_27), .z(tmp00_27_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030028(.x(x_28), .z(tmp00_28_3));
	booth_0010 #(.WIDTH(WIDTH)) mul00030029(.x(x_29), .z(tmp00_29_3));
	booth_0012 #(.WIDTH(WIDTH)) mul00030030(.x(x_30), .z(tmp00_30_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030031(.x(x_31), .z(tmp00_31_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030032(.x(x_32), .z(tmp00_32_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030033(.x(x_33), .z(tmp00_33_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030034(.x(x_34), .z(tmp00_34_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030035(.x(x_35), .z(tmp00_35_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030036(.x(x_36), .z(tmp00_36_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030037(.x(x_37), .z(tmp00_37_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030038(.x(x_38), .z(tmp00_38_3));
	booth_0002 #(.WIDTH(WIDTH)) mul00030039(.x(x_39), .z(tmp00_39_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030040(.x(x_40), .z(tmp00_40_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030041(.x(x_41), .z(tmp00_41_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030042(.x(x_42), .z(tmp00_42_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030043(.x(x_43), .z(tmp00_43_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030044(.x(x_44), .z(tmp00_44_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030045(.x(x_45), .z(tmp00_45_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030046(.x(x_46), .z(tmp00_46_3));
	booth_0002 #(.WIDTH(WIDTH)) mul00030047(.x(x_47), .z(tmp00_47_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030048(.x(x_48), .z(tmp00_48_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030049(.x(x_49), .z(tmp00_49_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030050(.x(x_50), .z(tmp00_50_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030051(.x(x_51), .z(tmp00_51_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030052(.x(x_52), .z(tmp00_52_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030053(.x(x_53), .z(tmp00_53_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030054(.x(x_54), .z(tmp00_54_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030055(.x(x_55), .z(tmp00_55_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030056(.x(x_56), .z(tmp00_56_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030057(.x(x_57), .z(tmp00_57_3));
	booth_0012 #(.WIDTH(WIDTH)) mul00030058(.x(x_58), .z(tmp00_58_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030059(.x(x_59), .z(tmp00_59_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030060(.x(x_60), .z(tmp00_60_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030061(.x(x_61), .z(tmp00_61_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030062(.x(x_62), .z(tmp00_62_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030063(.x(x_63), .z(tmp00_63_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030064(.x(x_64), .z(tmp00_64_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030065(.x(x_65), .z(tmp00_65_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030066(.x(x_66), .z(tmp00_66_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030067(.x(x_67), .z(tmp00_67_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030068(.x(x_68), .z(tmp00_68_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030069(.x(x_69), .z(tmp00_69_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030070(.x(x_70), .z(tmp00_70_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030071(.x(x_71), .z(tmp00_71_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030072(.x(x_72), .z(tmp00_72_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030073(.x(x_73), .z(tmp00_73_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030074(.x(x_74), .z(tmp00_74_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030075(.x(x_75), .z(tmp00_75_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030076(.x(x_76), .z(tmp00_76_3));
	booth_0012 #(.WIDTH(WIDTH)) mul00030077(.x(x_77), .z(tmp00_77_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030078(.x(x_78), .z(tmp00_78_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030079(.x(x_79), .z(tmp00_79_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030080(.x(x_80), .z(tmp00_80_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030081(.x(x_81), .z(tmp00_81_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030082(.x(x_82), .z(tmp00_82_3));
	booth_0002 #(.WIDTH(WIDTH)) mul00030083(.x(x_83), .z(tmp00_83_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030084(.x(x_84), .z(tmp00_84_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030085(.x(x_85), .z(tmp00_85_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030086(.x(x_86), .z(tmp00_86_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030087(.x(x_87), .z(tmp00_87_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030088(.x(x_88), .z(tmp00_88_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030089(.x(x_89), .z(tmp00_89_3));
	booth__010 #(.WIDTH(WIDTH)) mul00030090(.x(x_90), .z(tmp00_90_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030091(.x(x_91), .z(tmp00_91_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030092(.x(x_92), .z(tmp00_92_3));
	booth_0010 #(.WIDTH(WIDTH)) mul00030093(.x(x_93), .z(tmp00_93_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030094(.x(x_94), .z(tmp00_94_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030095(.x(x_95), .z(tmp00_95_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030096(.x(x_96), .z(tmp00_96_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030097(.x(x_97), .z(tmp00_97_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030098(.x(x_98), .z(tmp00_98_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030099(.x(x_99), .z(tmp00_99_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030100(.x(x_100), .z(tmp00_100_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030101(.x(x_101), .z(tmp00_101_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030102(.x(x_102), .z(tmp00_102_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030103(.x(x_103), .z(tmp00_103_3));
	booth_0012 #(.WIDTH(WIDTH)) mul00030104(.x(x_104), .z(tmp00_104_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030105(.x(x_105), .z(tmp00_105_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030106(.x(x_106), .z(tmp00_106_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030107(.x(x_107), .z(tmp00_107_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030108(.x(x_108), .z(tmp00_108_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030109(.x(x_109), .z(tmp00_109_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030110(.x(x_110), .z(tmp00_110_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030111(.x(x_111), .z(tmp00_111_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030112(.x(x_112), .z(tmp00_112_3));
	booth_0010 #(.WIDTH(WIDTH)) mul00030113(.x(x_113), .z(tmp00_113_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030114(.x(x_114), .z(tmp00_114_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030115(.x(x_115), .z(tmp00_115_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030116(.x(x_116), .z(tmp00_116_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030117(.x(x_117), .z(tmp00_117_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030118(.x(x_118), .z(tmp00_118_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030119(.x(x_119), .z(tmp00_119_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030120(.x(x_120), .z(tmp00_120_3));
	booth_0012 #(.WIDTH(WIDTH)) mul00030121(.x(x_121), .z(tmp00_121_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030122(.x(x_122), .z(tmp00_122_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030123(.x(x_123), .z(tmp00_123_3));
	booth_0010 #(.WIDTH(WIDTH)) mul00030124(.x(x_124), .z(tmp00_124_3));
	booth__010 #(.WIDTH(WIDTH)) mul00030125(.x(x_125), .z(tmp00_125_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030126(.x(x_126), .z(tmp00_126_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030127(.x(x_127), .z(tmp00_127_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00040000(.x(x_0), .z(tmp00_0_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040001(.x(x_1), .z(tmp00_1_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040002(.x(x_2), .z(tmp00_2_4));
	booth__006 #(.WIDTH(WIDTH)) mul00040003(.x(x_3), .z(tmp00_3_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040004(.x(x_4), .z(tmp00_4_4));
	booth_0010 #(.WIDTH(WIDTH)) mul00040005(.x(x_5), .z(tmp00_5_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040006(.x(x_6), .z(tmp00_6_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040007(.x(x_7), .z(tmp00_7_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040008(.x(x_8), .z(tmp00_8_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040009(.x(x_9), .z(tmp00_9_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040010(.x(x_10), .z(tmp00_10_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040011(.x(x_11), .z(tmp00_11_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040012(.x(x_12), .z(tmp00_12_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040013(.x(x_13), .z(tmp00_13_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040014(.x(x_14), .z(tmp00_14_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040015(.x(x_15), .z(tmp00_15_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040016(.x(x_16), .z(tmp00_16_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040017(.x(x_17), .z(tmp00_17_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040018(.x(x_18), .z(tmp00_18_4));
	booth__010 #(.WIDTH(WIDTH)) mul00040019(.x(x_19), .z(tmp00_19_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040020(.x(x_20), .z(tmp00_20_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040021(.x(x_21), .z(tmp00_21_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040022(.x(x_22), .z(tmp00_22_4));
	booth_0002 #(.WIDTH(WIDTH)) mul00040023(.x(x_23), .z(tmp00_23_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040024(.x(x_24), .z(tmp00_24_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040025(.x(x_25), .z(tmp00_25_4));
	booth__012 #(.WIDTH(WIDTH)) mul00040026(.x(x_26), .z(tmp00_26_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040027(.x(x_27), .z(tmp00_27_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040028(.x(x_28), .z(tmp00_28_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040029(.x(x_29), .z(tmp00_29_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040030(.x(x_30), .z(tmp00_30_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040031(.x(x_31), .z(tmp00_31_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040032(.x(x_32), .z(tmp00_32_4));
	booth_0006 #(.WIDTH(WIDTH)) mul00040033(.x(x_33), .z(tmp00_33_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040034(.x(x_34), .z(tmp00_34_4));
	booth_0012 #(.WIDTH(WIDTH)) mul00040035(.x(x_35), .z(tmp00_35_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040036(.x(x_36), .z(tmp00_36_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040037(.x(x_37), .z(tmp00_37_4));
	booth_0012 #(.WIDTH(WIDTH)) mul00040038(.x(x_38), .z(tmp00_38_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040039(.x(x_39), .z(tmp00_39_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040040(.x(x_40), .z(tmp00_40_4));
	booth_0012 #(.WIDTH(WIDTH)) mul00040041(.x(x_41), .z(tmp00_41_4));
	booth_0020 #(.WIDTH(WIDTH)) mul00040042(.x(x_42), .z(tmp00_42_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040043(.x(x_43), .z(tmp00_43_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040044(.x(x_44), .z(tmp00_44_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040045(.x(x_45), .z(tmp00_45_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040046(.x(x_46), .z(tmp00_46_4));
	booth_0012 #(.WIDTH(WIDTH)) mul00040047(.x(x_47), .z(tmp00_47_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040048(.x(x_48), .z(tmp00_48_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040049(.x(x_49), .z(tmp00_49_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040050(.x(x_50), .z(tmp00_50_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040051(.x(x_51), .z(tmp00_51_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040052(.x(x_52), .z(tmp00_52_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040053(.x(x_53), .z(tmp00_53_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040054(.x(x_54), .z(tmp00_54_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040055(.x(x_55), .z(tmp00_55_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040056(.x(x_56), .z(tmp00_56_4));
	booth__006 #(.WIDTH(WIDTH)) mul00040057(.x(x_57), .z(tmp00_57_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040058(.x(x_58), .z(tmp00_58_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040059(.x(x_59), .z(tmp00_59_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040060(.x(x_60), .z(tmp00_60_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040061(.x(x_61), .z(tmp00_61_4));
	booth_0006 #(.WIDTH(WIDTH)) mul00040062(.x(x_62), .z(tmp00_62_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040063(.x(x_63), .z(tmp00_63_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040064(.x(x_64), .z(tmp00_64_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040065(.x(x_65), .z(tmp00_65_4));
	booth_0014 #(.WIDTH(WIDTH)) mul00040066(.x(x_66), .z(tmp00_66_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040067(.x(x_67), .z(tmp00_67_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040068(.x(x_68), .z(tmp00_68_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040069(.x(x_69), .z(tmp00_69_4));
	booth__010 #(.WIDTH(WIDTH)) mul00040070(.x(x_70), .z(tmp00_70_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040071(.x(x_71), .z(tmp00_71_4));
	booth_0002 #(.WIDTH(WIDTH)) mul00040072(.x(x_72), .z(tmp00_72_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040073(.x(x_73), .z(tmp00_73_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040074(.x(x_74), .z(tmp00_74_4));
	booth__012 #(.WIDTH(WIDTH)) mul00040075(.x(x_75), .z(tmp00_75_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040076(.x(x_76), .z(tmp00_76_4));
	booth_0010 #(.WIDTH(WIDTH)) mul00040077(.x(x_77), .z(tmp00_77_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040078(.x(x_78), .z(tmp00_78_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040079(.x(x_79), .z(tmp00_79_4));
	booth_0016 #(.WIDTH(WIDTH)) mul00040080(.x(x_80), .z(tmp00_80_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040081(.x(x_81), .z(tmp00_81_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040082(.x(x_82), .z(tmp00_82_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040083(.x(x_83), .z(tmp00_83_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040084(.x(x_84), .z(tmp00_84_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040085(.x(x_85), .z(tmp00_85_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040086(.x(x_86), .z(tmp00_86_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040087(.x(x_87), .z(tmp00_87_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040088(.x(x_88), .z(tmp00_88_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040089(.x(x_89), .z(tmp00_89_4));
	booth_0012 #(.WIDTH(WIDTH)) mul00040090(.x(x_90), .z(tmp00_90_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040091(.x(x_91), .z(tmp00_91_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040092(.x(x_92), .z(tmp00_92_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040093(.x(x_93), .z(tmp00_93_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040094(.x(x_94), .z(tmp00_94_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040095(.x(x_95), .z(tmp00_95_4));
	booth__012 #(.WIDTH(WIDTH)) mul00040096(.x(x_96), .z(tmp00_96_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040097(.x(x_97), .z(tmp00_97_4));
	booth_0002 #(.WIDTH(WIDTH)) mul00040098(.x(x_98), .z(tmp00_98_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040099(.x(x_99), .z(tmp00_99_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040100(.x(x_100), .z(tmp00_100_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040101(.x(x_101), .z(tmp00_101_4));
	booth_0006 #(.WIDTH(WIDTH)) mul00040102(.x(x_102), .z(tmp00_102_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040103(.x(x_103), .z(tmp00_103_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040104(.x(x_104), .z(tmp00_104_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040105(.x(x_105), .z(tmp00_105_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040106(.x(x_106), .z(tmp00_106_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040107(.x(x_107), .z(tmp00_107_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040108(.x(x_108), .z(tmp00_108_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040109(.x(x_109), .z(tmp00_109_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040110(.x(x_110), .z(tmp00_110_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040111(.x(x_111), .z(tmp00_111_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040112(.x(x_112), .z(tmp00_112_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040113(.x(x_113), .z(tmp00_113_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040114(.x(x_114), .z(tmp00_114_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040115(.x(x_115), .z(tmp00_115_4));
	booth__012 #(.WIDTH(WIDTH)) mul00040116(.x(x_116), .z(tmp00_116_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040117(.x(x_117), .z(tmp00_117_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040118(.x(x_118), .z(tmp00_118_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040119(.x(x_119), .z(tmp00_119_4));
	booth__016 #(.WIDTH(WIDTH)) mul00040120(.x(x_120), .z(tmp00_120_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040121(.x(x_121), .z(tmp00_121_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040122(.x(x_122), .z(tmp00_122_4));
	booth__010 #(.WIDTH(WIDTH)) mul00040123(.x(x_123), .z(tmp00_123_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040124(.x(x_124), .z(tmp00_124_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040125(.x(x_125), .z(tmp00_125_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040126(.x(x_126), .z(tmp00_126_4));
	booth_0010 #(.WIDTH(WIDTH)) mul00040127(.x(x_127), .z(tmp00_127_4));
	booth__006 #(.WIDTH(WIDTH)) mul00050000(.x(x_0), .z(tmp00_0_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050001(.x(x_1), .z(tmp00_1_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050002(.x(x_2), .z(tmp00_2_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050003(.x(x_3), .z(tmp00_3_5));
	booth_0010 #(.WIDTH(WIDTH)) mul00050004(.x(x_4), .z(tmp00_4_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050005(.x(x_5), .z(tmp00_5_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050006(.x(x_6), .z(tmp00_6_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050007(.x(x_7), .z(tmp00_7_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050008(.x(x_8), .z(tmp00_8_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050009(.x(x_9), .z(tmp00_9_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050010(.x(x_10), .z(tmp00_10_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050011(.x(x_11), .z(tmp00_11_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050012(.x(x_12), .z(tmp00_12_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050013(.x(x_13), .z(tmp00_13_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050014(.x(x_14), .z(tmp00_14_5));
	booth__010 #(.WIDTH(WIDTH)) mul00050015(.x(x_15), .z(tmp00_15_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050016(.x(x_16), .z(tmp00_16_5));
	booth__010 #(.WIDTH(WIDTH)) mul00050017(.x(x_17), .z(tmp00_17_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050018(.x(x_18), .z(tmp00_18_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050019(.x(x_19), .z(tmp00_19_5));
	booth_0010 #(.WIDTH(WIDTH)) mul00050020(.x(x_20), .z(tmp00_20_5));
	booth_0012 #(.WIDTH(WIDTH)) mul00050021(.x(x_21), .z(tmp00_21_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050022(.x(x_22), .z(tmp00_22_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050023(.x(x_23), .z(tmp00_23_5));
	booth_0012 #(.WIDTH(WIDTH)) mul00050024(.x(x_24), .z(tmp00_24_5));
	booth__002 #(.WIDTH(WIDTH)) mul00050025(.x(x_25), .z(tmp00_25_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050026(.x(x_26), .z(tmp00_26_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050027(.x(x_27), .z(tmp00_27_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050028(.x(x_28), .z(tmp00_28_5));
	booth_0012 #(.WIDTH(WIDTH)) mul00050029(.x(x_29), .z(tmp00_29_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050030(.x(x_30), .z(tmp00_30_5));
	booth__002 #(.WIDTH(WIDTH)) mul00050031(.x(x_31), .z(tmp00_31_5));
	booth__002 #(.WIDTH(WIDTH)) mul00050032(.x(x_32), .z(tmp00_32_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050033(.x(x_33), .z(tmp00_33_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050034(.x(x_34), .z(tmp00_34_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050035(.x(x_35), .z(tmp00_35_5));
	booth__010 #(.WIDTH(WIDTH)) mul00050036(.x(x_36), .z(tmp00_36_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050037(.x(x_37), .z(tmp00_37_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050038(.x(x_38), .z(tmp00_38_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050039(.x(x_39), .z(tmp00_39_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050040(.x(x_40), .z(tmp00_40_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050041(.x(x_41), .z(tmp00_41_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050042(.x(x_42), .z(tmp00_42_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050043(.x(x_43), .z(tmp00_43_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050044(.x(x_44), .z(tmp00_44_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050045(.x(x_45), .z(tmp00_45_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050046(.x(x_46), .z(tmp00_46_5));
	booth_0006 #(.WIDTH(WIDTH)) mul00050047(.x(x_47), .z(tmp00_47_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050048(.x(x_48), .z(tmp00_48_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050049(.x(x_49), .z(tmp00_49_5));
	booth_0010 #(.WIDTH(WIDTH)) mul00050050(.x(x_50), .z(tmp00_50_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050051(.x(x_51), .z(tmp00_51_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050052(.x(x_52), .z(tmp00_52_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050053(.x(x_53), .z(tmp00_53_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050054(.x(x_54), .z(tmp00_54_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050055(.x(x_55), .z(tmp00_55_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050056(.x(x_56), .z(tmp00_56_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050057(.x(x_57), .z(tmp00_57_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050058(.x(x_58), .z(tmp00_58_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050059(.x(x_59), .z(tmp00_59_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050060(.x(x_60), .z(tmp00_60_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050061(.x(x_61), .z(tmp00_61_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050062(.x(x_62), .z(tmp00_62_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050063(.x(x_63), .z(tmp00_63_5));
	booth__002 #(.WIDTH(WIDTH)) mul00050064(.x(x_64), .z(tmp00_64_5));
	booth_0010 #(.WIDTH(WIDTH)) mul00050065(.x(x_65), .z(tmp00_65_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050066(.x(x_66), .z(tmp00_66_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050067(.x(x_67), .z(tmp00_67_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050068(.x(x_68), .z(tmp00_68_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050069(.x(x_69), .z(tmp00_69_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050070(.x(x_70), .z(tmp00_70_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050071(.x(x_71), .z(tmp00_71_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050072(.x(x_72), .z(tmp00_72_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050073(.x(x_73), .z(tmp00_73_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050074(.x(x_74), .z(tmp00_74_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050075(.x(x_75), .z(tmp00_75_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050076(.x(x_76), .z(tmp00_76_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050077(.x(x_77), .z(tmp00_77_5));
	booth_0010 #(.WIDTH(WIDTH)) mul00050078(.x(x_78), .z(tmp00_78_5));
	booth_0010 #(.WIDTH(WIDTH)) mul00050079(.x(x_79), .z(tmp00_79_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050080(.x(x_80), .z(tmp00_80_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050081(.x(x_81), .z(tmp00_81_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050082(.x(x_82), .z(tmp00_82_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050083(.x(x_83), .z(tmp00_83_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050084(.x(x_84), .z(tmp00_84_5));
	booth__010 #(.WIDTH(WIDTH)) mul00050085(.x(x_85), .z(tmp00_85_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050086(.x(x_86), .z(tmp00_86_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050087(.x(x_87), .z(tmp00_87_5));
	booth_0006 #(.WIDTH(WIDTH)) mul00050088(.x(x_88), .z(tmp00_88_5));
	booth_0012 #(.WIDTH(WIDTH)) mul00050089(.x(x_89), .z(tmp00_89_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050090(.x(x_90), .z(tmp00_90_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050091(.x(x_91), .z(tmp00_91_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050092(.x(x_92), .z(tmp00_92_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050093(.x(x_93), .z(tmp00_93_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050094(.x(x_94), .z(tmp00_94_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050095(.x(x_95), .z(tmp00_95_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050096(.x(x_96), .z(tmp00_96_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050097(.x(x_97), .z(tmp00_97_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050098(.x(x_98), .z(tmp00_98_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050099(.x(x_99), .z(tmp00_99_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050100(.x(x_100), .z(tmp00_100_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050101(.x(x_101), .z(tmp00_101_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050102(.x(x_102), .z(tmp00_102_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050103(.x(x_103), .z(tmp00_103_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050104(.x(x_104), .z(tmp00_104_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050105(.x(x_105), .z(tmp00_105_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050106(.x(x_106), .z(tmp00_106_5));
	booth_0012 #(.WIDTH(WIDTH)) mul00050107(.x(x_107), .z(tmp00_107_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050108(.x(x_108), .z(tmp00_108_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050109(.x(x_109), .z(tmp00_109_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050110(.x(x_110), .z(tmp00_110_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050111(.x(x_111), .z(tmp00_111_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050112(.x(x_112), .z(tmp00_112_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050113(.x(x_113), .z(tmp00_113_5));
	booth__008 #(.WIDTH(WIDTH)) mul00050114(.x(x_114), .z(tmp00_114_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050115(.x(x_115), .z(tmp00_115_5));
	booth__010 #(.WIDTH(WIDTH)) mul00050116(.x(x_116), .z(tmp00_116_5));
	booth__010 #(.WIDTH(WIDTH)) mul00050117(.x(x_117), .z(tmp00_117_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050118(.x(x_118), .z(tmp00_118_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050119(.x(x_119), .z(tmp00_119_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050120(.x(x_120), .z(tmp00_120_5));
	booth_0010 #(.WIDTH(WIDTH)) mul00050121(.x(x_121), .z(tmp00_121_5));
	booth__012 #(.WIDTH(WIDTH)) mul00050122(.x(x_122), .z(tmp00_122_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050123(.x(x_123), .z(tmp00_123_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050124(.x(x_124), .z(tmp00_124_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050125(.x(x_125), .z(tmp00_125_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050126(.x(x_126), .z(tmp00_126_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050127(.x(x_127), .z(tmp00_127_5));
	booth__008 #(.WIDTH(WIDTH)) mul00060000(.x(x_0), .z(tmp00_0_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060001(.x(x_1), .z(tmp00_1_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060002(.x(x_2), .z(tmp00_2_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060003(.x(x_3), .z(tmp00_3_6));
	booth_0016 #(.WIDTH(WIDTH)) mul00060004(.x(x_4), .z(tmp00_4_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060005(.x(x_5), .z(tmp00_5_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060006(.x(x_6), .z(tmp00_6_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060007(.x(x_7), .z(tmp00_7_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060008(.x(x_8), .z(tmp00_8_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060009(.x(x_9), .z(tmp00_9_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060010(.x(x_10), .z(tmp00_10_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060011(.x(x_11), .z(tmp00_11_6));
	booth_0010 #(.WIDTH(WIDTH)) mul00060012(.x(x_12), .z(tmp00_12_6));
	booth_0012 #(.WIDTH(WIDTH)) mul00060013(.x(x_13), .z(tmp00_13_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060014(.x(x_14), .z(tmp00_14_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060015(.x(x_15), .z(tmp00_15_6));
	booth__002 #(.WIDTH(WIDTH)) mul00060016(.x(x_16), .z(tmp00_16_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060017(.x(x_17), .z(tmp00_17_6));
	booth_0010 #(.WIDTH(WIDTH)) mul00060018(.x(x_18), .z(tmp00_18_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060019(.x(x_19), .z(tmp00_19_6));
	booth_0016 #(.WIDTH(WIDTH)) mul00060020(.x(x_20), .z(tmp00_20_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060021(.x(x_21), .z(tmp00_21_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060022(.x(x_22), .z(tmp00_22_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060023(.x(x_23), .z(tmp00_23_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060024(.x(x_24), .z(tmp00_24_6));
	booth__012 #(.WIDTH(WIDTH)) mul00060025(.x(x_25), .z(tmp00_25_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060026(.x(x_26), .z(tmp00_26_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060027(.x(x_27), .z(tmp00_27_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060028(.x(x_28), .z(tmp00_28_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060029(.x(x_29), .z(tmp00_29_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060030(.x(x_30), .z(tmp00_30_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060031(.x(x_31), .z(tmp00_31_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060032(.x(x_32), .z(tmp00_32_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060033(.x(x_33), .z(tmp00_33_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060034(.x(x_34), .z(tmp00_34_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060035(.x(x_35), .z(tmp00_35_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060036(.x(x_36), .z(tmp00_36_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060037(.x(x_37), .z(tmp00_37_6));
	booth__002 #(.WIDTH(WIDTH)) mul00060038(.x(x_38), .z(tmp00_38_6));
	booth__014 #(.WIDTH(WIDTH)) mul00060039(.x(x_39), .z(tmp00_39_6));
	booth_0010 #(.WIDTH(WIDTH)) mul00060040(.x(x_40), .z(tmp00_40_6));
	booth__006 #(.WIDTH(WIDTH)) mul00060041(.x(x_41), .z(tmp00_41_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060042(.x(x_42), .z(tmp00_42_6));
	booth__006 #(.WIDTH(WIDTH)) mul00060043(.x(x_43), .z(tmp00_43_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060044(.x(x_44), .z(tmp00_44_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060045(.x(x_45), .z(tmp00_45_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060046(.x(x_46), .z(tmp00_46_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060047(.x(x_47), .z(tmp00_47_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060048(.x(x_48), .z(tmp00_48_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060049(.x(x_49), .z(tmp00_49_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060050(.x(x_50), .z(tmp00_50_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060051(.x(x_51), .z(tmp00_51_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060052(.x(x_52), .z(tmp00_52_6));
	booth__010 #(.WIDTH(WIDTH)) mul00060053(.x(x_53), .z(tmp00_53_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060054(.x(x_54), .z(tmp00_54_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060055(.x(x_55), .z(tmp00_55_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060056(.x(x_56), .z(tmp00_56_6));
	booth_0012 #(.WIDTH(WIDTH)) mul00060057(.x(x_57), .z(tmp00_57_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060058(.x(x_58), .z(tmp00_58_6));
	booth__012 #(.WIDTH(WIDTH)) mul00060059(.x(x_59), .z(tmp00_59_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060060(.x(x_60), .z(tmp00_60_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060061(.x(x_61), .z(tmp00_61_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060062(.x(x_62), .z(tmp00_62_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060063(.x(x_63), .z(tmp00_63_6));
	booth_0006 #(.WIDTH(WIDTH)) mul00060064(.x(x_64), .z(tmp00_64_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060065(.x(x_65), .z(tmp00_65_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060066(.x(x_66), .z(tmp00_66_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060067(.x(x_67), .z(tmp00_67_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060068(.x(x_68), .z(tmp00_68_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060069(.x(x_69), .z(tmp00_69_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060070(.x(x_70), .z(tmp00_70_6));
	booth__002 #(.WIDTH(WIDTH)) mul00060071(.x(x_71), .z(tmp00_71_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060072(.x(x_72), .z(tmp00_72_6));
	booth_0010 #(.WIDTH(WIDTH)) mul00060073(.x(x_73), .z(tmp00_73_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060074(.x(x_74), .z(tmp00_74_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060075(.x(x_75), .z(tmp00_75_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060076(.x(x_76), .z(tmp00_76_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060077(.x(x_77), .z(tmp00_77_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060078(.x(x_78), .z(tmp00_78_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060079(.x(x_79), .z(tmp00_79_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060080(.x(x_80), .z(tmp00_80_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060081(.x(x_81), .z(tmp00_81_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060082(.x(x_82), .z(tmp00_82_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060083(.x(x_83), .z(tmp00_83_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060084(.x(x_84), .z(tmp00_84_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060085(.x(x_85), .z(tmp00_85_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060086(.x(x_86), .z(tmp00_86_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060087(.x(x_87), .z(tmp00_87_6));
	booth_0012 #(.WIDTH(WIDTH)) mul00060088(.x(x_88), .z(tmp00_88_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060089(.x(x_89), .z(tmp00_89_6));
	booth__002 #(.WIDTH(WIDTH)) mul00060090(.x(x_90), .z(tmp00_90_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060091(.x(x_91), .z(tmp00_91_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060092(.x(x_92), .z(tmp00_92_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060093(.x(x_93), .z(tmp00_93_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060094(.x(x_94), .z(tmp00_94_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060095(.x(x_95), .z(tmp00_95_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060096(.x(x_96), .z(tmp00_96_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060097(.x(x_97), .z(tmp00_97_6));
	booth_0006 #(.WIDTH(WIDTH)) mul00060098(.x(x_98), .z(tmp00_98_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060099(.x(x_99), .z(tmp00_99_6));
	booth_0012 #(.WIDTH(WIDTH)) mul00060100(.x(x_100), .z(tmp00_100_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060101(.x(x_101), .z(tmp00_101_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060102(.x(x_102), .z(tmp00_102_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060103(.x(x_103), .z(tmp00_103_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060104(.x(x_104), .z(tmp00_104_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060105(.x(x_105), .z(tmp00_105_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060106(.x(x_106), .z(tmp00_106_6));
	booth__006 #(.WIDTH(WIDTH)) mul00060107(.x(x_107), .z(tmp00_107_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060108(.x(x_108), .z(tmp00_108_6));
	booth_0016 #(.WIDTH(WIDTH)) mul00060109(.x(x_109), .z(tmp00_109_6));
	booth_0016 #(.WIDTH(WIDTH)) mul00060110(.x(x_110), .z(tmp00_110_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060111(.x(x_111), .z(tmp00_111_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060112(.x(x_112), .z(tmp00_112_6));
	booth__016 #(.WIDTH(WIDTH)) mul00060113(.x(x_113), .z(tmp00_113_6));
	booth__006 #(.WIDTH(WIDTH)) mul00060114(.x(x_114), .z(tmp00_114_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060115(.x(x_115), .z(tmp00_115_6));
	booth__002 #(.WIDTH(WIDTH)) mul00060116(.x(x_116), .z(tmp00_116_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060117(.x(x_117), .z(tmp00_117_6));
	booth_0012 #(.WIDTH(WIDTH)) mul00060118(.x(x_118), .z(tmp00_118_6));
	booth_0016 #(.WIDTH(WIDTH)) mul00060119(.x(x_119), .z(tmp00_119_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060120(.x(x_120), .z(tmp00_120_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060121(.x(x_121), .z(tmp00_121_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060122(.x(x_122), .z(tmp00_122_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060123(.x(x_123), .z(tmp00_123_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060124(.x(x_124), .z(tmp00_124_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060125(.x(x_125), .z(tmp00_125_6));
	booth__008 #(.WIDTH(WIDTH)) mul00060126(.x(x_126), .z(tmp00_126_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060127(.x(x_127), .z(tmp00_127_6));
	booth__004 #(.WIDTH(WIDTH)) mul00070000(.x(x_0), .z(tmp00_0_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070001(.x(x_1), .z(tmp00_1_7));
	booth_0002 #(.WIDTH(WIDTH)) mul00070002(.x(x_2), .z(tmp00_2_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070003(.x(x_3), .z(tmp00_3_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070004(.x(x_4), .z(tmp00_4_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070005(.x(x_5), .z(tmp00_5_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070006(.x(x_6), .z(tmp00_6_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070007(.x(x_7), .z(tmp00_7_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070008(.x(x_8), .z(tmp00_8_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070009(.x(x_9), .z(tmp00_9_7));
	booth__010 #(.WIDTH(WIDTH)) mul00070010(.x(x_10), .z(tmp00_10_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070011(.x(x_11), .z(tmp00_11_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070012(.x(x_12), .z(tmp00_12_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070013(.x(x_13), .z(tmp00_13_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070014(.x(x_14), .z(tmp00_14_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070015(.x(x_15), .z(tmp00_15_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070016(.x(x_16), .z(tmp00_16_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070017(.x(x_17), .z(tmp00_17_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070018(.x(x_18), .z(tmp00_18_7));
	booth__016 #(.WIDTH(WIDTH)) mul00070019(.x(x_19), .z(tmp00_19_7));
	booth__012 #(.WIDTH(WIDTH)) mul00070020(.x(x_20), .z(tmp00_20_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070021(.x(x_21), .z(tmp00_21_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070022(.x(x_22), .z(tmp00_22_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070023(.x(x_23), .z(tmp00_23_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070024(.x(x_24), .z(tmp00_24_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070025(.x(x_25), .z(tmp00_25_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070026(.x(x_26), .z(tmp00_26_7));
	booth__010 #(.WIDTH(WIDTH)) mul00070027(.x(x_27), .z(tmp00_27_7));
	booth_0002 #(.WIDTH(WIDTH)) mul00070028(.x(x_28), .z(tmp00_28_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070029(.x(x_29), .z(tmp00_29_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070030(.x(x_30), .z(tmp00_30_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070031(.x(x_31), .z(tmp00_31_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070032(.x(x_32), .z(tmp00_32_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070033(.x(x_33), .z(tmp00_33_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070034(.x(x_34), .z(tmp00_34_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070035(.x(x_35), .z(tmp00_35_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070036(.x(x_36), .z(tmp00_36_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070037(.x(x_37), .z(tmp00_37_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070038(.x(x_38), .z(tmp00_38_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070039(.x(x_39), .z(tmp00_39_7));
	booth__002 #(.WIDTH(WIDTH)) mul00070040(.x(x_40), .z(tmp00_40_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070041(.x(x_41), .z(tmp00_41_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070042(.x(x_42), .z(tmp00_42_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070043(.x(x_43), .z(tmp00_43_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070044(.x(x_44), .z(tmp00_44_7));
	booth__010 #(.WIDTH(WIDTH)) mul00070045(.x(x_45), .z(tmp00_45_7));
	booth__016 #(.WIDTH(WIDTH)) mul00070046(.x(x_46), .z(tmp00_46_7));
	booth_0012 #(.WIDTH(WIDTH)) mul00070047(.x(x_47), .z(tmp00_47_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070048(.x(x_48), .z(tmp00_48_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070049(.x(x_49), .z(tmp00_49_7));
	booth__010 #(.WIDTH(WIDTH)) mul00070050(.x(x_50), .z(tmp00_50_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070051(.x(x_51), .z(tmp00_51_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070052(.x(x_52), .z(tmp00_52_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070053(.x(x_53), .z(tmp00_53_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070054(.x(x_54), .z(tmp00_54_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070055(.x(x_55), .z(tmp00_55_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070056(.x(x_56), .z(tmp00_56_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070057(.x(x_57), .z(tmp00_57_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070058(.x(x_58), .z(tmp00_58_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070059(.x(x_59), .z(tmp00_59_7));
	booth__006 #(.WIDTH(WIDTH)) mul00070060(.x(x_60), .z(tmp00_60_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070061(.x(x_61), .z(tmp00_61_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070062(.x(x_62), .z(tmp00_62_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070063(.x(x_63), .z(tmp00_63_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070064(.x(x_64), .z(tmp00_64_7));
	booth__012 #(.WIDTH(WIDTH)) mul00070065(.x(x_65), .z(tmp00_65_7));
	booth__002 #(.WIDTH(WIDTH)) mul00070066(.x(x_66), .z(tmp00_66_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070067(.x(x_67), .z(tmp00_67_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070068(.x(x_68), .z(tmp00_68_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070069(.x(x_69), .z(tmp00_69_7));
	booth__002 #(.WIDTH(WIDTH)) mul00070070(.x(x_70), .z(tmp00_70_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070071(.x(x_71), .z(tmp00_71_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070072(.x(x_72), .z(tmp00_72_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070073(.x(x_73), .z(tmp00_73_7));
	booth_0012 #(.WIDTH(WIDTH)) mul00070074(.x(x_74), .z(tmp00_74_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070075(.x(x_75), .z(tmp00_75_7));
	booth_0012 #(.WIDTH(WIDTH)) mul00070076(.x(x_76), .z(tmp00_76_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070077(.x(x_77), .z(tmp00_77_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070078(.x(x_78), .z(tmp00_78_7));
	booth__006 #(.WIDTH(WIDTH)) mul00070079(.x(x_79), .z(tmp00_79_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070080(.x(x_80), .z(tmp00_80_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070081(.x(x_81), .z(tmp00_81_7));
	booth_0010 #(.WIDTH(WIDTH)) mul00070082(.x(x_82), .z(tmp00_82_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070083(.x(x_83), .z(tmp00_83_7));
	booth__006 #(.WIDTH(WIDTH)) mul00070084(.x(x_84), .z(tmp00_84_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070085(.x(x_85), .z(tmp00_85_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070086(.x(x_86), .z(tmp00_86_7));
	booth_0012 #(.WIDTH(WIDTH)) mul00070087(.x(x_87), .z(tmp00_87_7));
	booth_0012 #(.WIDTH(WIDTH)) mul00070088(.x(x_88), .z(tmp00_88_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070089(.x(x_89), .z(tmp00_89_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070090(.x(x_90), .z(tmp00_90_7));
	booth__012 #(.WIDTH(WIDTH)) mul00070091(.x(x_91), .z(tmp00_91_7));
	booth_0012 #(.WIDTH(WIDTH)) mul00070092(.x(x_92), .z(tmp00_92_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070093(.x(x_93), .z(tmp00_93_7));
	booth__012 #(.WIDTH(WIDTH)) mul00070094(.x(x_94), .z(tmp00_94_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070095(.x(x_95), .z(tmp00_95_7));
	booth__012 #(.WIDTH(WIDTH)) mul00070096(.x(x_96), .z(tmp00_96_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070097(.x(x_97), .z(tmp00_97_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070098(.x(x_98), .z(tmp00_98_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070099(.x(x_99), .z(tmp00_99_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070100(.x(x_100), .z(tmp00_100_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070101(.x(x_101), .z(tmp00_101_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070102(.x(x_102), .z(tmp00_102_7));
	booth_0010 #(.WIDTH(WIDTH)) mul00070103(.x(x_103), .z(tmp00_103_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070104(.x(x_104), .z(tmp00_104_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070105(.x(x_105), .z(tmp00_105_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070106(.x(x_106), .z(tmp00_106_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070107(.x(x_107), .z(tmp00_107_7));
	booth_0012 #(.WIDTH(WIDTH)) mul00070108(.x(x_108), .z(tmp00_108_7));
	booth__012 #(.WIDTH(WIDTH)) mul00070109(.x(x_109), .z(tmp00_109_7));
	booth__002 #(.WIDTH(WIDTH)) mul00070110(.x(x_110), .z(tmp00_110_7));
	booth_0010 #(.WIDTH(WIDTH)) mul00070111(.x(x_111), .z(tmp00_111_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070112(.x(x_112), .z(tmp00_112_7));
	booth_0014 #(.WIDTH(WIDTH)) mul00070113(.x(x_113), .z(tmp00_113_7));
	booth_0016 #(.WIDTH(WIDTH)) mul00070114(.x(x_114), .z(tmp00_114_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070115(.x(x_115), .z(tmp00_115_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070116(.x(x_116), .z(tmp00_116_7));
	booth_0002 #(.WIDTH(WIDTH)) mul00070117(.x(x_117), .z(tmp00_117_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070118(.x(x_118), .z(tmp00_118_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070119(.x(x_119), .z(tmp00_119_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070120(.x(x_120), .z(tmp00_120_7));
	booth_0002 #(.WIDTH(WIDTH)) mul00070121(.x(x_121), .z(tmp00_121_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070122(.x(x_122), .z(tmp00_122_7));
	booth_0008 #(.WIDTH(WIDTH)) mul00070123(.x(x_123), .z(tmp00_123_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070124(.x(x_124), .z(tmp00_124_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070125(.x(x_125), .z(tmp00_125_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070126(.x(x_126), .z(tmp00_126_7));
	booth__008 #(.WIDTH(WIDTH)) mul00070127(.x(x_127), .z(tmp00_127_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00080000(.x(x_0), .z(tmp00_0_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080001(.x(x_1), .z(tmp00_1_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080002(.x(x_2), .z(tmp00_2_8));
	booth_0012 #(.WIDTH(WIDTH)) mul00080003(.x(x_3), .z(tmp00_3_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080004(.x(x_4), .z(tmp00_4_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080005(.x(x_5), .z(tmp00_5_8));
	booth_0006 #(.WIDTH(WIDTH)) mul00080006(.x(x_6), .z(tmp00_6_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080007(.x(x_7), .z(tmp00_7_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080008(.x(x_8), .z(tmp00_8_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080009(.x(x_9), .z(tmp00_9_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080010(.x(x_10), .z(tmp00_10_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080011(.x(x_11), .z(tmp00_11_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080012(.x(x_12), .z(tmp00_12_8));
	booth__002 #(.WIDTH(WIDTH)) mul00080013(.x(x_13), .z(tmp00_13_8));
	booth_0006 #(.WIDTH(WIDTH)) mul00080014(.x(x_14), .z(tmp00_14_8));
	booth_0006 #(.WIDTH(WIDTH)) mul00080015(.x(x_15), .z(tmp00_15_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080016(.x(x_16), .z(tmp00_16_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080017(.x(x_17), .z(tmp00_17_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080018(.x(x_18), .z(tmp00_18_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080019(.x(x_19), .z(tmp00_19_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080020(.x(x_20), .z(tmp00_20_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080021(.x(x_21), .z(tmp00_21_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080022(.x(x_22), .z(tmp00_22_8));
	booth__006 #(.WIDTH(WIDTH)) mul00080023(.x(x_23), .z(tmp00_23_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080024(.x(x_24), .z(tmp00_24_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080025(.x(x_25), .z(tmp00_25_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080026(.x(x_26), .z(tmp00_26_8));
	booth__012 #(.WIDTH(WIDTH)) mul00080027(.x(x_27), .z(tmp00_27_8));
	booth__010 #(.WIDTH(WIDTH)) mul00080028(.x(x_28), .z(tmp00_28_8));
	booth_0010 #(.WIDTH(WIDTH)) mul00080029(.x(x_29), .z(tmp00_29_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080030(.x(x_30), .z(tmp00_30_8));
	booth_0010 #(.WIDTH(WIDTH)) mul00080031(.x(x_31), .z(tmp00_31_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080032(.x(x_32), .z(tmp00_32_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080033(.x(x_33), .z(tmp00_33_8));
	booth_0010 #(.WIDTH(WIDTH)) mul00080034(.x(x_34), .z(tmp00_34_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080035(.x(x_35), .z(tmp00_35_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080036(.x(x_36), .z(tmp00_36_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080037(.x(x_37), .z(tmp00_37_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080038(.x(x_38), .z(tmp00_38_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080039(.x(x_39), .z(tmp00_39_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080040(.x(x_40), .z(tmp00_40_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080041(.x(x_41), .z(tmp00_41_8));
	booth__002 #(.WIDTH(WIDTH)) mul00080042(.x(x_42), .z(tmp00_42_8));
	booth__006 #(.WIDTH(WIDTH)) mul00080043(.x(x_43), .z(tmp00_43_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080044(.x(x_44), .z(tmp00_44_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080045(.x(x_45), .z(tmp00_45_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080046(.x(x_46), .z(tmp00_46_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080047(.x(x_47), .z(tmp00_47_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080048(.x(x_48), .z(tmp00_48_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080049(.x(x_49), .z(tmp00_49_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080050(.x(x_50), .z(tmp00_50_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080051(.x(x_51), .z(tmp00_51_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080052(.x(x_52), .z(tmp00_52_8));
	booth__010 #(.WIDTH(WIDTH)) mul00080053(.x(x_53), .z(tmp00_53_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080054(.x(x_54), .z(tmp00_54_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080055(.x(x_55), .z(tmp00_55_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080056(.x(x_56), .z(tmp00_56_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080057(.x(x_57), .z(tmp00_57_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080058(.x(x_58), .z(tmp00_58_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080059(.x(x_59), .z(tmp00_59_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080060(.x(x_60), .z(tmp00_60_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080061(.x(x_61), .z(tmp00_61_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080062(.x(x_62), .z(tmp00_62_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080063(.x(x_63), .z(tmp00_63_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080064(.x(x_64), .z(tmp00_64_8));
	booth_0006 #(.WIDTH(WIDTH)) mul00080065(.x(x_65), .z(tmp00_65_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080066(.x(x_66), .z(tmp00_66_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080067(.x(x_67), .z(tmp00_67_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080068(.x(x_68), .z(tmp00_68_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080069(.x(x_69), .z(tmp00_69_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080070(.x(x_70), .z(tmp00_70_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080071(.x(x_71), .z(tmp00_71_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080072(.x(x_72), .z(tmp00_72_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080073(.x(x_73), .z(tmp00_73_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080074(.x(x_74), .z(tmp00_74_8));
	booth_0006 #(.WIDTH(WIDTH)) mul00080075(.x(x_75), .z(tmp00_75_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080076(.x(x_76), .z(tmp00_76_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080077(.x(x_77), .z(tmp00_77_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080078(.x(x_78), .z(tmp00_78_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080079(.x(x_79), .z(tmp00_79_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080080(.x(x_80), .z(tmp00_80_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080081(.x(x_81), .z(tmp00_81_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080082(.x(x_82), .z(tmp00_82_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080083(.x(x_83), .z(tmp00_83_8));
	booth_0010 #(.WIDTH(WIDTH)) mul00080084(.x(x_84), .z(tmp00_84_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080085(.x(x_85), .z(tmp00_85_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080086(.x(x_86), .z(tmp00_86_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080087(.x(x_87), .z(tmp00_87_8));
	booth_0010 #(.WIDTH(WIDTH)) mul00080088(.x(x_88), .z(tmp00_88_8));
	booth__002 #(.WIDTH(WIDTH)) mul00080089(.x(x_89), .z(tmp00_89_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080090(.x(x_90), .z(tmp00_90_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080091(.x(x_91), .z(tmp00_91_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080092(.x(x_92), .z(tmp00_92_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080093(.x(x_93), .z(tmp00_93_8));
	booth__002 #(.WIDTH(WIDTH)) mul00080094(.x(x_94), .z(tmp00_94_8));
	booth_0010 #(.WIDTH(WIDTH)) mul00080095(.x(x_95), .z(tmp00_95_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080096(.x(x_96), .z(tmp00_96_8));
	booth__010 #(.WIDTH(WIDTH)) mul00080097(.x(x_97), .z(tmp00_97_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080098(.x(x_98), .z(tmp00_98_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080099(.x(x_99), .z(tmp00_99_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080100(.x(x_100), .z(tmp00_100_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080101(.x(x_101), .z(tmp00_101_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080102(.x(x_102), .z(tmp00_102_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080103(.x(x_103), .z(tmp00_103_8));
	booth_0012 #(.WIDTH(WIDTH)) mul00080104(.x(x_104), .z(tmp00_104_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080105(.x(x_105), .z(tmp00_105_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080106(.x(x_106), .z(tmp00_106_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080107(.x(x_107), .z(tmp00_107_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080108(.x(x_108), .z(tmp00_108_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080109(.x(x_109), .z(tmp00_109_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080110(.x(x_110), .z(tmp00_110_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080111(.x(x_111), .z(tmp00_111_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080112(.x(x_112), .z(tmp00_112_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080113(.x(x_113), .z(tmp00_113_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080114(.x(x_114), .z(tmp00_114_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080115(.x(x_115), .z(tmp00_115_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080116(.x(x_116), .z(tmp00_116_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080117(.x(x_117), .z(tmp00_117_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080118(.x(x_118), .z(tmp00_118_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080119(.x(x_119), .z(tmp00_119_8));
	booth_0010 #(.WIDTH(WIDTH)) mul00080120(.x(x_120), .z(tmp00_120_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080121(.x(x_121), .z(tmp00_121_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080122(.x(x_122), .z(tmp00_122_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080123(.x(x_123), .z(tmp00_123_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080124(.x(x_124), .z(tmp00_124_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080125(.x(x_125), .z(tmp00_125_8));
	booth_0006 #(.WIDTH(WIDTH)) mul00080126(.x(x_126), .z(tmp00_126_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080127(.x(x_127), .z(tmp00_127_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00090000(.x(x_0), .z(tmp00_0_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090001(.x(x_1), .z(tmp00_1_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090002(.x(x_2), .z(tmp00_2_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090003(.x(x_3), .z(tmp00_3_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090004(.x(x_4), .z(tmp00_4_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090005(.x(x_5), .z(tmp00_5_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090006(.x(x_6), .z(tmp00_6_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090007(.x(x_7), .z(tmp00_7_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090008(.x(x_8), .z(tmp00_8_9));
	booth_0012 #(.WIDTH(WIDTH)) mul00090009(.x(x_9), .z(tmp00_9_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090010(.x(x_10), .z(tmp00_10_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090011(.x(x_11), .z(tmp00_11_9));
	booth_0012 #(.WIDTH(WIDTH)) mul00090012(.x(x_12), .z(tmp00_12_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090013(.x(x_13), .z(tmp00_13_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090014(.x(x_14), .z(tmp00_14_9));
	booth__010 #(.WIDTH(WIDTH)) mul00090015(.x(x_15), .z(tmp00_15_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090016(.x(x_16), .z(tmp00_16_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090017(.x(x_17), .z(tmp00_17_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090018(.x(x_18), .z(tmp00_18_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090019(.x(x_19), .z(tmp00_19_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090020(.x(x_20), .z(tmp00_20_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090021(.x(x_21), .z(tmp00_21_9));
	booth_0014 #(.WIDTH(WIDTH)) mul00090022(.x(x_22), .z(tmp00_22_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090023(.x(x_23), .z(tmp00_23_9));
	booth_0010 #(.WIDTH(WIDTH)) mul00090024(.x(x_24), .z(tmp00_24_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090025(.x(x_25), .z(tmp00_25_9));
	booth_0012 #(.WIDTH(WIDTH)) mul00090026(.x(x_26), .z(tmp00_26_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090027(.x(x_27), .z(tmp00_27_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090028(.x(x_28), .z(tmp00_28_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090029(.x(x_29), .z(tmp00_29_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090030(.x(x_30), .z(tmp00_30_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090031(.x(x_31), .z(tmp00_31_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090032(.x(x_32), .z(tmp00_32_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090033(.x(x_33), .z(tmp00_33_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090034(.x(x_34), .z(tmp00_34_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090035(.x(x_35), .z(tmp00_35_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090036(.x(x_36), .z(tmp00_36_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090037(.x(x_37), .z(tmp00_37_9));
	booth__012 #(.WIDTH(WIDTH)) mul00090038(.x(x_38), .z(tmp00_38_9));
	booth_0016 #(.WIDTH(WIDTH)) mul00090039(.x(x_39), .z(tmp00_39_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090040(.x(x_40), .z(tmp00_40_9));
	booth__012 #(.WIDTH(WIDTH)) mul00090041(.x(x_41), .z(tmp00_41_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090042(.x(x_42), .z(tmp00_42_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090043(.x(x_43), .z(tmp00_43_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090044(.x(x_44), .z(tmp00_44_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090045(.x(x_45), .z(tmp00_45_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090046(.x(x_46), .z(tmp00_46_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090047(.x(x_47), .z(tmp00_47_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090048(.x(x_48), .z(tmp00_48_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090049(.x(x_49), .z(tmp00_49_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090050(.x(x_50), .z(tmp00_50_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090051(.x(x_51), .z(tmp00_51_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090052(.x(x_52), .z(tmp00_52_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090053(.x(x_53), .z(tmp00_53_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090054(.x(x_54), .z(tmp00_54_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090055(.x(x_55), .z(tmp00_55_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090056(.x(x_56), .z(tmp00_56_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090057(.x(x_57), .z(tmp00_57_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090058(.x(x_58), .z(tmp00_58_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090059(.x(x_59), .z(tmp00_59_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090060(.x(x_60), .z(tmp00_60_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090061(.x(x_61), .z(tmp00_61_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090062(.x(x_62), .z(tmp00_62_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090063(.x(x_63), .z(tmp00_63_9));
	booth__010 #(.WIDTH(WIDTH)) mul00090064(.x(x_64), .z(tmp00_64_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090065(.x(x_65), .z(tmp00_65_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090066(.x(x_66), .z(tmp00_66_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090067(.x(x_67), .z(tmp00_67_9));
	booth_0014 #(.WIDTH(WIDTH)) mul00090068(.x(x_68), .z(tmp00_68_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090069(.x(x_69), .z(tmp00_69_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090070(.x(x_70), .z(tmp00_70_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090071(.x(x_71), .z(tmp00_71_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090072(.x(x_72), .z(tmp00_72_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090073(.x(x_73), .z(tmp00_73_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090074(.x(x_74), .z(tmp00_74_9));
	booth_0010 #(.WIDTH(WIDTH)) mul00090075(.x(x_75), .z(tmp00_75_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090076(.x(x_76), .z(tmp00_76_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090077(.x(x_77), .z(tmp00_77_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090078(.x(x_78), .z(tmp00_78_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090079(.x(x_79), .z(tmp00_79_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090080(.x(x_80), .z(tmp00_80_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090081(.x(x_81), .z(tmp00_81_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090082(.x(x_82), .z(tmp00_82_9));
	booth__010 #(.WIDTH(WIDTH)) mul00090083(.x(x_83), .z(tmp00_83_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090084(.x(x_84), .z(tmp00_84_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090085(.x(x_85), .z(tmp00_85_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090086(.x(x_86), .z(tmp00_86_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090087(.x(x_87), .z(tmp00_87_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090088(.x(x_88), .z(tmp00_88_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090089(.x(x_89), .z(tmp00_89_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090090(.x(x_90), .z(tmp00_90_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090091(.x(x_91), .z(tmp00_91_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090092(.x(x_92), .z(tmp00_92_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090093(.x(x_93), .z(tmp00_93_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090094(.x(x_94), .z(tmp00_94_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090095(.x(x_95), .z(tmp00_95_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090096(.x(x_96), .z(tmp00_96_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090097(.x(x_97), .z(tmp00_97_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090098(.x(x_98), .z(tmp00_98_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090099(.x(x_99), .z(tmp00_99_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090100(.x(x_100), .z(tmp00_100_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090101(.x(x_101), .z(tmp00_101_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090102(.x(x_102), .z(tmp00_102_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090103(.x(x_103), .z(tmp00_103_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090104(.x(x_104), .z(tmp00_104_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090105(.x(x_105), .z(tmp00_105_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090106(.x(x_106), .z(tmp00_106_9));
	booth__010 #(.WIDTH(WIDTH)) mul00090107(.x(x_107), .z(tmp00_107_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090108(.x(x_108), .z(tmp00_108_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090109(.x(x_109), .z(tmp00_109_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090110(.x(x_110), .z(tmp00_110_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090111(.x(x_111), .z(tmp00_111_9));
	booth_0010 #(.WIDTH(WIDTH)) mul00090112(.x(x_112), .z(tmp00_112_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090113(.x(x_113), .z(tmp00_113_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090114(.x(x_114), .z(tmp00_114_9));
	booth_0012 #(.WIDTH(WIDTH)) mul00090115(.x(x_115), .z(tmp00_115_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090116(.x(x_116), .z(tmp00_116_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090117(.x(x_117), .z(tmp00_117_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090118(.x(x_118), .z(tmp00_118_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090119(.x(x_119), .z(tmp00_119_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090120(.x(x_120), .z(tmp00_120_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090121(.x(x_121), .z(tmp00_121_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090122(.x(x_122), .z(tmp00_122_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090123(.x(x_123), .z(tmp00_123_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090124(.x(x_124), .z(tmp00_124_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090125(.x(x_125), .z(tmp00_125_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090126(.x(x_126), .z(tmp00_126_9));
	booth_0012 #(.WIDTH(WIDTH)) mul00090127(.x(x_127), .z(tmp00_127_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00100000(.x(x_0), .z(tmp00_0_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100001(.x(x_1), .z(tmp00_1_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100002(.x(x_2), .z(tmp00_2_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100003(.x(x_3), .z(tmp00_3_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100004(.x(x_4), .z(tmp00_4_10));
	booth__012 #(.WIDTH(WIDTH)) mul00100005(.x(x_5), .z(tmp00_5_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100006(.x(x_6), .z(tmp00_6_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100007(.x(x_7), .z(tmp00_7_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100008(.x(x_8), .z(tmp00_8_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100009(.x(x_9), .z(tmp00_9_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100010(.x(x_10), .z(tmp00_10_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100011(.x(x_11), .z(tmp00_11_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100012(.x(x_12), .z(tmp00_12_10));
	booth_0006 #(.WIDTH(WIDTH)) mul00100013(.x(x_13), .z(tmp00_13_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100014(.x(x_14), .z(tmp00_14_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100015(.x(x_15), .z(tmp00_15_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100016(.x(x_16), .z(tmp00_16_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100017(.x(x_17), .z(tmp00_17_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100018(.x(x_18), .z(tmp00_18_10));
	booth__010 #(.WIDTH(WIDTH)) mul00100019(.x(x_19), .z(tmp00_19_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100020(.x(x_20), .z(tmp00_20_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100021(.x(x_21), .z(tmp00_21_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100022(.x(x_22), .z(tmp00_22_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100023(.x(x_23), .z(tmp00_23_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100024(.x(x_24), .z(tmp00_24_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100025(.x(x_25), .z(tmp00_25_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100026(.x(x_26), .z(tmp00_26_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100027(.x(x_27), .z(tmp00_27_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100028(.x(x_28), .z(tmp00_28_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100029(.x(x_29), .z(tmp00_29_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100030(.x(x_30), .z(tmp00_30_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100031(.x(x_31), .z(tmp00_31_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100032(.x(x_32), .z(tmp00_32_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100033(.x(x_33), .z(tmp00_33_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100034(.x(x_34), .z(tmp00_34_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100035(.x(x_35), .z(tmp00_35_10));
	booth__010 #(.WIDTH(WIDTH)) mul00100036(.x(x_36), .z(tmp00_36_10));
	booth_0006 #(.WIDTH(WIDTH)) mul00100037(.x(x_37), .z(tmp00_37_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100038(.x(x_38), .z(tmp00_38_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100039(.x(x_39), .z(tmp00_39_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100040(.x(x_40), .z(tmp00_40_10));
	booth_0010 #(.WIDTH(WIDTH)) mul00100041(.x(x_41), .z(tmp00_41_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100042(.x(x_42), .z(tmp00_42_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100043(.x(x_43), .z(tmp00_43_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100044(.x(x_44), .z(tmp00_44_10));
	booth__002 #(.WIDTH(WIDTH)) mul00100045(.x(x_45), .z(tmp00_45_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100046(.x(x_46), .z(tmp00_46_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100047(.x(x_47), .z(tmp00_47_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100048(.x(x_48), .z(tmp00_48_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100049(.x(x_49), .z(tmp00_49_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100050(.x(x_50), .z(tmp00_50_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100051(.x(x_51), .z(tmp00_51_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100052(.x(x_52), .z(tmp00_52_10));
	booth_0012 #(.WIDTH(WIDTH)) mul00100053(.x(x_53), .z(tmp00_53_10));
	booth__010 #(.WIDTH(WIDTH)) mul00100054(.x(x_54), .z(tmp00_54_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100055(.x(x_55), .z(tmp00_55_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100056(.x(x_56), .z(tmp00_56_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100057(.x(x_57), .z(tmp00_57_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100058(.x(x_58), .z(tmp00_58_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100059(.x(x_59), .z(tmp00_59_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100060(.x(x_60), .z(tmp00_60_10));
	booth__010 #(.WIDTH(WIDTH)) mul00100061(.x(x_61), .z(tmp00_61_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100062(.x(x_62), .z(tmp00_62_10));
	booth_0002 #(.WIDTH(WIDTH)) mul00100063(.x(x_63), .z(tmp00_63_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100064(.x(x_64), .z(tmp00_64_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100065(.x(x_65), .z(tmp00_65_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100066(.x(x_66), .z(tmp00_66_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100067(.x(x_67), .z(tmp00_67_10));
	booth_0002 #(.WIDTH(WIDTH)) mul00100068(.x(x_68), .z(tmp00_68_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100069(.x(x_69), .z(tmp00_69_10));
	booth__006 #(.WIDTH(WIDTH)) mul00100070(.x(x_70), .z(tmp00_70_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100071(.x(x_71), .z(tmp00_71_10));
	booth__006 #(.WIDTH(WIDTH)) mul00100072(.x(x_72), .z(tmp00_72_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100073(.x(x_73), .z(tmp00_73_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100074(.x(x_74), .z(tmp00_74_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100075(.x(x_75), .z(tmp00_75_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100076(.x(x_76), .z(tmp00_76_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100077(.x(x_77), .z(tmp00_77_10));
	booth__006 #(.WIDTH(WIDTH)) mul00100078(.x(x_78), .z(tmp00_78_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100079(.x(x_79), .z(tmp00_79_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100080(.x(x_80), .z(tmp00_80_10));
	booth__002 #(.WIDTH(WIDTH)) mul00100081(.x(x_81), .z(tmp00_81_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100082(.x(x_82), .z(tmp00_82_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100083(.x(x_83), .z(tmp00_83_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100084(.x(x_84), .z(tmp00_84_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100085(.x(x_85), .z(tmp00_85_10));
	booth__006 #(.WIDTH(WIDTH)) mul00100086(.x(x_86), .z(tmp00_86_10));
	booth_0010 #(.WIDTH(WIDTH)) mul00100087(.x(x_87), .z(tmp00_87_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100088(.x(x_88), .z(tmp00_88_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100089(.x(x_89), .z(tmp00_89_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100090(.x(x_90), .z(tmp00_90_10));
	booth_0006 #(.WIDTH(WIDTH)) mul00100091(.x(x_91), .z(tmp00_91_10));
	booth__010 #(.WIDTH(WIDTH)) mul00100092(.x(x_92), .z(tmp00_92_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100093(.x(x_93), .z(tmp00_93_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100094(.x(x_94), .z(tmp00_94_10));
	booth_0006 #(.WIDTH(WIDTH)) mul00100095(.x(x_95), .z(tmp00_95_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100096(.x(x_96), .z(tmp00_96_10));
	booth__006 #(.WIDTH(WIDTH)) mul00100097(.x(x_97), .z(tmp00_97_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100098(.x(x_98), .z(tmp00_98_10));
	booth_0010 #(.WIDTH(WIDTH)) mul00100099(.x(x_99), .z(tmp00_99_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100100(.x(x_100), .z(tmp00_100_10));
	booth__012 #(.WIDTH(WIDTH)) mul00100101(.x(x_101), .z(tmp00_101_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100102(.x(x_102), .z(tmp00_102_10));
	booth__002 #(.WIDTH(WIDTH)) mul00100103(.x(x_103), .z(tmp00_103_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100104(.x(x_104), .z(tmp00_104_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100105(.x(x_105), .z(tmp00_105_10));
	booth__010 #(.WIDTH(WIDTH)) mul00100106(.x(x_106), .z(tmp00_106_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100107(.x(x_107), .z(tmp00_107_10));
	booth_0008 #(.WIDTH(WIDTH)) mul00100108(.x(x_108), .z(tmp00_108_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100109(.x(x_109), .z(tmp00_109_10));
	booth_0004 #(.WIDTH(WIDTH)) mul00100110(.x(x_110), .z(tmp00_110_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100111(.x(x_111), .z(tmp00_111_10));
	booth_0006 #(.WIDTH(WIDTH)) mul00100112(.x(x_112), .z(tmp00_112_10));
	booth__010 #(.WIDTH(WIDTH)) mul00100113(.x(x_113), .z(tmp00_113_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100114(.x(x_114), .z(tmp00_114_10));
	booth_0006 #(.WIDTH(WIDTH)) mul00100115(.x(x_115), .z(tmp00_115_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100116(.x(x_116), .z(tmp00_116_10));
	booth__010 #(.WIDTH(WIDTH)) mul00100117(.x(x_117), .z(tmp00_117_10));
	booth_0010 #(.WIDTH(WIDTH)) mul00100118(.x(x_118), .z(tmp00_118_10));
	booth__004 #(.WIDTH(WIDTH)) mul00100119(.x(x_119), .z(tmp00_119_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100120(.x(x_120), .z(tmp00_120_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100121(.x(x_121), .z(tmp00_121_10));
	booth_0010 #(.WIDTH(WIDTH)) mul00100122(.x(x_122), .z(tmp00_122_10));
	booth__008 #(.WIDTH(WIDTH)) mul00100123(.x(x_123), .z(tmp00_123_10));
	booth_0002 #(.WIDTH(WIDTH)) mul00100124(.x(x_124), .z(tmp00_124_10));
	booth__002 #(.WIDTH(WIDTH)) mul00100125(.x(x_125), .z(tmp00_125_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100126(.x(x_126), .z(tmp00_126_10));
	booth_0000 #(.WIDTH(WIDTH)) mul00100127(.x(x_127), .z(tmp00_127_10));
	booth__010 #(.WIDTH(WIDTH)) mul00110000(.x(x_0), .z(tmp00_0_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110001(.x(x_1), .z(tmp00_1_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110002(.x(x_2), .z(tmp00_2_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110003(.x(x_3), .z(tmp00_3_11));
	booth__006 #(.WIDTH(WIDTH)) mul00110004(.x(x_4), .z(tmp00_4_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110005(.x(x_5), .z(tmp00_5_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110006(.x(x_6), .z(tmp00_6_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110007(.x(x_7), .z(tmp00_7_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110008(.x(x_8), .z(tmp00_8_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110009(.x(x_9), .z(tmp00_9_11));
	booth_0002 #(.WIDTH(WIDTH)) mul00110010(.x(x_10), .z(tmp00_10_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110011(.x(x_11), .z(tmp00_11_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110012(.x(x_12), .z(tmp00_12_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110013(.x(x_13), .z(tmp00_13_11));
	booth__006 #(.WIDTH(WIDTH)) mul00110014(.x(x_14), .z(tmp00_14_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110015(.x(x_15), .z(tmp00_15_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110016(.x(x_16), .z(tmp00_16_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110017(.x(x_17), .z(tmp00_17_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110018(.x(x_18), .z(tmp00_18_11));
	booth_0006 #(.WIDTH(WIDTH)) mul00110019(.x(x_19), .z(tmp00_19_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110020(.x(x_20), .z(tmp00_20_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110021(.x(x_21), .z(tmp00_21_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110022(.x(x_22), .z(tmp00_22_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110023(.x(x_23), .z(tmp00_23_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110024(.x(x_24), .z(tmp00_24_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110025(.x(x_25), .z(tmp00_25_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110026(.x(x_26), .z(tmp00_26_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110027(.x(x_27), .z(tmp00_27_11));
	booth_0010 #(.WIDTH(WIDTH)) mul00110028(.x(x_28), .z(tmp00_28_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110029(.x(x_29), .z(tmp00_29_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110030(.x(x_30), .z(tmp00_30_11));
	booth__006 #(.WIDTH(WIDTH)) mul00110031(.x(x_31), .z(tmp00_31_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110032(.x(x_32), .z(tmp00_32_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110033(.x(x_33), .z(tmp00_33_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110034(.x(x_34), .z(tmp00_34_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110035(.x(x_35), .z(tmp00_35_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110036(.x(x_36), .z(tmp00_36_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110037(.x(x_37), .z(tmp00_37_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110038(.x(x_38), .z(tmp00_38_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110039(.x(x_39), .z(tmp00_39_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110040(.x(x_40), .z(tmp00_40_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110041(.x(x_41), .z(tmp00_41_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110042(.x(x_42), .z(tmp00_42_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110043(.x(x_43), .z(tmp00_43_11));
	booth__006 #(.WIDTH(WIDTH)) mul00110044(.x(x_44), .z(tmp00_44_11));
	booth__002 #(.WIDTH(WIDTH)) mul00110045(.x(x_45), .z(tmp00_45_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110046(.x(x_46), .z(tmp00_46_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110047(.x(x_47), .z(tmp00_47_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110048(.x(x_48), .z(tmp00_48_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110049(.x(x_49), .z(tmp00_49_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110050(.x(x_50), .z(tmp00_50_11));
	booth_0006 #(.WIDTH(WIDTH)) mul00110051(.x(x_51), .z(tmp00_51_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110052(.x(x_52), .z(tmp00_52_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110053(.x(x_53), .z(tmp00_53_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110054(.x(x_54), .z(tmp00_54_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110055(.x(x_55), .z(tmp00_55_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110056(.x(x_56), .z(tmp00_56_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110057(.x(x_57), .z(tmp00_57_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110058(.x(x_58), .z(tmp00_58_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110059(.x(x_59), .z(tmp00_59_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110060(.x(x_60), .z(tmp00_60_11));
	booth__002 #(.WIDTH(WIDTH)) mul00110061(.x(x_61), .z(tmp00_61_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110062(.x(x_62), .z(tmp00_62_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110063(.x(x_63), .z(tmp00_63_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110064(.x(x_64), .z(tmp00_64_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110065(.x(x_65), .z(tmp00_65_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110066(.x(x_66), .z(tmp00_66_11));
	booth__010 #(.WIDTH(WIDTH)) mul00110067(.x(x_67), .z(tmp00_67_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110068(.x(x_68), .z(tmp00_68_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110069(.x(x_69), .z(tmp00_69_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110070(.x(x_70), .z(tmp00_70_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110071(.x(x_71), .z(tmp00_71_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110072(.x(x_72), .z(tmp00_72_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110073(.x(x_73), .z(tmp00_73_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110074(.x(x_74), .z(tmp00_74_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110075(.x(x_75), .z(tmp00_75_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110076(.x(x_76), .z(tmp00_76_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110077(.x(x_77), .z(tmp00_77_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110078(.x(x_78), .z(tmp00_78_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110079(.x(x_79), .z(tmp00_79_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110080(.x(x_80), .z(tmp00_80_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110081(.x(x_81), .z(tmp00_81_11));
	booth__010 #(.WIDTH(WIDTH)) mul00110082(.x(x_82), .z(tmp00_82_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110083(.x(x_83), .z(tmp00_83_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110084(.x(x_84), .z(tmp00_84_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110085(.x(x_85), .z(tmp00_85_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110086(.x(x_86), .z(tmp00_86_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110087(.x(x_87), .z(tmp00_87_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110088(.x(x_88), .z(tmp00_88_11));
	booth__002 #(.WIDTH(WIDTH)) mul00110089(.x(x_89), .z(tmp00_89_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110090(.x(x_90), .z(tmp00_90_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110091(.x(x_91), .z(tmp00_91_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110092(.x(x_92), .z(tmp00_92_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110093(.x(x_93), .z(tmp00_93_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110094(.x(x_94), .z(tmp00_94_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110095(.x(x_95), .z(tmp00_95_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110096(.x(x_96), .z(tmp00_96_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110097(.x(x_97), .z(tmp00_97_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110098(.x(x_98), .z(tmp00_98_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110099(.x(x_99), .z(tmp00_99_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110100(.x(x_100), .z(tmp00_100_11));
	booth_0010 #(.WIDTH(WIDTH)) mul00110101(.x(x_101), .z(tmp00_101_11));
	booth_0010 #(.WIDTH(WIDTH)) mul00110102(.x(x_102), .z(tmp00_102_11));
	booth_0006 #(.WIDTH(WIDTH)) mul00110103(.x(x_103), .z(tmp00_103_11));
	booth_0008 #(.WIDTH(WIDTH)) mul00110104(.x(x_104), .z(tmp00_104_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110105(.x(x_105), .z(tmp00_105_11));
	booth__002 #(.WIDTH(WIDTH)) mul00110106(.x(x_106), .z(tmp00_106_11));
	booth_0010 #(.WIDTH(WIDTH)) mul00110107(.x(x_107), .z(tmp00_107_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110108(.x(x_108), .z(tmp00_108_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110109(.x(x_109), .z(tmp00_109_11));
	booth_0006 #(.WIDTH(WIDTH)) mul00110110(.x(x_110), .z(tmp00_110_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110111(.x(x_111), .z(tmp00_111_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110112(.x(x_112), .z(tmp00_112_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110113(.x(x_113), .z(tmp00_113_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110114(.x(x_114), .z(tmp00_114_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110115(.x(x_115), .z(tmp00_115_11));
	booth__010 #(.WIDTH(WIDTH)) mul00110116(.x(x_116), .z(tmp00_116_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110117(.x(x_117), .z(tmp00_117_11));
	booth__002 #(.WIDTH(WIDTH)) mul00110118(.x(x_118), .z(tmp00_118_11));
	booth__004 #(.WIDTH(WIDTH)) mul00110119(.x(x_119), .z(tmp00_119_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110120(.x(x_120), .z(tmp00_120_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110121(.x(x_121), .z(tmp00_121_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00110122(.x(x_122), .z(tmp00_122_11));
	booth_0006 #(.WIDTH(WIDTH)) mul00110123(.x(x_123), .z(tmp00_123_11));
	booth_0010 #(.WIDTH(WIDTH)) mul00110124(.x(x_124), .z(tmp00_124_11));
	booth__008 #(.WIDTH(WIDTH)) mul00110125(.x(x_125), .z(tmp00_125_11));
	booth_0010 #(.WIDTH(WIDTH)) mul00110126(.x(x_126), .z(tmp00_126_11));
	booth_0004 #(.WIDTH(WIDTH)) mul00110127(.x(x_127), .z(tmp00_127_11));
	booth_0000 #(.WIDTH(WIDTH)) mul00120000(.x(x_0), .z(tmp00_0_12));
	booth__002 #(.WIDTH(WIDTH)) mul00120001(.x(x_1), .z(tmp00_1_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120002(.x(x_2), .z(tmp00_2_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120003(.x(x_3), .z(tmp00_3_12));
	booth_0008 #(.WIDTH(WIDTH)) mul00120004(.x(x_4), .z(tmp00_4_12));
	booth_0002 #(.WIDTH(WIDTH)) mul00120005(.x(x_5), .z(tmp00_5_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120006(.x(x_6), .z(tmp00_6_12));
	booth_0010 #(.WIDTH(WIDTH)) mul00120007(.x(x_7), .z(tmp00_7_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120008(.x(x_8), .z(tmp00_8_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120009(.x(x_9), .z(tmp00_9_12));
	booth__006 #(.WIDTH(WIDTH)) mul00120010(.x(x_10), .z(tmp00_10_12));
	booth__006 #(.WIDTH(WIDTH)) mul00120011(.x(x_11), .z(tmp00_11_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120012(.x(x_12), .z(tmp00_12_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120013(.x(x_13), .z(tmp00_13_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120014(.x(x_14), .z(tmp00_14_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120015(.x(x_15), .z(tmp00_15_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120016(.x(x_16), .z(tmp00_16_12));
	booth_0008 #(.WIDTH(WIDTH)) mul00120017(.x(x_17), .z(tmp00_17_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120018(.x(x_18), .z(tmp00_18_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120019(.x(x_19), .z(tmp00_19_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120020(.x(x_20), .z(tmp00_20_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120021(.x(x_21), .z(tmp00_21_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120022(.x(x_22), .z(tmp00_22_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120023(.x(x_23), .z(tmp00_23_12));
	booth__002 #(.WIDTH(WIDTH)) mul00120024(.x(x_24), .z(tmp00_24_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120025(.x(x_25), .z(tmp00_25_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120026(.x(x_26), .z(tmp00_26_12));
	booth__010 #(.WIDTH(WIDTH)) mul00120027(.x(x_27), .z(tmp00_27_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120028(.x(x_28), .z(tmp00_28_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120029(.x(x_29), .z(tmp00_29_12));
	booth_0006 #(.WIDTH(WIDTH)) mul00120030(.x(x_30), .z(tmp00_30_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120031(.x(x_31), .z(tmp00_31_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120032(.x(x_32), .z(tmp00_32_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120033(.x(x_33), .z(tmp00_33_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120034(.x(x_34), .z(tmp00_34_12));
	booth__006 #(.WIDTH(WIDTH)) mul00120035(.x(x_35), .z(tmp00_35_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120036(.x(x_36), .z(tmp00_36_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120037(.x(x_37), .z(tmp00_37_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120038(.x(x_38), .z(tmp00_38_12));
	booth__010 #(.WIDTH(WIDTH)) mul00120039(.x(x_39), .z(tmp00_39_12));
	booth__006 #(.WIDTH(WIDTH)) mul00120040(.x(x_40), .z(tmp00_40_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120041(.x(x_41), .z(tmp00_41_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120042(.x(x_42), .z(tmp00_42_12));
	booth__012 #(.WIDTH(WIDTH)) mul00120043(.x(x_43), .z(tmp00_43_12));
	booth_0008 #(.WIDTH(WIDTH)) mul00120044(.x(x_44), .z(tmp00_44_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120045(.x(x_45), .z(tmp00_45_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120046(.x(x_46), .z(tmp00_46_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120047(.x(x_47), .z(tmp00_47_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120048(.x(x_48), .z(tmp00_48_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120049(.x(x_49), .z(tmp00_49_12));
	booth__010 #(.WIDTH(WIDTH)) mul00120050(.x(x_50), .z(tmp00_50_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120051(.x(x_51), .z(tmp00_51_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120052(.x(x_52), .z(tmp00_52_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120053(.x(x_53), .z(tmp00_53_12));
	booth_0006 #(.WIDTH(WIDTH)) mul00120054(.x(x_54), .z(tmp00_54_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120055(.x(x_55), .z(tmp00_55_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120056(.x(x_56), .z(tmp00_56_12));
	booth__010 #(.WIDTH(WIDTH)) mul00120057(.x(x_57), .z(tmp00_57_12));
	booth__002 #(.WIDTH(WIDTH)) mul00120058(.x(x_58), .z(tmp00_58_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120059(.x(x_59), .z(tmp00_59_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120060(.x(x_60), .z(tmp00_60_12));
	booth__010 #(.WIDTH(WIDTH)) mul00120061(.x(x_61), .z(tmp00_61_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120062(.x(x_62), .z(tmp00_62_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120063(.x(x_63), .z(tmp00_63_12));
	booth_0012 #(.WIDTH(WIDTH)) mul00120064(.x(x_64), .z(tmp00_64_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120065(.x(x_65), .z(tmp00_65_12));
	booth__006 #(.WIDTH(WIDTH)) mul00120066(.x(x_66), .z(tmp00_66_12));
	booth__002 #(.WIDTH(WIDTH)) mul00120067(.x(x_67), .z(tmp00_67_12));
	booth_0010 #(.WIDTH(WIDTH)) mul00120068(.x(x_68), .z(tmp00_68_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120069(.x(x_69), .z(tmp00_69_12));
	booth_0006 #(.WIDTH(WIDTH)) mul00120070(.x(x_70), .z(tmp00_70_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120071(.x(x_71), .z(tmp00_71_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120072(.x(x_72), .z(tmp00_72_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120073(.x(x_73), .z(tmp00_73_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120074(.x(x_74), .z(tmp00_74_12));
	booth_0006 #(.WIDTH(WIDTH)) mul00120075(.x(x_75), .z(tmp00_75_12));
	booth_0002 #(.WIDTH(WIDTH)) mul00120076(.x(x_76), .z(tmp00_76_12));
	booth_0008 #(.WIDTH(WIDTH)) mul00120077(.x(x_77), .z(tmp00_77_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120078(.x(x_78), .z(tmp00_78_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120079(.x(x_79), .z(tmp00_79_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120080(.x(x_80), .z(tmp00_80_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120081(.x(x_81), .z(tmp00_81_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120082(.x(x_82), .z(tmp00_82_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120083(.x(x_83), .z(tmp00_83_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120084(.x(x_84), .z(tmp00_84_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120085(.x(x_85), .z(tmp00_85_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120086(.x(x_86), .z(tmp00_86_12));
	booth__006 #(.WIDTH(WIDTH)) mul00120087(.x(x_87), .z(tmp00_87_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120088(.x(x_88), .z(tmp00_88_12));
	booth__002 #(.WIDTH(WIDTH)) mul00120089(.x(x_89), .z(tmp00_89_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120090(.x(x_90), .z(tmp00_90_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120091(.x(x_91), .z(tmp00_91_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120092(.x(x_92), .z(tmp00_92_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120093(.x(x_93), .z(tmp00_93_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120094(.x(x_94), .z(tmp00_94_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120095(.x(x_95), .z(tmp00_95_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120096(.x(x_96), .z(tmp00_96_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120097(.x(x_97), .z(tmp00_97_12));
	booth__002 #(.WIDTH(WIDTH)) mul00120098(.x(x_98), .z(tmp00_98_12));
	booth__002 #(.WIDTH(WIDTH)) mul00120099(.x(x_99), .z(tmp00_99_12));
	booth_0006 #(.WIDTH(WIDTH)) mul00120100(.x(x_100), .z(tmp00_100_12));
	booth_0012 #(.WIDTH(WIDTH)) mul00120101(.x(x_101), .z(tmp00_101_12));
	booth__012 #(.WIDTH(WIDTH)) mul00120102(.x(x_102), .z(tmp00_102_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120103(.x(x_103), .z(tmp00_103_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120104(.x(x_104), .z(tmp00_104_12));
	booth_0008 #(.WIDTH(WIDTH)) mul00120105(.x(x_105), .z(tmp00_105_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120106(.x(x_106), .z(tmp00_106_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120107(.x(x_107), .z(tmp00_107_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120108(.x(x_108), .z(tmp00_108_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120109(.x(x_109), .z(tmp00_109_12));
	booth__004 #(.WIDTH(WIDTH)) mul00120110(.x(x_110), .z(tmp00_110_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120111(.x(x_111), .z(tmp00_111_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120112(.x(x_112), .z(tmp00_112_12));
	booth__006 #(.WIDTH(WIDTH)) mul00120113(.x(x_113), .z(tmp00_113_12));
	booth__002 #(.WIDTH(WIDTH)) mul00120114(.x(x_114), .z(tmp00_114_12));
	booth_0006 #(.WIDTH(WIDTH)) mul00120115(.x(x_115), .z(tmp00_115_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120116(.x(x_116), .z(tmp00_116_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120117(.x(x_117), .z(tmp00_117_12));
	booth_0010 #(.WIDTH(WIDTH)) mul00120118(.x(x_118), .z(tmp00_118_12));
	booth__008 #(.WIDTH(WIDTH)) mul00120119(.x(x_119), .z(tmp00_119_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120120(.x(x_120), .z(tmp00_120_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120121(.x(x_121), .z(tmp00_121_12));
	booth_0006 #(.WIDTH(WIDTH)) mul00120122(.x(x_122), .z(tmp00_122_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120123(.x(x_123), .z(tmp00_123_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00120124(.x(x_124), .z(tmp00_124_12));
	booth__006 #(.WIDTH(WIDTH)) mul00120125(.x(x_125), .z(tmp00_125_12));
	booth_0006 #(.WIDTH(WIDTH)) mul00120126(.x(x_126), .z(tmp00_126_12));
	booth_0004 #(.WIDTH(WIDTH)) mul00120127(.x(x_127), .z(tmp00_127_12));
	booth_0000 #(.WIDTH(WIDTH)) mul00130000(.x(x_0), .z(tmp00_0_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130001(.x(x_1), .z(tmp00_1_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130002(.x(x_2), .z(tmp00_2_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130003(.x(x_3), .z(tmp00_3_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130004(.x(x_4), .z(tmp00_4_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130005(.x(x_5), .z(tmp00_5_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130006(.x(x_6), .z(tmp00_6_13));
	booth__006 #(.WIDTH(WIDTH)) mul00130007(.x(x_7), .z(tmp00_7_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130008(.x(x_8), .z(tmp00_8_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130009(.x(x_9), .z(tmp00_9_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130010(.x(x_10), .z(tmp00_10_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130011(.x(x_11), .z(tmp00_11_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130012(.x(x_12), .z(tmp00_12_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130013(.x(x_13), .z(tmp00_13_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130014(.x(x_14), .z(tmp00_14_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130015(.x(x_15), .z(tmp00_15_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130016(.x(x_16), .z(tmp00_16_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130017(.x(x_17), .z(tmp00_17_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130018(.x(x_18), .z(tmp00_18_13));
	booth__006 #(.WIDTH(WIDTH)) mul00130019(.x(x_19), .z(tmp00_19_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130020(.x(x_20), .z(tmp00_20_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130021(.x(x_21), .z(tmp00_21_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130022(.x(x_22), .z(tmp00_22_13));
	booth_0014 #(.WIDTH(WIDTH)) mul00130023(.x(x_23), .z(tmp00_23_13));
	booth_0010 #(.WIDTH(WIDTH)) mul00130024(.x(x_24), .z(tmp00_24_13));
	booth_0012 #(.WIDTH(WIDTH)) mul00130025(.x(x_25), .z(tmp00_25_13));
	booth_0006 #(.WIDTH(WIDTH)) mul00130026(.x(x_26), .z(tmp00_26_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130027(.x(x_27), .z(tmp00_27_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130028(.x(x_28), .z(tmp00_28_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130029(.x(x_29), .z(tmp00_29_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130030(.x(x_30), .z(tmp00_30_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130031(.x(x_31), .z(tmp00_31_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130032(.x(x_32), .z(tmp00_32_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130033(.x(x_33), .z(tmp00_33_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130034(.x(x_34), .z(tmp00_34_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130035(.x(x_35), .z(tmp00_35_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130036(.x(x_36), .z(tmp00_36_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130037(.x(x_37), .z(tmp00_37_13));
	booth__006 #(.WIDTH(WIDTH)) mul00130038(.x(x_38), .z(tmp00_38_13));
	booth__012 #(.WIDTH(WIDTH)) mul00130039(.x(x_39), .z(tmp00_39_13));
	booth_0006 #(.WIDTH(WIDTH)) mul00130040(.x(x_40), .z(tmp00_40_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130041(.x(x_41), .z(tmp00_41_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130042(.x(x_42), .z(tmp00_42_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130043(.x(x_43), .z(tmp00_43_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130044(.x(x_44), .z(tmp00_44_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130045(.x(x_45), .z(tmp00_45_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130046(.x(x_46), .z(tmp00_46_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130047(.x(x_47), .z(tmp00_47_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130048(.x(x_48), .z(tmp00_48_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130049(.x(x_49), .z(tmp00_49_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130050(.x(x_50), .z(tmp00_50_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130051(.x(x_51), .z(tmp00_51_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130052(.x(x_52), .z(tmp00_52_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130053(.x(x_53), .z(tmp00_53_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130054(.x(x_54), .z(tmp00_54_13));
	booth_0006 #(.WIDTH(WIDTH)) mul00130055(.x(x_55), .z(tmp00_55_13));
	booth_0014 #(.WIDTH(WIDTH)) mul00130056(.x(x_56), .z(tmp00_56_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130057(.x(x_57), .z(tmp00_57_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130058(.x(x_58), .z(tmp00_58_13));
	booth_0016 #(.WIDTH(WIDTH)) mul00130059(.x(x_59), .z(tmp00_59_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130060(.x(x_60), .z(tmp00_60_13));
	booth__006 #(.WIDTH(WIDTH)) mul00130061(.x(x_61), .z(tmp00_61_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130062(.x(x_62), .z(tmp00_62_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130063(.x(x_63), .z(tmp00_63_13));
	booth_0010 #(.WIDTH(WIDTH)) mul00130064(.x(x_64), .z(tmp00_64_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130065(.x(x_65), .z(tmp00_65_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130066(.x(x_66), .z(tmp00_66_13));
	booth_0010 #(.WIDTH(WIDTH)) mul00130067(.x(x_67), .z(tmp00_67_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130068(.x(x_68), .z(tmp00_68_13));
	booth_0010 #(.WIDTH(WIDTH)) mul00130069(.x(x_69), .z(tmp00_69_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130070(.x(x_70), .z(tmp00_70_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130071(.x(x_71), .z(tmp00_71_13));
	booth_0012 #(.WIDTH(WIDTH)) mul00130072(.x(x_72), .z(tmp00_72_13));
	booth_0006 #(.WIDTH(WIDTH)) mul00130073(.x(x_73), .z(tmp00_73_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130074(.x(x_74), .z(tmp00_74_13));
	booth__010 #(.WIDTH(WIDTH)) mul00130075(.x(x_75), .z(tmp00_75_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130076(.x(x_76), .z(tmp00_76_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130077(.x(x_77), .z(tmp00_77_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130078(.x(x_78), .z(tmp00_78_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130079(.x(x_79), .z(tmp00_79_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130080(.x(x_80), .z(tmp00_80_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130081(.x(x_81), .z(tmp00_81_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130082(.x(x_82), .z(tmp00_82_13));
	booth_0010 #(.WIDTH(WIDTH)) mul00130083(.x(x_83), .z(tmp00_83_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130084(.x(x_84), .z(tmp00_84_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130085(.x(x_85), .z(tmp00_85_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130086(.x(x_86), .z(tmp00_86_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130087(.x(x_87), .z(tmp00_87_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130088(.x(x_88), .z(tmp00_88_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130089(.x(x_89), .z(tmp00_89_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130090(.x(x_90), .z(tmp00_90_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130091(.x(x_91), .z(tmp00_91_13));
	booth__002 #(.WIDTH(WIDTH)) mul00130092(.x(x_92), .z(tmp00_92_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130093(.x(x_93), .z(tmp00_93_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130094(.x(x_94), .z(tmp00_94_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130095(.x(x_95), .z(tmp00_95_13));
	booth__010 #(.WIDTH(WIDTH)) mul00130096(.x(x_96), .z(tmp00_96_13));
	booth_0006 #(.WIDTH(WIDTH)) mul00130097(.x(x_97), .z(tmp00_97_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130098(.x(x_98), .z(tmp00_98_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130099(.x(x_99), .z(tmp00_99_13));
	booth_0012 #(.WIDTH(WIDTH)) mul00130100(.x(x_100), .z(tmp00_100_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130101(.x(x_101), .z(tmp00_101_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130102(.x(x_102), .z(tmp00_102_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130103(.x(x_103), .z(tmp00_103_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130104(.x(x_104), .z(tmp00_104_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130105(.x(x_105), .z(tmp00_105_13));
	booth__010 #(.WIDTH(WIDTH)) mul00130106(.x(x_106), .z(tmp00_106_13));
	booth_0004 #(.WIDTH(WIDTH)) mul00130107(.x(x_107), .z(tmp00_107_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130108(.x(x_108), .z(tmp00_108_13));
	booth__002 #(.WIDTH(WIDTH)) mul00130109(.x(x_109), .z(tmp00_109_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130110(.x(x_110), .z(tmp00_110_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130111(.x(x_111), .z(tmp00_111_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130112(.x(x_112), .z(tmp00_112_13));
	booth_0016 #(.WIDTH(WIDTH)) mul00130113(.x(x_113), .z(tmp00_113_13));
	booth_0014 #(.WIDTH(WIDTH)) mul00130114(.x(x_114), .z(tmp00_114_13));
	booth_0012 #(.WIDTH(WIDTH)) mul00130115(.x(x_115), .z(tmp00_115_13));
	booth_0002 #(.WIDTH(WIDTH)) mul00130116(.x(x_116), .z(tmp00_116_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130117(.x(x_117), .z(tmp00_117_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130118(.x(x_118), .z(tmp00_118_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130119(.x(x_119), .z(tmp00_119_13));
	booth_0016 #(.WIDTH(WIDTH)) mul00130120(.x(x_120), .z(tmp00_120_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130121(.x(x_121), .z(tmp00_121_13));
	booth_0010 #(.WIDTH(WIDTH)) mul00130122(.x(x_122), .z(tmp00_122_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130123(.x(x_123), .z(tmp00_123_13));
	booth_0008 #(.WIDTH(WIDTH)) mul00130124(.x(x_124), .z(tmp00_124_13));
	booth__008 #(.WIDTH(WIDTH)) mul00130125(.x(x_125), .z(tmp00_125_13));
	booth__004 #(.WIDTH(WIDTH)) mul00130126(.x(x_126), .z(tmp00_126_13));
	booth_0000 #(.WIDTH(WIDTH)) mul00130127(.x(x_127), .z(tmp00_127_13));
	booth__006 #(.WIDTH(WIDTH)) mul00140000(.x(x_0), .z(tmp00_0_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140001(.x(x_1), .z(tmp00_1_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140002(.x(x_2), .z(tmp00_2_14));
	booth_0006 #(.WIDTH(WIDTH)) mul00140003(.x(x_3), .z(tmp00_3_14));
	booth_0010 #(.WIDTH(WIDTH)) mul00140004(.x(x_4), .z(tmp00_4_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140005(.x(x_5), .z(tmp00_5_14));
	booth_0012 #(.WIDTH(WIDTH)) mul00140006(.x(x_6), .z(tmp00_6_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140007(.x(x_7), .z(tmp00_7_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140008(.x(x_8), .z(tmp00_8_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140009(.x(x_9), .z(tmp00_9_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140010(.x(x_10), .z(tmp00_10_14));
	booth_0002 #(.WIDTH(WIDTH)) mul00140011(.x(x_11), .z(tmp00_11_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140012(.x(x_12), .z(tmp00_12_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140013(.x(x_13), .z(tmp00_13_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140014(.x(x_14), .z(tmp00_14_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140015(.x(x_15), .z(tmp00_15_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140016(.x(x_16), .z(tmp00_16_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140017(.x(x_17), .z(tmp00_17_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140018(.x(x_18), .z(tmp00_18_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140019(.x(x_19), .z(tmp00_19_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140020(.x(x_20), .z(tmp00_20_14));
	booth__010 #(.WIDTH(WIDTH)) mul00140021(.x(x_21), .z(tmp00_21_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140022(.x(x_22), .z(tmp00_22_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140023(.x(x_23), .z(tmp00_23_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140024(.x(x_24), .z(tmp00_24_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140025(.x(x_25), .z(tmp00_25_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140026(.x(x_26), .z(tmp00_26_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140027(.x(x_27), .z(tmp00_27_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140028(.x(x_28), .z(tmp00_28_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140029(.x(x_29), .z(tmp00_29_14));
	booth__010 #(.WIDTH(WIDTH)) mul00140030(.x(x_30), .z(tmp00_30_14));
	booth_0006 #(.WIDTH(WIDTH)) mul00140031(.x(x_31), .z(tmp00_31_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140032(.x(x_32), .z(tmp00_32_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140033(.x(x_33), .z(tmp00_33_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140034(.x(x_34), .z(tmp00_34_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140035(.x(x_35), .z(tmp00_35_14));
	booth_0012 #(.WIDTH(WIDTH)) mul00140036(.x(x_36), .z(tmp00_36_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140037(.x(x_37), .z(tmp00_37_14));
	booth_0010 #(.WIDTH(WIDTH)) mul00140038(.x(x_38), .z(tmp00_38_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140039(.x(x_39), .z(tmp00_39_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140040(.x(x_40), .z(tmp00_40_14));
	booth_0012 #(.WIDTH(WIDTH)) mul00140041(.x(x_41), .z(tmp00_41_14));
	booth_0016 #(.WIDTH(WIDTH)) mul00140042(.x(x_42), .z(tmp00_42_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140043(.x(x_43), .z(tmp00_43_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140044(.x(x_44), .z(tmp00_44_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140045(.x(x_45), .z(tmp00_45_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140046(.x(x_46), .z(tmp00_46_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140047(.x(x_47), .z(tmp00_47_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140048(.x(x_48), .z(tmp00_48_14));
	booth_0006 #(.WIDTH(WIDTH)) mul00140049(.x(x_49), .z(tmp00_49_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140050(.x(x_50), .z(tmp00_50_14));
	booth__006 #(.WIDTH(WIDTH)) mul00140051(.x(x_51), .z(tmp00_51_14));
	booth_0002 #(.WIDTH(WIDTH)) mul00140052(.x(x_52), .z(tmp00_52_14));
	booth__012 #(.WIDTH(WIDTH)) mul00140053(.x(x_53), .z(tmp00_53_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140054(.x(x_54), .z(tmp00_54_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140055(.x(x_55), .z(tmp00_55_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140056(.x(x_56), .z(tmp00_56_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140057(.x(x_57), .z(tmp00_57_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140058(.x(x_58), .z(tmp00_58_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140059(.x(x_59), .z(tmp00_59_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140060(.x(x_60), .z(tmp00_60_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140061(.x(x_61), .z(tmp00_61_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140062(.x(x_62), .z(tmp00_62_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140063(.x(x_63), .z(tmp00_63_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140064(.x(x_64), .z(tmp00_64_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140065(.x(x_65), .z(tmp00_65_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140066(.x(x_66), .z(tmp00_66_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140067(.x(x_67), .z(tmp00_67_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140068(.x(x_68), .z(tmp00_68_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140069(.x(x_69), .z(tmp00_69_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140070(.x(x_70), .z(tmp00_70_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140071(.x(x_71), .z(tmp00_71_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140072(.x(x_72), .z(tmp00_72_14));
	booth_0010 #(.WIDTH(WIDTH)) mul00140073(.x(x_73), .z(tmp00_73_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140074(.x(x_74), .z(tmp00_74_14));
	booth__012 #(.WIDTH(WIDTH)) mul00140075(.x(x_75), .z(tmp00_75_14));
	booth_0006 #(.WIDTH(WIDTH)) mul00140076(.x(x_76), .z(tmp00_76_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140077(.x(x_77), .z(tmp00_77_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140078(.x(x_78), .z(tmp00_78_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140079(.x(x_79), .z(tmp00_79_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140080(.x(x_80), .z(tmp00_80_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140081(.x(x_81), .z(tmp00_81_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140082(.x(x_82), .z(tmp00_82_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140083(.x(x_83), .z(tmp00_83_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140084(.x(x_84), .z(tmp00_84_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140085(.x(x_85), .z(tmp00_85_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140086(.x(x_86), .z(tmp00_86_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140087(.x(x_87), .z(tmp00_87_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140088(.x(x_88), .z(tmp00_88_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140089(.x(x_89), .z(tmp00_89_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140090(.x(x_90), .z(tmp00_90_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140091(.x(x_91), .z(tmp00_91_14));
	booth__012 #(.WIDTH(WIDTH)) mul00140092(.x(x_92), .z(tmp00_92_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140093(.x(x_93), .z(tmp00_93_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140094(.x(x_94), .z(tmp00_94_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140095(.x(x_95), .z(tmp00_95_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140096(.x(x_96), .z(tmp00_96_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140097(.x(x_97), .z(tmp00_97_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140098(.x(x_98), .z(tmp00_98_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140099(.x(x_99), .z(tmp00_99_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140100(.x(x_100), .z(tmp00_100_14));
	booth__010 #(.WIDTH(WIDTH)) mul00140101(.x(x_101), .z(tmp00_101_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140102(.x(x_102), .z(tmp00_102_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140103(.x(x_103), .z(tmp00_103_14));
	booth_0002 #(.WIDTH(WIDTH)) mul00140104(.x(x_104), .z(tmp00_104_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140105(.x(x_105), .z(tmp00_105_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140106(.x(x_106), .z(tmp00_106_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140107(.x(x_107), .z(tmp00_107_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140108(.x(x_108), .z(tmp00_108_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140109(.x(x_109), .z(tmp00_109_14));
	booth_0010 #(.WIDTH(WIDTH)) mul00140110(.x(x_110), .z(tmp00_110_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140111(.x(x_111), .z(tmp00_111_14));
	booth_0006 #(.WIDTH(WIDTH)) mul00140112(.x(x_112), .z(tmp00_112_14));
	booth_0012 #(.WIDTH(WIDTH)) mul00140113(.x(x_113), .z(tmp00_113_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140114(.x(x_114), .z(tmp00_114_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140115(.x(x_115), .z(tmp00_115_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140116(.x(x_116), .z(tmp00_116_14));
	booth__004 #(.WIDTH(WIDTH)) mul00140117(.x(x_117), .z(tmp00_117_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140118(.x(x_118), .z(tmp00_118_14));
	booth_0004 #(.WIDTH(WIDTH)) mul00140119(.x(x_119), .z(tmp00_119_14));
	booth__008 #(.WIDTH(WIDTH)) mul00140120(.x(x_120), .z(tmp00_120_14));
	booth_0008 #(.WIDTH(WIDTH)) mul00140121(.x(x_121), .z(tmp00_121_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140122(.x(x_122), .z(tmp00_122_14));
	booth_0010 #(.WIDTH(WIDTH)) mul00140123(.x(x_123), .z(tmp00_123_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140124(.x(x_124), .z(tmp00_124_14));
	booth__006 #(.WIDTH(WIDTH)) mul00140125(.x(x_125), .z(tmp00_125_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140126(.x(x_126), .z(tmp00_126_14));
	booth_0000 #(.WIDTH(WIDTH)) mul00140127(.x(x_127), .z(tmp00_127_14));
	booth__006 #(.WIDTH(WIDTH)) mul00150000(.x(x_0), .z(tmp00_0_15));
	booth__006 #(.WIDTH(WIDTH)) mul00150001(.x(x_1), .z(tmp00_1_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150002(.x(x_2), .z(tmp00_2_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150003(.x(x_3), .z(tmp00_3_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150004(.x(x_4), .z(tmp00_4_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150005(.x(x_5), .z(tmp00_5_15));
	booth__012 #(.WIDTH(WIDTH)) mul00150006(.x(x_6), .z(tmp00_6_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150007(.x(x_7), .z(tmp00_7_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150008(.x(x_8), .z(tmp00_8_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150009(.x(x_9), .z(tmp00_9_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150010(.x(x_10), .z(tmp00_10_15));
	booth_0006 #(.WIDTH(WIDTH)) mul00150011(.x(x_11), .z(tmp00_11_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150012(.x(x_12), .z(tmp00_12_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150013(.x(x_13), .z(tmp00_13_15));
	booth__006 #(.WIDTH(WIDTH)) mul00150014(.x(x_14), .z(tmp00_14_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150015(.x(x_15), .z(tmp00_15_15));
	booth__002 #(.WIDTH(WIDTH)) mul00150016(.x(x_16), .z(tmp00_16_15));
	booth_0010 #(.WIDTH(WIDTH)) mul00150017(.x(x_17), .z(tmp00_17_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150018(.x(x_18), .z(tmp00_18_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150019(.x(x_19), .z(tmp00_19_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150020(.x(x_20), .z(tmp00_20_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150021(.x(x_21), .z(tmp00_21_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150022(.x(x_22), .z(tmp00_22_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150023(.x(x_23), .z(tmp00_23_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150024(.x(x_24), .z(tmp00_24_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150025(.x(x_25), .z(tmp00_25_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150026(.x(x_26), .z(tmp00_26_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150027(.x(x_27), .z(tmp00_27_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150028(.x(x_28), .z(tmp00_28_15));
	booth_0006 #(.WIDTH(WIDTH)) mul00150029(.x(x_29), .z(tmp00_29_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150030(.x(x_30), .z(tmp00_30_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150031(.x(x_31), .z(tmp00_31_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150032(.x(x_32), .z(tmp00_32_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150033(.x(x_33), .z(tmp00_33_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150034(.x(x_34), .z(tmp00_34_15));
	booth__002 #(.WIDTH(WIDTH)) mul00150035(.x(x_35), .z(tmp00_35_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150036(.x(x_36), .z(tmp00_36_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150037(.x(x_37), .z(tmp00_37_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150038(.x(x_38), .z(tmp00_38_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150039(.x(x_39), .z(tmp00_39_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150040(.x(x_40), .z(tmp00_40_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150041(.x(x_41), .z(tmp00_41_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150042(.x(x_42), .z(tmp00_42_15));
	booth_0010 #(.WIDTH(WIDTH)) mul00150043(.x(x_43), .z(tmp00_43_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150044(.x(x_44), .z(tmp00_44_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150045(.x(x_45), .z(tmp00_45_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150046(.x(x_46), .z(tmp00_46_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150047(.x(x_47), .z(tmp00_47_15));
	booth_0010 #(.WIDTH(WIDTH)) mul00150048(.x(x_48), .z(tmp00_48_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150049(.x(x_49), .z(tmp00_49_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150050(.x(x_50), .z(tmp00_50_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150051(.x(x_51), .z(tmp00_51_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150052(.x(x_52), .z(tmp00_52_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150053(.x(x_53), .z(tmp00_53_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150054(.x(x_54), .z(tmp00_54_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150055(.x(x_55), .z(tmp00_55_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150056(.x(x_56), .z(tmp00_56_15));
	booth_0010 #(.WIDTH(WIDTH)) mul00150057(.x(x_57), .z(tmp00_57_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150058(.x(x_58), .z(tmp00_58_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150059(.x(x_59), .z(tmp00_59_15));
	booth__002 #(.WIDTH(WIDTH)) mul00150060(.x(x_60), .z(tmp00_60_15));
	booth_0010 #(.WIDTH(WIDTH)) mul00150061(.x(x_61), .z(tmp00_61_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150062(.x(x_62), .z(tmp00_62_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150063(.x(x_63), .z(tmp00_63_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150064(.x(x_64), .z(tmp00_64_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150065(.x(x_65), .z(tmp00_65_15));
	booth_0010 #(.WIDTH(WIDTH)) mul00150066(.x(x_66), .z(tmp00_66_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150067(.x(x_67), .z(tmp00_67_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150068(.x(x_68), .z(tmp00_68_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150069(.x(x_69), .z(tmp00_69_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150070(.x(x_70), .z(tmp00_70_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150071(.x(x_71), .z(tmp00_71_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150072(.x(x_72), .z(tmp00_72_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150073(.x(x_73), .z(tmp00_73_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150074(.x(x_74), .z(tmp00_74_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150075(.x(x_75), .z(tmp00_75_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150076(.x(x_76), .z(tmp00_76_15));
	booth__002 #(.WIDTH(WIDTH)) mul00150077(.x(x_77), .z(tmp00_77_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150078(.x(x_78), .z(tmp00_78_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150079(.x(x_79), .z(tmp00_79_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150080(.x(x_80), .z(tmp00_80_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150081(.x(x_81), .z(tmp00_81_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150082(.x(x_82), .z(tmp00_82_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150083(.x(x_83), .z(tmp00_83_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150084(.x(x_84), .z(tmp00_84_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150085(.x(x_85), .z(tmp00_85_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150086(.x(x_86), .z(tmp00_86_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150087(.x(x_87), .z(tmp00_87_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150088(.x(x_88), .z(tmp00_88_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150089(.x(x_89), .z(tmp00_89_15));
	booth__006 #(.WIDTH(WIDTH)) mul00150090(.x(x_90), .z(tmp00_90_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150091(.x(x_91), .z(tmp00_91_15));
	booth__006 #(.WIDTH(WIDTH)) mul00150092(.x(x_92), .z(tmp00_92_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150093(.x(x_93), .z(tmp00_93_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150094(.x(x_94), .z(tmp00_94_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150095(.x(x_95), .z(tmp00_95_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150096(.x(x_96), .z(tmp00_96_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150097(.x(x_97), .z(tmp00_97_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150098(.x(x_98), .z(tmp00_98_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150099(.x(x_99), .z(tmp00_99_15));
	booth__006 #(.WIDTH(WIDTH)) mul00150100(.x(x_100), .z(tmp00_100_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150101(.x(x_101), .z(tmp00_101_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150102(.x(x_102), .z(tmp00_102_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150103(.x(x_103), .z(tmp00_103_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00150104(.x(x_104), .z(tmp00_104_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150105(.x(x_105), .z(tmp00_105_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150106(.x(x_106), .z(tmp00_106_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150107(.x(x_107), .z(tmp00_107_15));
	booth__002 #(.WIDTH(WIDTH)) mul00150108(.x(x_108), .z(tmp00_108_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150109(.x(x_109), .z(tmp00_109_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150110(.x(x_110), .z(tmp00_110_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150111(.x(x_111), .z(tmp00_111_15));
	booth__010 #(.WIDTH(WIDTH)) mul00150112(.x(x_112), .z(tmp00_112_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150113(.x(x_113), .z(tmp00_113_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150114(.x(x_114), .z(tmp00_114_15));
	booth__002 #(.WIDTH(WIDTH)) mul00150115(.x(x_115), .z(tmp00_115_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150116(.x(x_116), .z(tmp00_116_15));
	booth__004 #(.WIDTH(WIDTH)) mul00150117(.x(x_117), .z(tmp00_117_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150118(.x(x_118), .z(tmp00_118_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150119(.x(x_119), .z(tmp00_119_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150120(.x(x_120), .z(tmp00_120_15));
	booth_0008 #(.WIDTH(WIDTH)) mul00150121(.x(x_121), .z(tmp00_121_15));
	booth_0010 #(.WIDTH(WIDTH)) mul00150122(.x(x_122), .z(tmp00_122_15));
	booth__008 #(.WIDTH(WIDTH)) mul00150123(.x(x_123), .z(tmp00_123_15));
	booth_0002 #(.WIDTH(WIDTH)) mul00150124(.x(x_124), .z(tmp00_124_15));
	booth_0000 #(.WIDTH(WIDTH)) mul00150125(.x(x_125), .z(tmp00_125_15));
	booth_0006 #(.WIDTH(WIDTH)) mul00150126(.x(x_126), .z(tmp00_126_15));
	booth__006 #(.WIDTH(WIDTH)) mul00150127(.x(x_127), .z(tmp00_127_15));
	booth_0004 #(.WIDTH(WIDTH)) mul00160000(.x(x_0), .z(tmp00_0_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160001(.x(x_1), .z(tmp00_1_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160002(.x(x_2), .z(tmp00_2_16));
	booth__006 #(.WIDTH(WIDTH)) mul00160003(.x(x_3), .z(tmp00_3_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160004(.x(x_4), .z(tmp00_4_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160005(.x(x_5), .z(tmp00_5_16));
	booth__010 #(.WIDTH(WIDTH)) mul00160006(.x(x_6), .z(tmp00_6_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160007(.x(x_7), .z(tmp00_7_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160008(.x(x_8), .z(tmp00_8_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160009(.x(x_9), .z(tmp00_9_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160010(.x(x_10), .z(tmp00_10_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160011(.x(x_11), .z(tmp00_11_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160012(.x(x_12), .z(tmp00_12_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160013(.x(x_13), .z(tmp00_13_16));
	booth_0010 #(.WIDTH(WIDTH)) mul00160014(.x(x_14), .z(tmp00_14_16));
	booth__010 #(.WIDTH(WIDTH)) mul00160015(.x(x_15), .z(tmp00_15_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160016(.x(x_16), .z(tmp00_16_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160017(.x(x_17), .z(tmp00_17_16));
	booth__006 #(.WIDTH(WIDTH)) mul00160018(.x(x_18), .z(tmp00_18_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160019(.x(x_19), .z(tmp00_19_16));
	booth_0006 #(.WIDTH(WIDTH)) mul00160020(.x(x_20), .z(tmp00_20_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160021(.x(x_21), .z(tmp00_21_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160022(.x(x_22), .z(tmp00_22_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160023(.x(x_23), .z(tmp00_23_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160024(.x(x_24), .z(tmp00_24_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160025(.x(x_25), .z(tmp00_25_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160026(.x(x_26), .z(tmp00_26_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160027(.x(x_27), .z(tmp00_27_16));
	booth_0002 #(.WIDTH(WIDTH)) mul00160028(.x(x_28), .z(tmp00_28_16));
	booth__010 #(.WIDTH(WIDTH)) mul00160029(.x(x_29), .z(tmp00_29_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160030(.x(x_30), .z(tmp00_30_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160031(.x(x_31), .z(tmp00_31_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160032(.x(x_32), .z(tmp00_32_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160033(.x(x_33), .z(tmp00_33_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160034(.x(x_34), .z(tmp00_34_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160035(.x(x_35), .z(tmp00_35_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160036(.x(x_36), .z(tmp00_36_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160037(.x(x_37), .z(tmp00_37_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160038(.x(x_38), .z(tmp00_38_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160039(.x(x_39), .z(tmp00_39_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160040(.x(x_40), .z(tmp00_40_16));
	booth_0010 #(.WIDTH(WIDTH)) mul00160041(.x(x_41), .z(tmp00_41_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160042(.x(x_42), .z(tmp00_42_16));
	booth__006 #(.WIDTH(WIDTH)) mul00160043(.x(x_43), .z(tmp00_43_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160044(.x(x_44), .z(tmp00_44_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160045(.x(x_45), .z(tmp00_45_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160046(.x(x_46), .z(tmp00_46_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160047(.x(x_47), .z(tmp00_47_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160048(.x(x_48), .z(tmp00_48_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160049(.x(x_49), .z(tmp00_49_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160050(.x(x_50), .z(tmp00_50_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160051(.x(x_51), .z(tmp00_51_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160052(.x(x_52), .z(tmp00_52_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160053(.x(x_53), .z(tmp00_53_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160054(.x(x_54), .z(tmp00_54_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160055(.x(x_55), .z(tmp00_55_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160056(.x(x_56), .z(tmp00_56_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160057(.x(x_57), .z(tmp00_57_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160058(.x(x_58), .z(tmp00_58_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160059(.x(x_59), .z(tmp00_59_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160060(.x(x_60), .z(tmp00_60_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160061(.x(x_61), .z(tmp00_61_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160062(.x(x_62), .z(tmp00_62_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160063(.x(x_63), .z(tmp00_63_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160064(.x(x_64), .z(tmp00_64_16));
	booth_0010 #(.WIDTH(WIDTH)) mul00160065(.x(x_65), .z(tmp00_65_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160066(.x(x_66), .z(tmp00_66_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160067(.x(x_67), .z(tmp00_67_16));
	booth__010 #(.WIDTH(WIDTH)) mul00160068(.x(x_68), .z(tmp00_68_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160069(.x(x_69), .z(tmp00_69_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160070(.x(x_70), .z(tmp00_70_16));
	booth_0006 #(.WIDTH(WIDTH)) mul00160071(.x(x_71), .z(tmp00_71_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160072(.x(x_72), .z(tmp00_72_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160073(.x(x_73), .z(tmp00_73_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160074(.x(x_74), .z(tmp00_74_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160075(.x(x_75), .z(tmp00_75_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160076(.x(x_76), .z(tmp00_76_16));
	booth_0010 #(.WIDTH(WIDTH)) mul00160077(.x(x_77), .z(tmp00_77_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160078(.x(x_78), .z(tmp00_78_16));
	booth_0010 #(.WIDTH(WIDTH)) mul00160079(.x(x_79), .z(tmp00_79_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160080(.x(x_80), .z(tmp00_80_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160081(.x(x_81), .z(tmp00_81_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160082(.x(x_82), .z(tmp00_82_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160083(.x(x_83), .z(tmp00_83_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160084(.x(x_84), .z(tmp00_84_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160085(.x(x_85), .z(tmp00_85_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160086(.x(x_86), .z(tmp00_86_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160087(.x(x_87), .z(tmp00_87_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160088(.x(x_88), .z(tmp00_88_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160089(.x(x_89), .z(tmp00_89_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160090(.x(x_90), .z(tmp00_90_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160091(.x(x_91), .z(tmp00_91_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160092(.x(x_92), .z(tmp00_92_16));
	booth__010 #(.WIDTH(WIDTH)) mul00160093(.x(x_93), .z(tmp00_93_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160094(.x(x_94), .z(tmp00_94_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160095(.x(x_95), .z(tmp00_95_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160096(.x(x_96), .z(tmp00_96_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160097(.x(x_97), .z(tmp00_97_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160098(.x(x_98), .z(tmp00_98_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160099(.x(x_99), .z(tmp00_99_16));
	booth_0002 #(.WIDTH(WIDTH)) mul00160100(.x(x_100), .z(tmp00_100_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160101(.x(x_101), .z(tmp00_101_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160102(.x(x_102), .z(tmp00_102_16));
	booth_0006 #(.WIDTH(WIDTH)) mul00160103(.x(x_103), .z(tmp00_103_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160104(.x(x_104), .z(tmp00_104_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160105(.x(x_105), .z(tmp00_105_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160106(.x(x_106), .z(tmp00_106_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160107(.x(x_107), .z(tmp00_107_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160108(.x(x_108), .z(tmp00_108_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160109(.x(x_109), .z(tmp00_109_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160110(.x(x_110), .z(tmp00_110_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160111(.x(x_111), .z(tmp00_111_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160112(.x(x_112), .z(tmp00_112_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160113(.x(x_113), .z(tmp00_113_16));
	booth_0006 #(.WIDTH(WIDTH)) mul00160114(.x(x_114), .z(tmp00_114_16));
	booth__008 #(.WIDTH(WIDTH)) mul00160115(.x(x_115), .z(tmp00_115_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00160116(.x(x_116), .z(tmp00_116_16));
	booth__002 #(.WIDTH(WIDTH)) mul00160117(.x(x_117), .z(tmp00_117_16));
	booth_0002 #(.WIDTH(WIDTH)) mul00160118(.x(x_118), .z(tmp00_118_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160119(.x(x_119), .z(tmp00_119_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160120(.x(x_120), .z(tmp00_120_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160121(.x(x_121), .z(tmp00_121_16));
	booth_0004 #(.WIDTH(WIDTH)) mul00160122(.x(x_122), .z(tmp00_122_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160123(.x(x_123), .z(tmp00_123_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160124(.x(x_124), .z(tmp00_124_16));
	booth__004 #(.WIDTH(WIDTH)) mul00160125(.x(x_125), .z(tmp00_125_16));
	booth_0000 #(.WIDTH(WIDTH)) mul00160126(.x(x_126), .z(tmp00_126_16));
	booth_0010 #(.WIDTH(WIDTH)) mul00160127(.x(x_127), .z(tmp00_127_16));
	booth_0008 #(.WIDTH(WIDTH)) mul00170000(.x(x_0), .z(tmp00_0_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170001(.x(x_1), .z(tmp00_1_17));
	booth__012 #(.WIDTH(WIDTH)) mul00170002(.x(x_2), .z(tmp00_2_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170003(.x(x_3), .z(tmp00_3_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170004(.x(x_4), .z(tmp00_4_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170005(.x(x_5), .z(tmp00_5_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170006(.x(x_6), .z(tmp00_6_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00170007(.x(x_7), .z(tmp00_7_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170008(.x(x_8), .z(tmp00_8_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170009(.x(x_9), .z(tmp00_9_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00170010(.x(x_10), .z(tmp00_10_17));
	booth_0002 #(.WIDTH(WIDTH)) mul00170011(.x(x_11), .z(tmp00_11_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170012(.x(x_12), .z(tmp00_12_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170013(.x(x_13), .z(tmp00_13_17));
	booth_0006 #(.WIDTH(WIDTH)) mul00170014(.x(x_14), .z(tmp00_14_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170015(.x(x_15), .z(tmp00_15_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170016(.x(x_16), .z(tmp00_16_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170017(.x(x_17), .z(tmp00_17_17));
	booth__006 #(.WIDTH(WIDTH)) mul00170018(.x(x_18), .z(tmp00_18_17));
	booth__016 #(.WIDTH(WIDTH)) mul00170019(.x(x_19), .z(tmp00_19_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170020(.x(x_20), .z(tmp00_20_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170021(.x(x_21), .z(tmp00_21_17));
	booth_0014 #(.WIDTH(WIDTH)) mul00170022(.x(x_22), .z(tmp00_22_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170023(.x(x_23), .z(tmp00_23_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170024(.x(x_24), .z(tmp00_24_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170025(.x(x_25), .z(tmp00_25_17));
	booth__010 #(.WIDTH(WIDTH)) mul00170026(.x(x_26), .z(tmp00_26_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170027(.x(x_27), .z(tmp00_27_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170028(.x(x_28), .z(tmp00_28_17));
	booth__010 #(.WIDTH(WIDTH)) mul00170029(.x(x_29), .z(tmp00_29_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00170030(.x(x_30), .z(tmp00_30_17));
	booth_0010 #(.WIDTH(WIDTH)) mul00170031(.x(x_31), .z(tmp00_31_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170032(.x(x_32), .z(tmp00_32_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00170033(.x(x_33), .z(tmp00_33_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170034(.x(x_34), .z(tmp00_34_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00170035(.x(x_35), .z(tmp00_35_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170036(.x(x_36), .z(tmp00_36_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170037(.x(x_37), .z(tmp00_37_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170038(.x(x_38), .z(tmp00_38_17));
	booth_0028 #(.WIDTH(WIDTH)) mul00170039(.x(x_39), .z(tmp00_39_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170040(.x(x_40), .z(tmp00_40_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170041(.x(x_41), .z(tmp00_41_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170042(.x(x_42), .z(tmp00_42_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170043(.x(x_43), .z(tmp00_43_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170044(.x(x_44), .z(tmp00_44_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170045(.x(x_45), .z(tmp00_45_17));
	booth__012 #(.WIDTH(WIDTH)) mul00170046(.x(x_46), .z(tmp00_46_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170047(.x(x_47), .z(tmp00_47_17));
	booth_0014 #(.WIDTH(WIDTH)) mul00170048(.x(x_48), .z(tmp00_48_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170049(.x(x_49), .z(tmp00_49_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170050(.x(x_50), .z(tmp00_50_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170051(.x(x_51), .z(tmp00_51_17));
	booth__012 #(.WIDTH(WIDTH)) mul00170052(.x(x_52), .z(tmp00_52_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170053(.x(x_53), .z(tmp00_53_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170054(.x(x_54), .z(tmp00_54_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170055(.x(x_55), .z(tmp00_55_17));
	booth__016 #(.WIDTH(WIDTH)) mul00170056(.x(x_56), .z(tmp00_56_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170057(.x(x_57), .z(tmp00_57_17));
	booth__012 #(.WIDTH(WIDTH)) mul00170058(.x(x_58), .z(tmp00_58_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170059(.x(x_59), .z(tmp00_59_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170060(.x(x_60), .z(tmp00_60_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170061(.x(x_61), .z(tmp00_61_17));
	booth__002 #(.WIDTH(WIDTH)) mul00170062(.x(x_62), .z(tmp00_62_17));
	booth__012 #(.WIDTH(WIDTH)) mul00170063(.x(x_63), .z(tmp00_63_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170064(.x(x_64), .z(tmp00_64_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170065(.x(x_65), .z(tmp00_65_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170066(.x(x_66), .z(tmp00_66_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170067(.x(x_67), .z(tmp00_67_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00170068(.x(x_68), .z(tmp00_68_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170069(.x(x_69), .z(tmp00_69_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170070(.x(x_70), .z(tmp00_70_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00170071(.x(x_71), .z(tmp00_71_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170072(.x(x_72), .z(tmp00_72_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170073(.x(x_73), .z(tmp00_73_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170074(.x(x_74), .z(tmp00_74_17));
	booth_0014 #(.WIDTH(WIDTH)) mul00170075(.x(x_75), .z(tmp00_75_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170076(.x(x_76), .z(tmp00_76_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170077(.x(x_77), .z(tmp00_77_17));
	booth_0010 #(.WIDTH(WIDTH)) mul00170078(.x(x_78), .z(tmp00_78_17));
	booth__006 #(.WIDTH(WIDTH)) mul00170079(.x(x_79), .z(tmp00_79_17));
	booth_0014 #(.WIDTH(WIDTH)) mul00170080(.x(x_80), .z(tmp00_80_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170081(.x(x_81), .z(tmp00_81_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170082(.x(x_82), .z(tmp00_82_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170083(.x(x_83), .z(tmp00_83_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170084(.x(x_84), .z(tmp00_84_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170085(.x(x_85), .z(tmp00_85_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170086(.x(x_86), .z(tmp00_86_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170087(.x(x_87), .z(tmp00_87_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170088(.x(x_88), .z(tmp00_88_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170089(.x(x_89), .z(tmp00_89_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170090(.x(x_90), .z(tmp00_90_17));
	booth_0016 #(.WIDTH(WIDTH)) mul00170091(.x(x_91), .z(tmp00_91_17));
	booth_0016 #(.WIDTH(WIDTH)) mul00170092(.x(x_92), .z(tmp00_92_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170093(.x(x_93), .z(tmp00_93_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170094(.x(x_94), .z(tmp00_94_17));
	booth_0010 #(.WIDTH(WIDTH)) mul00170095(.x(x_95), .z(tmp00_95_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170096(.x(x_96), .z(tmp00_96_17));
	booth_0006 #(.WIDTH(WIDTH)) mul00170097(.x(x_97), .z(tmp00_97_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170098(.x(x_98), .z(tmp00_98_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170099(.x(x_99), .z(tmp00_99_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170100(.x(x_100), .z(tmp00_100_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170101(.x(x_101), .z(tmp00_101_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170102(.x(x_102), .z(tmp00_102_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00170103(.x(x_103), .z(tmp00_103_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170104(.x(x_104), .z(tmp00_104_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170105(.x(x_105), .z(tmp00_105_17));
	booth__004 #(.WIDTH(WIDTH)) mul00170106(.x(x_106), .z(tmp00_106_17));
	booth_0010 #(.WIDTH(WIDTH)) mul00170107(.x(x_107), .z(tmp00_107_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170108(.x(x_108), .z(tmp00_108_17));
	booth__012 #(.WIDTH(WIDTH)) mul00170109(.x(x_109), .z(tmp00_109_17));
	booth__002 #(.WIDTH(WIDTH)) mul00170110(.x(x_110), .z(tmp00_110_17));
	booth__002 #(.WIDTH(WIDTH)) mul00170111(.x(x_111), .z(tmp00_111_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170112(.x(x_112), .z(tmp00_112_17));
	booth_0016 #(.WIDTH(WIDTH)) mul00170113(.x(x_113), .z(tmp00_113_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170114(.x(x_114), .z(tmp00_114_17));
	booth__012 #(.WIDTH(WIDTH)) mul00170115(.x(x_115), .z(tmp00_115_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170116(.x(x_116), .z(tmp00_116_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170117(.x(x_117), .z(tmp00_117_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170118(.x(x_118), .z(tmp00_118_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170119(.x(x_119), .z(tmp00_119_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170120(.x(x_120), .z(tmp00_120_17));
	booth_0004 #(.WIDTH(WIDTH)) mul00170121(.x(x_121), .z(tmp00_121_17));
	booth__008 #(.WIDTH(WIDTH)) mul00170122(.x(x_122), .z(tmp00_122_17));
	booth_0010 #(.WIDTH(WIDTH)) mul00170123(.x(x_123), .z(tmp00_123_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170124(.x(x_124), .z(tmp00_124_17));
	booth__006 #(.WIDTH(WIDTH)) mul00170125(.x(x_125), .z(tmp00_125_17));
	booth_0012 #(.WIDTH(WIDTH)) mul00170126(.x(x_126), .z(tmp00_126_17));
	booth_0000 #(.WIDTH(WIDTH)) mul00170127(.x(x_127), .z(tmp00_127_17));
	booth_0008 #(.WIDTH(WIDTH)) mul00180000(.x(x_0), .z(tmp00_0_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180001(.x(x_1), .z(tmp00_1_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180002(.x(x_2), .z(tmp00_2_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180003(.x(x_3), .z(tmp00_3_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180004(.x(x_4), .z(tmp00_4_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180005(.x(x_5), .z(tmp00_5_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180006(.x(x_6), .z(tmp00_6_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180007(.x(x_7), .z(tmp00_7_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180008(.x(x_8), .z(tmp00_8_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180009(.x(x_9), .z(tmp00_9_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180010(.x(x_10), .z(tmp00_10_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180011(.x(x_11), .z(tmp00_11_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180012(.x(x_12), .z(tmp00_12_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180013(.x(x_13), .z(tmp00_13_18));
	booth__006 #(.WIDTH(WIDTH)) mul00180014(.x(x_14), .z(tmp00_14_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180015(.x(x_15), .z(tmp00_15_18));
	booth__010 #(.WIDTH(WIDTH)) mul00180016(.x(x_16), .z(tmp00_16_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180017(.x(x_17), .z(tmp00_17_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180018(.x(x_18), .z(tmp00_18_18));
	booth__012 #(.WIDTH(WIDTH)) mul00180019(.x(x_19), .z(tmp00_19_18));
	booth__006 #(.WIDTH(WIDTH)) mul00180020(.x(x_20), .z(tmp00_20_18));
	booth__008 #(.WIDTH(WIDTH)) mul00180021(.x(x_21), .z(tmp00_21_18));
	booth__008 #(.WIDTH(WIDTH)) mul00180022(.x(x_22), .z(tmp00_22_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180023(.x(x_23), .z(tmp00_23_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180024(.x(x_24), .z(tmp00_24_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180025(.x(x_25), .z(tmp00_25_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180026(.x(x_26), .z(tmp00_26_18));
	booth__008 #(.WIDTH(WIDTH)) mul00180027(.x(x_27), .z(tmp00_27_18));
	booth_0002 #(.WIDTH(WIDTH)) mul00180028(.x(x_28), .z(tmp00_28_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180029(.x(x_29), .z(tmp00_29_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180030(.x(x_30), .z(tmp00_30_18));
	booth__006 #(.WIDTH(WIDTH)) mul00180031(.x(x_31), .z(tmp00_31_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180032(.x(x_32), .z(tmp00_32_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180033(.x(x_33), .z(tmp00_33_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180034(.x(x_34), .z(tmp00_34_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180035(.x(x_35), .z(tmp00_35_18));
	booth_0010 #(.WIDTH(WIDTH)) mul00180036(.x(x_36), .z(tmp00_36_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180037(.x(x_37), .z(tmp00_37_18));
	booth_0002 #(.WIDTH(WIDTH)) mul00180038(.x(x_38), .z(tmp00_38_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180039(.x(x_39), .z(tmp00_39_18));
	booth_0006 #(.WIDTH(WIDTH)) mul00180040(.x(x_40), .z(tmp00_40_18));
	booth_0002 #(.WIDTH(WIDTH)) mul00180041(.x(x_41), .z(tmp00_41_18));
	booth_0014 #(.WIDTH(WIDTH)) mul00180042(.x(x_42), .z(tmp00_42_18));
	booth__012 #(.WIDTH(WIDTH)) mul00180043(.x(x_43), .z(tmp00_43_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180044(.x(x_44), .z(tmp00_44_18));
	booth_0002 #(.WIDTH(WIDTH)) mul00180045(.x(x_45), .z(tmp00_45_18));
	booth__012 #(.WIDTH(WIDTH)) mul00180046(.x(x_46), .z(tmp00_46_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180047(.x(x_47), .z(tmp00_47_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180048(.x(x_48), .z(tmp00_48_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180049(.x(x_49), .z(tmp00_49_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180050(.x(x_50), .z(tmp00_50_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180051(.x(x_51), .z(tmp00_51_18));
	booth__012 #(.WIDTH(WIDTH)) mul00180052(.x(x_52), .z(tmp00_52_18));
	booth_0002 #(.WIDTH(WIDTH)) mul00180053(.x(x_53), .z(tmp00_53_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180054(.x(x_54), .z(tmp00_54_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180055(.x(x_55), .z(tmp00_55_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180056(.x(x_56), .z(tmp00_56_18));
	booth__010 #(.WIDTH(WIDTH)) mul00180057(.x(x_57), .z(tmp00_57_18));
	booth_0006 #(.WIDTH(WIDTH)) mul00180058(.x(x_58), .z(tmp00_58_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180059(.x(x_59), .z(tmp00_59_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180060(.x(x_60), .z(tmp00_60_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180061(.x(x_61), .z(tmp00_61_18));
	booth__010 #(.WIDTH(WIDTH)) mul00180062(.x(x_62), .z(tmp00_62_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180063(.x(x_63), .z(tmp00_63_18));
	booth_0006 #(.WIDTH(WIDTH)) mul00180064(.x(x_64), .z(tmp00_64_18));
	booth__008 #(.WIDTH(WIDTH)) mul00180065(.x(x_65), .z(tmp00_65_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180066(.x(x_66), .z(tmp00_66_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180067(.x(x_67), .z(tmp00_67_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180068(.x(x_68), .z(tmp00_68_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180069(.x(x_69), .z(tmp00_69_18));
	booth_0012 #(.WIDTH(WIDTH)) mul00180070(.x(x_70), .z(tmp00_70_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180071(.x(x_71), .z(tmp00_71_18));
	booth__008 #(.WIDTH(WIDTH)) mul00180072(.x(x_72), .z(tmp00_72_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180073(.x(x_73), .z(tmp00_73_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180074(.x(x_74), .z(tmp00_74_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180075(.x(x_75), .z(tmp00_75_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180076(.x(x_76), .z(tmp00_76_18));
	booth_0012 #(.WIDTH(WIDTH)) mul00180077(.x(x_77), .z(tmp00_77_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180078(.x(x_78), .z(tmp00_78_18));
	booth__008 #(.WIDTH(WIDTH)) mul00180079(.x(x_79), .z(tmp00_79_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180080(.x(x_80), .z(tmp00_80_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180081(.x(x_81), .z(tmp00_81_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180082(.x(x_82), .z(tmp00_82_18));
	booth_0010 #(.WIDTH(WIDTH)) mul00180083(.x(x_83), .z(tmp00_83_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180084(.x(x_84), .z(tmp00_84_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180085(.x(x_85), .z(tmp00_85_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180086(.x(x_86), .z(tmp00_86_18));
	booth_0012 #(.WIDTH(WIDTH)) mul00180087(.x(x_87), .z(tmp00_87_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180088(.x(x_88), .z(tmp00_88_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180089(.x(x_89), .z(tmp00_89_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180090(.x(x_90), .z(tmp00_90_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180091(.x(x_91), .z(tmp00_91_18));
	booth__006 #(.WIDTH(WIDTH)) mul00180092(.x(x_92), .z(tmp00_92_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180093(.x(x_93), .z(tmp00_93_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180094(.x(x_94), .z(tmp00_94_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180095(.x(x_95), .z(tmp00_95_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180096(.x(x_96), .z(tmp00_96_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180097(.x(x_97), .z(tmp00_97_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180098(.x(x_98), .z(tmp00_98_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180099(.x(x_99), .z(tmp00_99_18));
	booth__012 #(.WIDTH(WIDTH)) mul00180100(.x(x_100), .z(tmp00_100_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180101(.x(x_101), .z(tmp00_101_18));
	booth__012 #(.WIDTH(WIDTH)) mul00180102(.x(x_102), .z(tmp00_102_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180103(.x(x_103), .z(tmp00_103_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180104(.x(x_104), .z(tmp00_104_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180105(.x(x_105), .z(tmp00_105_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180106(.x(x_106), .z(tmp00_106_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180107(.x(x_107), .z(tmp00_107_18));
	booth_0012 #(.WIDTH(WIDTH)) mul00180108(.x(x_108), .z(tmp00_108_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180109(.x(x_109), .z(tmp00_109_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180110(.x(x_110), .z(tmp00_110_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180111(.x(x_111), .z(tmp00_111_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180112(.x(x_112), .z(tmp00_112_18));
	booth_0002 #(.WIDTH(WIDTH)) mul00180113(.x(x_113), .z(tmp00_113_18));
	booth_0002 #(.WIDTH(WIDTH)) mul00180114(.x(x_114), .z(tmp00_114_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180115(.x(x_115), .z(tmp00_115_18));
	booth__004 #(.WIDTH(WIDTH)) mul00180116(.x(x_116), .z(tmp00_116_18));
	booth_0008 #(.WIDTH(WIDTH)) mul00180117(.x(x_117), .z(tmp00_117_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180118(.x(x_118), .z(tmp00_118_18));
	booth_0002 #(.WIDTH(WIDTH)) mul00180119(.x(x_119), .z(tmp00_119_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180120(.x(x_120), .z(tmp00_120_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180121(.x(x_121), .z(tmp00_121_18));
	booth__008 #(.WIDTH(WIDTH)) mul00180122(.x(x_122), .z(tmp00_122_18));
	booth__010 #(.WIDTH(WIDTH)) mul00180123(.x(x_123), .z(tmp00_123_18));
	booth__014 #(.WIDTH(WIDTH)) mul00180124(.x(x_124), .z(tmp00_124_18));
	booth_0004 #(.WIDTH(WIDTH)) mul00180125(.x(x_125), .z(tmp00_125_18));
	booth__002 #(.WIDTH(WIDTH)) mul00180126(.x(x_126), .z(tmp00_126_18));
	booth_0000 #(.WIDTH(WIDTH)) mul00180127(.x(x_127), .z(tmp00_127_18));
	booth__010 #(.WIDTH(WIDTH)) mul00190000(.x(x_0), .z(tmp00_0_19));
	booth_0010 #(.WIDTH(WIDTH)) mul00190001(.x(x_1), .z(tmp00_1_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190002(.x(x_2), .z(tmp00_2_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190003(.x(x_3), .z(tmp00_3_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190004(.x(x_4), .z(tmp00_4_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190005(.x(x_5), .z(tmp00_5_19));
	booth_0010 #(.WIDTH(WIDTH)) mul00190006(.x(x_6), .z(tmp00_6_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190007(.x(x_7), .z(tmp00_7_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190008(.x(x_8), .z(tmp00_8_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190009(.x(x_9), .z(tmp00_9_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190010(.x(x_10), .z(tmp00_10_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190011(.x(x_11), .z(tmp00_11_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190012(.x(x_12), .z(tmp00_12_19));
	booth_0010 #(.WIDTH(WIDTH)) mul00190013(.x(x_13), .z(tmp00_13_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190014(.x(x_14), .z(tmp00_14_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190015(.x(x_15), .z(tmp00_15_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190016(.x(x_16), .z(tmp00_16_19));
	booth__002 #(.WIDTH(WIDTH)) mul00190017(.x(x_17), .z(tmp00_17_19));
	booth__010 #(.WIDTH(WIDTH)) mul00190018(.x(x_18), .z(tmp00_18_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190019(.x(x_19), .z(tmp00_19_19));
	booth_0012 #(.WIDTH(WIDTH)) mul00190020(.x(x_20), .z(tmp00_20_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190021(.x(x_21), .z(tmp00_21_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190022(.x(x_22), .z(tmp00_22_19));
	booth_0002 #(.WIDTH(WIDTH)) mul00190023(.x(x_23), .z(tmp00_23_19));
	booth__010 #(.WIDTH(WIDTH)) mul00190024(.x(x_24), .z(tmp00_24_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190025(.x(x_25), .z(tmp00_25_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190026(.x(x_26), .z(tmp00_26_19));
	booth_0010 #(.WIDTH(WIDTH)) mul00190027(.x(x_27), .z(tmp00_27_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190028(.x(x_28), .z(tmp00_28_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190029(.x(x_29), .z(tmp00_29_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190030(.x(x_30), .z(tmp00_30_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190031(.x(x_31), .z(tmp00_31_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190032(.x(x_32), .z(tmp00_32_19));
	booth__010 #(.WIDTH(WIDTH)) mul00190033(.x(x_33), .z(tmp00_33_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190034(.x(x_34), .z(tmp00_34_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190035(.x(x_35), .z(tmp00_35_19));
	booth__006 #(.WIDTH(WIDTH)) mul00190036(.x(x_36), .z(tmp00_36_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190037(.x(x_37), .z(tmp00_37_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190038(.x(x_38), .z(tmp00_38_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190039(.x(x_39), .z(tmp00_39_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190040(.x(x_40), .z(tmp00_40_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190041(.x(x_41), .z(tmp00_41_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190042(.x(x_42), .z(tmp00_42_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190043(.x(x_43), .z(tmp00_43_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190044(.x(x_44), .z(tmp00_44_19));
	booth_0002 #(.WIDTH(WIDTH)) mul00190045(.x(x_45), .z(tmp00_45_19));
	booth__002 #(.WIDTH(WIDTH)) mul00190046(.x(x_46), .z(tmp00_46_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190047(.x(x_47), .z(tmp00_47_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190048(.x(x_48), .z(tmp00_48_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190049(.x(x_49), .z(tmp00_49_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190050(.x(x_50), .z(tmp00_50_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190051(.x(x_51), .z(tmp00_51_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190052(.x(x_52), .z(tmp00_52_19));
	booth__010 #(.WIDTH(WIDTH)) mul00190053(.x(x_53), .z(tmp00_53_19));
	booth__002 #(.WIDTH(WIDTH)) mul00190054(.x(x_54), .z(tmp00_54_19));
	booth_0002 #(.WIDTH(WIDTH)) mul00190055(.x(x_55), .z(tmp00_55_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190056(.x(x_56), .z(tmp00_56_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190057(.x(x_57), .z(tmp00_57_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190058(.x(x_58), .z(tmp00_58_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190059(.x(x_59), .z(tmp00_59_19));
	booth__006 #(.WIDTH(WIDTH)) mul00190060(.x(x_60), .z(tmp00_60_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190061(.x(x_61), .z(tmp00_61_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190062(.x(x_62), .z(tmp00_62_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190063(.x(x_63), .z(tmp00_63_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190064(.x(x_64), .z(tmp00_64_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190065(.x(x_65), .z(tmp00_65_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190066(.x(x_66), .z(tmp00_66_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190067(.x(x_67), .z(tmp00_67_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190068(.x(x_68), .z(tmp00_68_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190069(.x(x_69), .z(tmp00_69_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190070(.x(x_70), .z(tmp00_70_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190071(.x(x_71), .z(tmp00_71_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190072(.x(x_72), .z(tmp00_72_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190073(.x(x_73), .z(tmp00_73_19));
	booth__004 #(.WIDTH(WIDTH)) mul00190074(.x(x_74), .z(tmp00_74_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190075(.x(x_75), .z(tmp00_75_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190076(.x(x_76), .z(tmp00_76_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190077(.x(x_77), .z(tmp00_77_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190078(.x(x_78), .z(tmp00_78_19));
	booth__006 #(.WIDTH(WIDTH)) mul00190079(.x(x_79), .z(tmp00_79_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190080(.x(x_80), .z(tmp00_80_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190081(.x(x_81), .z(tmp00_81_19));
	booth_0002 #(.WIDTH(WIDTH)) mul00190082(.x(x_82), .z(tmp00_82_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190083(.x(x_83), .z(tmp00_83_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190084(.x(x_84), .z(tmp00_84_19));
	booth__006 #(.WIDTH(WIDTH)) mul00190085(.x(x_85), .z(tmp00_85_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190086(.x(x_86), .z(tmp00_86_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190087(.x(x_87), .z(tmp00_87_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190088(.x(x_88), .z(tmp00_88_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190089(.x(x_89), .z(tmp00_89_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190090(.x(x_90), .z(tmp00_90_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190091(.x(x_91), .z(tmp00_91_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190092(.x(x_92), .z(tmp00_92_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190093(.x(x_93), .z(tmp00_93_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190094(.x(x_94), .z(tmp00_94_19));
	booth_0002 #(.WIDTH(WIDTH)) mul00190095(.x(x_95), .z(tmp00_95_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190096(.x(x_96), .z(tmp00_96_19));
	booth_0010 #(.WIDTH(WIDTH)) mul00190097(.x(x_97), .z(tmp00_97_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190098(.x(x_98), .z(tmp00_98_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190099(.x(x_99), .z(tmp00_99_19));
	booth_0002 #(.WIDTH(WIDTH)) mul00190100(.x(x_100), .z(tmp00_100_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190101(.x(x_101), .z(tmp00_101_19));
	booth__002 #(.WIDTH(WIDTH)) mul00190102(.x(x_102), .z(tmp00_102_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190103(.x(x_103), .z(tmp00_103_19));
	booth_0010 #(.WIDTH(WIDTH)) mul00190104(.x(x_104), .z(tmp00_104_19));
	booth_0010 #(.WIDTH(WIDTH)) mul00190105(.x(x_105), .z(tmp00_105_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190106(.x(x_106), .z(tmp00_106_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190107(.x(x_107), .z(tmp00_107_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190108(.x(x_108), .z(tmp00_108_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190109(.x(x_109), .z(tmp00_109_19));
	booth__012 #(.WIDTH(WIDTH)) mul00190110(.x(x_110), .z(tmp00_110_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190111(.x(x_111), .z(tmp00_111_19));
	booth_0002 #(.WIDTH(WIDTH)) mul00190112(.x(x_112), .z(tmp00_112_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190113(.x(x_113), .z(tmp00_113_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190114(.x(x_114), .z(tmp00_114_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190115(.x(x_115), .z(tmp00_115_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190116(.x(x_116), .z(tmp00_116_19));
	booth_0000 #(.WIDTH(WIDTH)) mul00190117(.x(x_117), .z(tmp00_117_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00190118(.x(x_118), .z(tmp00_118_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190119(.x(x_119), .z(tmp00_119_19));
	booth__002 #(.WIDTH(WIDTH)) mul00190120(.x(x_120), .z(tmp00_120_19));
	booth_0004 #(.WIDTH(WIDTH)) mul00190121(.x(x_121), .z(tmp00_121_19));
	booth_0010 #(.WIDTH(WIDTH)) mul00190122(.x(x_122), .z(tmp00_122_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190123(.x(x_123), .z(tmp00_123_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190124(.x(x_124), .z(tmp00_124_19));
	booth_0008 #(.WIDTH(WIDTH)) mul00190125(.x(x_125), .z(tmp00_125_19));
	booth__006 #(.WIDTH(WIDTH)) mul00190126(.x(x_126), .z(tmp00_126_19));
	booth__008 #(.WIDTH(WIDTH)) mul00190127(.x(x_127), .z(tmp00_127_19));
	booth_0006 #(.WIDTH(WIDTH)) mul00200000(.x(x_0), .z(tmp00_0_20));
	booth_0004 #(.WIDTH(WIDTH)) mul00200001(.x(x_1), .z(tmp00_1_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200002(.x(x_2), .z(tmp00_2_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200003(.x(x_3), .z(tmp00_3_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200004(.x(x_4), .z(tmp00_4_20));
	booth_0006 #(.WIDTH(WIDTH)) mul00200005(.x(x_5), .z(tmp00_5_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200006(.x(x_6), .z(tmp00_6_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200007(.x(x_7), .z(tmp00_7_20));
	booth__006 #(.WIDTH(WIDTH)) mul00200008(.x(x_8), .z(tmp00_8_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200009(.x(x_9), .z(tmp00_9_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200010(.x(x_10), .z(tmp00_10_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200011(.x(x_11), .z(tmp00_11_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200012(.x(x_12), .z(tmp00_12_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200013(.x(x_13), .z(tmp00_13_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200014(.x(x_14), .z(tmp00_14_20));
	booth_0006 #(.WIDTH(WIDTH)) mul00200015(.x(x_15), .z(tmp00_15_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200016(.x(x_16), .z(tmp00_16_20));
	booth_0004 #(.WIDTH(WIDTH)) mul00200017(.x(x_17), .z(tmp00_17_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200018(.x(x_18), .z(tmp00_18_20));
	booth_0016 #(.WIDTH(WIDTH)) mul00200019(.x(x_19), .z(tmp00_19_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200020(.x(x_20), .z(tmp00_20_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200021(.x(x_21), .z(tmp00_21_20));
	booth_0002 #(.WIDTH(WIDTH)) mul00200022(.x(x_22), .z(tmp00_22_20));
	booth_0016 #(.WIDTH(WIDTH)) mul00200023(.x(x_23), .z(tmp00_23_20));
	booth_0020 #(.WIDTH(WIDTH)) mul00200024(.x(x_24), .z(tmp00_24_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200025(.x(x_25), .z(tmp00_25_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200026(.x(x_26), .z(tmp00_26_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200027(.x(x_27), .z(tmp00_27_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200028(.x(x_28), .z(tmp00_28_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200029(.x(x_29), .z(tmp00_29_20));
	booth__002 #(.WIDTH(WIDTH)) mul00200030(.x(x_30), .z(tmp00_30_20));
	booth_0004 #(.WIDTH(WIDTH)) mul00200031(.x(x_31), .z(tmp00_31_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200032(.x(x_32), .z(tmp00_32_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200033(.x(x_33), .z(tmp00_33_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200034(.x(x_34), .z(tmp00_34_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200035(.x(x_35), .z(tmp00_35_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200036(.x(x_36), .z(tmp00_36_20));
	booth_0012 #(.WIDTH(WIDTH)) mul00200037(.x(x_37), .z(tmp00_37_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200038(.x(x_38), .z(tmp00_38_20));
	booth__022 #(.WIDTH(WIDTH)) mul00200039(.x(x_39), .z(tmp00_39_20));
	booth_0010 #(.WIDTH(WIDTH)) mul00200040(.x(x_40), .z(tmp00_40_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200041(.x(x_41), .z(tmp00_41_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200042(.x(x_42), .z(tmp00_42_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200043(.x(x_43), .z(tmp00_43_20));
	booth__016 #(.WIDTH(WIDTH)) mul00200044(.x(x_44), .z(tmp00_44_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200045(.x(x_45), .z(tmp00_45_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200046(.x(x_46), .z(tmp00_46_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200047(.x(x_47), .z(tmp00_47_20));
	booth__002 #(.WIDTH(WIDTH)) mul00200048(.x(x_48), .z(tmp00_48_20));
	booth_0004 #(.WIDTH(WIDTH)) mul00200049(.x(x_49), .z(tmp00_49_20));
	booth_0006 #(.WIDTH(WIDTH)) mul00200050(.x(x_50), .z(tmp00_50_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200051(.x(x_51), .z(tmp00_51_20));
	booth_0012 #(.WIDTH(WIDTH)) mul00200052(.x(x_52), .z(tmp00_52_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200053(.x(x_53), .z(tmp00_53_20));
	booth__012 #(.WIDTH(WIDTH)) mul00200054(.x(x_54), .z(tmp00_54_20));
	booth_0016 #(.WIDTH(WIDTH)) mul00200055(.x(x_55), .z(tmp00_55_20));
	booth_0016 #(.WIDTH(WIDTH)) mul00200056(.x(x_56), .z(tmp00_56_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200057(.x(x_57), .z(tmp00_57_20));
	booth_0012 #(.WIDTH(WIDTH)) mul00200058(.x(x_58), .z(tmp00_58_20));
	booth_0020 #(.WIDTH(WIDTH)) mul00200059(.x(x_59), .z(tmp00_59_20));
	booth_0010 #(.WIDTH(WIDTH)) mul00200060(.x(x_60), .z(tmp00_60_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200061(.x(x_61), .z(tmp00_61_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200062(.x(x_62), .z(tmp00_62_20));
	booth_0014 #(.WIDTH(WIDTH)) mul00200063(.x(x_63), .z(tmp00_63_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200064(.x(x_64), .z(tmp00_64_20));
	booth_0004 #(.WIDTH(WIDTH)) mul00200065(.x(x_65), .z(tmp00_65_20));
	booth_0014 #(.WIDTH(WIDTH)) mul00200066(.x(x_66), .z(tmp00_66_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200067(.x(x_67), .z(tmp00_67_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200068(.x(x_68), .z(tmp00_68_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200069(.x(x_69), .z(tmp00_69_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200070(.x(x_70), .z(tmp00_70_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200071(.x(x_71), .z(tmp00_71_20));
	booth_0012 #(.WIDTH(WIDTH)) mul00200072(.x(x_72), .z(tmp00_72_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200073(.x(x_73), .z(tmp00_73_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200074(.x(x_74), .z(tmp00_74_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200075(.x(x_75), .z(tmp00_75_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200076(.x(x_76), .z(tmp00_76_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200077(.x(x_77), .z(tmp00_77_20));
	booth_0002 #(.WIDTH(WIDTH)) mul00200078(.x(x_78), .z(tmp00_78_20));
	booth_0010 #(.WIDTH(WIDTH)) mul00200079(.x(x_79), .z(tmp00_79_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200080(.x(x_80), .z(tmp00_80_20));
	booth_0016 #(.WIDTH(WIDTH)) mul00200081(.x(x_81), .z(tmp00_81_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200082(.x(x_82), .z(tmp00_82_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200083(.x(x_83), .z(tmp00_83_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200084(.x(x_84), .z(tmp00_84_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200085(.x(x_85), .z(tmp00_85_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200086(.x(x_86), .z(tmp00_86_20));
	booth__010 #(.WIDTH(WIDTH)) mul00200087(.x(x_87), .z(tmp00_87_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200088(.x(x_88), .z(tmp00_88_20));
	booth_0006 #(.WIDTH(WIDTH)) mul00200089(.x(x_89), .z(tmp00_89_20));
	booth__012 #(.WIDTH(WIDTH)) mul00200090(.x(x_90), .z(tmp00_90_20));
	booth_0002 #(.WIDTH(WIDTH)) mul00200091(.x(x_91), .z(tmp00_91_20));
	booth__012 #(.WIDTH(WIDTH)) mul00200092(.x(x_92), .z(tmp00_92_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200093(.x(x_93), .z(tmp00_93_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200094(.x(x_94), .z(tmp00_94_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200095(.x(x_95), .z(tmp00_95_20));
	booth__006 #(.WIDTH(WIDTH)) mul00200096(.x(x_96), .z(tmp00_96_20));
	booth__012 #(.WIDTH(WIDTH)) mul00200097(.x(x_97), .z(tmp00_97_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200098(.x(x_98), .z(tmp00_98_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200099(.x(x_99), .z(tmp00_99_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200100(.x(x_100), .z(tmp00_100_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200101(.x(x_101), .z(tmp00_101_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200102(.x(x_102), .z(tmp00_102_20));
	booth_0010 #(.WIDTH(WIDTH)) mul00200103(.x(x_103), .z(tmp00_103_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200104(.x(x_104), .z(tmp00_104_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200105(.x(x_105), .z(tmp00_105_20));
	booth__002 #(.WIDTH(WIDTH)) mul00200106(.x(x_106), .z(tmp00_106_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200107(.x(x_107), .z(tmp00_107_20));
	booth__002 #(.WIDTH(WIDTH)) mul00200108(.x(x_108), .z(tmp00_108_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200109(.x(x_109), .z(tmp00_109_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200110(.x(x_110), .z(tmp00_110_20));
	booth_0002 #(.WIDTH(WIDTH)) mul00200111(.x(x_111), .z(tmp00_111_20));
	booth__016 #(.WIDTH(WIDTH)) mul00200112(.x(x_112), .z(tmp00_112_20));
	booth_0018 #(.WIDTH(WIDTH)) mul00200113(.x(x_113), .z(tmp00_113_20));
	booth_0006 #(.WIDTH(WIDTH)) mul00200114(.x(x_114), .z(tmp00_114_20));
	booth_0016 #(.WIDTH(WIDTH)) mul00200115(.x(x_115), .z(tmp00_115_20));
	booth__002 #(.WIDTH(WIDTH)) mul00200116(.x(x_116), .z(tmp00_116_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200117(.x(x_117), .z(tmp00_117_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200118(.x(x_118), .z(tmp00_118_20));
	booth__008 #(.WIDTH(WIDTH)) mul00200119(.x(x_119), .z(tmp00_119_20));
	booth_0016 #(.WIDTH(WIDTH)) mul00200120(.x(x_120), .z(tmp00_120_20));
	booth_0014 #(.WIDTH(WIDTH)) mul00200121(.x(x_121), .z(tmp00_121_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200122(.x(x_122), .z(tmp00_122_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200123(.x(x_123), .z(tmp00_123_20));
	booth_0008 #(.WIDTH(WIDTH)) mul00200124(.x(x_124), .z(tmp00_124_20));
	booth__004 #(.WIDTH(WIDTH)) mul00200125(.x(x_125), .z(tmp00_125_20));
	booth_0000 #(.WIDTH(WIDTH)) mul00200126(.x(x_126), .z(tmp00_126_20));
	booth__002 #(.WIDTH(WIDTH)) mul00200127(.x(x_127), .z(tmp00_127_20));
	booth_0004 #(.WIDTH(WIDTH)) mul00210000(.x(x_0), .z(tmp00_0_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210001(.x(x_1), .z(tmp00_1_21));
	booth_0010 #(.WIDTH(WIDTH)) mul00210002(.x(x_2), .z(tmp00_2_21));
	booth_0010 #(.WIDTH(WIDTH)) mul00210003(.x(x_3), .z(tmp00_3_21));
	booth__006 #(.WIDTH(WIDTH)) mul00210004(.x(x_4), .z(tmp00_4_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210005(.x(x_5), .z(tmp00_5_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210006(.x(x_6), .z(tmp00_6_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210007(.x(x_7), .z(tmp00_7_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210008(.x(x_8), .z(tmp00_8_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210009(.x(x_9), .z(tmp00_9_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210010(.x(x_10), .z(tmp00_10_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210011(.x(x_11), .z(tmp00_11_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210012(.x(x_12), .z(tmp00_12_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210013(.x(x_13), .z(tmp00_13_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210014(.x(x_14), .z(tmp00_14_21));
	booth_0010 #(.WIDTH(WIDTH)) mul00210015(.x(x_15), .z(tmp00_15_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210016(.x(x_16), .z(tmp00_16_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210017(.x(x_17), .z(tmp00_17_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210018(.x(x_18), .z(tmp00_18_21));
	booth_0010 #(.WIDTH(WIDTH)) mul00210019(.x(x_19), .z(tmp00_19_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210020(.x(x_20), .z(tmp00_20_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210021(.x(x_21), .z(tmp00_21_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210022(.x(x_22), .z(tmp00_22_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210023(.x(x_23), .z(tmp00_23_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210024(.x(x_24), .z(tmp00_24_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210025(.x(x_25), .z(tmp00_25_21));
	booth_0002 #(.WIDTH(WIDTH)) mul00210026(.x(x_26), .z(tmp00_26_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210027(.x(x_27), .z(tmp00_27_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210028(.x(x_28), .z(tmp00_28_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210029(.x(x_29), .z(tmp00_29_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210030(.x(x_30), .z(tmp00_30_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210031(.x(x_31), .z(tmp00_31_21));
	booth__006 #(.WIDTH(WIDTH)) mul00210032(.x(x_32), .z(tmp00_32_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210033(.x(x_33), .z(tmp00_33_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210034(.x(x_34), .z(tmp00_34_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210035(.x(x_35), .z(tmp00_35_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210036(.x(x_36), .z(tmp00_36_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210037(.x(x_37), .z(tmp00_37_21));
	booth_0006 #(.WIDTH(WIDTH)) mul00210038(.x(x_38), .z(tmp00_38_21));
	booth__006 #(.WIDTH(WIDTH)) mul00210039(.x(x_39), .z(tmp00_39_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210040(.x(x_40), .z(tmp00_40_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210041(.x(x_41), .z(tmp00_41_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210042(.x(x_42), .z(tmp00_42_21));
	booth__006 #(.WIDTH(WIDTH)) mul00210043(.x(x_43), .z(tmp00_43_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210044(.x(x_44), .z(tmp00_44_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210045(.x(x_45), .z(tmp00_45_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210046(.x(x_46), .z(tmp00_46_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210047(.x(x_47), .z(tmp00_47_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210048(.x(x_48), .z(tmp00_48_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210049(.x(x_49), .z(tmp00_49_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210050(.x(x_50), .z(tmp00_50_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210051(.x(x_51), .z(tmp00_51_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210052(.x(x_52), .z(tmp00_52_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210053(.x(x_53), .z(tmp00_53_21));
	booth__010 #(.WIDTH(WIDTH)) mul00210054(.x(x_54), .z(tmp00_54_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210055(.x(x_55), .z(tmp00_55_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210056(.x(x_56), .z(tmp00_56_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210057(.x(x_57), .z(tmp00_57_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210058(.x(x_58), .z(tmp00_58_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210059(.x(x_59), .z(tmp00_59_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210060(.x(x_60), .z(tmp00_60_21));
	booth__010 #(.WIDTH(WIDTH)) mul00210061(.x(x_61), .z(tmp00_61_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210062(.x(x_62), .z(tmp00_62_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210063(.x(x_63), .z(tmp00_63_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210064(.x(x_64), .z(tmp00_64_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210065(.x(x_65), .z(tmp00_65_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210066(.x(x_66), .z(tmp00_66_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210067(.x(x_67), .z(tmp00_67_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210068(.x(x_68), .z(tmp00_68_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210069(.x(x_69), .z(tmp00_69_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210070(.x(x_70), .z(tmp00_70_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210071(.x(x_71), .z(tmp00_71_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210072(.x(x_72), .z(tmp00_72_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210073(.x(x_73), .z(tmp00_73_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210074(.x(x_74), .z(tmp00_74_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210075(.x(x_75), .z(tmp00_75_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210076(.x(x_76), .z(tmp00_76_21));
	booth_0006 #(.WIDTH(WIDTH)) mul00210077(.x(x_77), .z(tmp00_77_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210078(.x(x_78), .z(tmp00_78_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210079(.x(x_79), .z(tmp00_79_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210080(.x(x_80), .z(tmp00_80_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210081(.x(x_81), .z(tmp00_81_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210082(.x(x_82), .z(tmp00_82_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210083(.x(x_83), .z(tmp00_83_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210084(.x(x_84), .z(tmp00_84_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210085(.x(x_85), .z(tmp00_85_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210086(.x(x_86), .z(tmp00_86_21));
	booth_0006 #(.WIDTH(WIDTH)) mul00210087(.x(x_87), .z(tmp00_87_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210088(.x(x_88), .z(tmp00_88_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210089(.x(x_89), .z(tmp00_89_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210090(.x(x_90), .z(tmp00_90_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210091(.x(x_91), .z(tmp00_91_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210092(.x(x_92), .z(tmp00_92_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210093(.x(x_93), .z(tmp00_93_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210094(.x(x_94), .z(tmp00_94_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210095(.x(x_95), .z(tmp00_95_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210096(.x(x_96), .z(tmp00_96_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210097(.x(x_97), .z(tmp00_97_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210098(.x(x_98), .z(tmp00_98_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210099(.x(x_99), .z(tmp00_99_21));
	booth_0006 #(.WIDTH(WIDTH)) mul00210100(.x(x_100), .z(tmp00_100_21));
	booth__010 #(.WIDTH(WIDTH)) mul00210101(.x(x_101), .z(tmp00_101_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210102(.x(x_102), .z(tmp00_102_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210103(.x(x_103), .z(tmp00_103_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210104(.x(x_104), .z(tmp00_104_21));
	booth_0004 #(.WIDTH(WIDTH)) mul00210105(.x(x_105), .z(tmp00_105_21));
	booth_0010 #(.WIDTH(WIDTH)) mul00210106(.x(x_106), .z(tmp00_106_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00210107(.x(x_107), .z(tmp00_107_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210108(.x(x_108), .z(tmp00_108_21));
	booth__002 #(.WIDTH(WIDTH)) mul00210109(.x(x_109), .z(tmp00_109_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210110(.x(x_110), .z(tmp00_110_21));
	booth_0002 #(.WIDTH(WIDTH)) mul00210111(.x(x_111), .z(tmp00_111_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210112(.x(x_112), .z(tmp00_112_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210113(.x(x_113), .z(tmp00_113_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210114(.x(x_114), .z(tmp00_114_21));
	booth_0006 #(.WIDTH(WIDTH)) mul00210115(.x(x_115), .z(tmp00_115_21));
	booth_0012 #(.WIDTH(WIDTH)) mul00210116(.x(x_116), .z(tmp00_116_21));
	booth_0010 #(.WIDTH(WIDTH)) mul00210117(.x(x_117), .z(tmp00_117_21));
	booth__004 #(.WIDTH(WIDTH)) mul00210118(.x(x_118), .z(tmp00_118_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210119(.x(x_119), .z(tmp00_119_21));
	booth_0002 #(.WIDTH(WIDTH)) mul00210120(.x(x_120), .z(tmp00_120_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210121(.x(x_121), .z(tmp00_121_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210122(.x(x_122), .z(tmp00_122_21));
	booth_0002 #(.WIDTH(WIDTH)) mul00210123(.x(x_123), .z(tmp00_123_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210124(.x(x_124), .z(tmp00_124_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210125(.x(x_125), .z(tmp00_125_21));
	booth__008 #(.WIDTH(WIDTH)) mul00210126(.x(x_126), .z(tmp00_126_21));
	booth_0000 #(.WIDTH(WIDTH)) mul00210127(.x(x_127), .z(tmp00_127_21));
	booth_0008 #(.WIDTH(WIDTH)) mul00220000(.x(x_0), .z(tmp00_0_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220001(.x(x_1), .z(tmp00_1_22));
	booth_0012 #(.WIDTH(WIDTH)) mul00220002(.x(x_2), .z(tmp00_2_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220003(.x(x_3), .z(tmp00_3_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220004(.x(x_4), .z(tmp00_4_22));
	booth__002 #(.WIDTH(WIDTH)) mul00220005(.x(x_5), .z(tmp00_5_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220006(.x(x_6), .z(tmp00_6_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220007(.x(x_7), .z(tmp00_7_22));
	booth__012 #(.WIDTH(WIDTH)) mul00220008(.x(x_8), .z(tmp00_8_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220009(.x(x_9), .z(tmp00_9_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220010(.x(x_10), .z(tmp00_10_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220011(.x(x_11), .z(tmp00_11_22));
	booth__012 #(.WIDTH(WIDTH)) mul00220012(.x(x_12), .z(tmp00_12_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220013(.x(x_13), .z(tmp00_13_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220014(.x(x_14), .z(tmp00_14_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220015(.x(x_15), .z(tmp00_15_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220016(.x(x_16), .z(tmp00_16_22));
	booth__010 #(.WIDTH(WIDTH)) mul00220017(.x(x_17), .z(tmp00_17_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220018(.x(x_18), .z(tmp00_18_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220019(.x(x_19), .z(tmp00_19_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220020(.x(x_20), .z(tmp00_20_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220021(.x(x_21), .z(tmp00_21_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220022(.x(x_22), .z(tmp00_22_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220023(.x(x_23), .z(tmp00_23_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220024(.x(x_24), .z(tmp00_24_22));
	booth_0016 #(.WIDTH(WIDTH)) mul00220025(.x(x_25), .z(tmp00_25_22));
	booth_0006 #(.WIDTH(WIDTH)) mul00220026(.x(x_26), .z(tmp00_26_22));
	booth__006 #(.WIDTH(WIDTH)) mul00220027(.x(x_27), .z(tmp00_27_22));
	booth_0010 #(.WIDTH(WIDTH)) mul00220028(.x(x_28), .z(tmp00_28_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220029(.x(x_29), .z(tmp00_29_22));
	booth__002 #(.WIDTH(WIDTH)) mul00220030(.x(x_30), .z(tmp00_30_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220031(.x(x_31), .z(tmp00_31_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220032(.x(x_32), .z(tmp00_32_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220033(.x(x_33), .z(tmp00_33_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220034(.x(x_34), .z(tmp00_34_22));
	booth_0006 #(.WIDTH(WIDTH)) mul00220035(.x(x_35), .z(tmp00_35_22));
	booth_0012 #(.WIDTH(WIDTH)) mul00220036(.x(x_36), .z(tmp00_36_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220037(.x(x_37), .z(tmp00_37_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220038(.x(x_38), .z(tmp00_38_22));
	booth__020 #(.WIDTH(WIDTH)) mul00220039(.x(x_39), .z(tmp00_39_22));
	booth_0012 #(.WIDTH(WIDTH)) mul00220040(.x(x_40), .z(tmp00_40_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220041(.x(x_41), .z(tmp00_41_22));
	booth_0016 #(.WIDTH(WIDTH)) mul00220042(.x(x_42), .z(tmp00_42_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220043(.x(x_43), .z(tmp00_43_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220044(.x(x_44), .z(tmp00_44_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220045(.x(x_45), .z(tmp00_45_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220046(.x(x_46), .z(tmp00_46_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220047(.x(x_47), .z(tmp00_47_22));
	booth__002 #(.WIDTH(WIDTH)) mul00220048(.x(x_48), .z(tmp00_48_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220049(.x(x_49), .z(tmp00_49_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220050(.x(x_50), .z(tmp00_50_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220051(.x(x_51), .z(tmp00_51_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220052(.x(x_52), .z(tmp00_52_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220053(.x(x_53), .z(tmp00_53_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220054(.x(x_54), .z(tmp00_54_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220055(.x(x_55), .z(tmp00_55_22));
	booth_0010 #(.WIDTH(WIDTH)) mul00220056(.x(x_56), .z(tmp00_56_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220057(.x(x_57), .z(tmp00_57_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220058(.x(x_58), .z(tmp00_58_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220059(.x(x_59), .z(tmp00_59_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220060(.x(x_60), .z(tmp00_60_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220061(.x(x_61), .z(tmp00_61_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220062(.x(x_62), .z(tmp00_62_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220063(.x(x_63), .z(tmp00_63_22));
	booth_0006 #(.WIDTH(WIDTH)) mul00220064(.x(x_64), .z(tmp00_64_22));
	booth__006 #(.WIDTH(WIDTH)) mul00220065(.x(x_65), .z(tmp00_65_22));
	booth_0012 #(.WIDTH(WIDTH)) mul00220066(.x(x_66), .z(tmp00_66_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220067(.x(x_67), .z(tmp00_67_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220068(.x(x_68), .z(tmp00_68_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220069(.x(x_69), .z(tmp00_69_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220070(.x(x_70), .z(tmp00_70_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220071(.x(x_71), .z(tmp00_71_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220072(.x(x_72), .z(tmp00_72_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220073(.x(x_73), .z(tmp00_73_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220074(.x(x_74), .z(tmp00_74_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220075(.x(x_75), .z(tmp00_75_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220076(.x(x_76), .z(tmp00_76_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220077(.x(x_77), .z(tmp00_77_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220078(.x(x_78), .z(tmp00_78_22));
	booth__006 #(.WIDTH(WIDTH)) mul00220079(.x(x_79), .z(tmp00_79_22));
	booth__002 #(.WIDTH(WIDTH)) mul00220080(.x(x_80), .z(tmp00_80_22));
	booth_0016 #(.WIDTH(WIDTH)) mul00220081(.x(x_81), .z(tmp00_81_22));
	booth__010 #(.WIDTH(WIDTH)) mul00220082(.x(x_82), .z(tmp00_82_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220083(.x(x_83), .z(tmp00_83_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220084(.x(x_84), .z(tmp00_84_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220085(.x(x_85), .z(tmp00_85_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220086(.x(x_86), .z(tmp00_86_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220087(.x(x_87), .z(tmp00_87_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220088(.x(x_88), .z(tmp00_88_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220089(.x(x_89), .z(tmp00_89_22));
	booth_0016 #(.WIDTH(WIDTH)) mul00220090(.x(x_90), .z(tmp00_90_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220091(.x(x_91), .z(tmp00_91_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220092(.x(x_92), .z(tmp00_92_22));
	booth__010 #(.WIDTH(WIDTH)) mul00220093(.x(x_93), .z(tmp00_93_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220094(.x(x_94), .z(tmp00_94_22));
	booth_0006 #(.WIDTH(WIDTH)) mul00220095(.x(x_95), .z(tmp00_95_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220096(.x(x_96), .z(tmp00_96_22));
	booth_0008 #(.WIDTH(WIDTH)) mul00220097(.x(x_97), .z(tmp00_97_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220098(.x(x_98), .z(tmp00_98_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220099(.x(x_99), .z(tmp00_99_22));
	booth_0002 #(.WIDTH(WIDTH)) mul00220100(.x(x_100), .z(tmp00_100_22));
	booth__004 #(.WIDTH(WIDTH)) mul00220101(.x(x_101), .z(tmp00_101_22));
	booth__014 #(.WIDTH(WIDTH)) mul00220102(.x(x_102), .z(tmp00_102_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220103(.x(x_103), .z(tmp00_103_22));
	booth__010 #(.WIDTH(WIDTH)) mul00220104(.x(x_104), .z(tmp00_104_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220105(.x(x_105), .z(tmp00_105_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220106(.x(x_106), .z(tmp00_106_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220107(.x(x_107), .z(tmp00_107_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220108(.x(x_108), .z(tmp00_108_22));
	booth__012 #(.WIDTH(WIDTH)) mul00220109(.x(x_109), .z(tmp00_109_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220110(.x(x_110), .z(tmp00_110_22));
	booth_0012 #(.WIDTH(WIDTH)) mul00220111(.x(x_111), .z(tmp00_111_22));
	booth__002 #(.WIDTH(WIDTH)) mul00220112(.x(x_112), .z(tmp00_112_22));
	booth_0014 #(.WIDTH(WIDTH)) mul00220113(.x(x_113), .z(tmp00_113_22));
	booth_0010 #(.WIDTH(WIDTH)) mul00220114(.x(x_114), .z(tmp00_114_22));
	booth_0014 #(.WIDTH(WIDTH)) mul00220115(.x(x_115), .z(tmp00_115_22));
	booth__010 #(.WIDTH(WIDTH)) mul00220116(.x(x_116), .z(tmp00_116_22));
	booth__002 #(.WIDTH(WIDTH)) mul00220117(.x(x_117), .z(tmp00_117_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220118(.x(x_118), .z(tmp00_118_22));
	booth_0016 #(.WIDTH(WIDTH)) mul00220119(.x(x_119), .z(tmp00_119_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220120(.x(x_120), .z(tmp00_120_22));
	booth__008 #(.WIDTH(WIDTH)) mul00220121(.x(x_121), .z(tmp00_121_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220122(.x(x_122), .z(tmp00_122_22));
	booth__010 #(.WIDTH(WIDTH)) mul00220123(.x(x_123), .z(tmp00_123_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220124(.x(x_124), .z(tmp00_124_22));
	booth_0004 #(.WIDTH(WIDTH)) mul00220125(.x(x_125), .z(tmp00_125_22));
	booth__002 #(.WIDTH(WIDTH)) mul00220126(.x(x_126), .z(tmp00_126_22));
	booth_0000 #(.WIDTH(WIDTH)) mul00220127(.x(x_127), .z(tmp00_127_22));
	booth__006 #(.WIDTH(WIDTH)) mul00230000(.x(x_0), .z(tmp00_0_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230001(.x(x_1), .z(tmp00_1_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230002(.x(x_2), .z(tmp00_2_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230003(.x(x_3), .z(tmp00_3_23));
	booth_0006 #(.WIDTH(WIDTH)) mul00230004(.x(x_4), .z(tmp00_4_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230005(.x(x_5), .z(tmp00_5_23));
	booth__006 #(.WIDTH(WIDTH)) mul00230006(.x(x_6), .z(tmp00_6_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230007(.x(x_7), .z(tmp00_7_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230008(.x(x_8), .z(tmp00_8_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230009(.x(x_9), .z(tmp00_9_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230010(.x(x_10), .z(tmp00_10_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230011(.x(x_11), .z(tmp00_11_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230012(.x(x_12), .z(tmp00_12_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230013(.x(x_13), .z(tmp00_13_23));
	booth_0006 #(.WIDTH(WIDTH)) mul00230014(.x(x_14), .z(tmp00_14_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230015(.x(x_15), .z(tmp00_15_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230016(.x(x_16), .z(tmp00_16_23));
	booth_0010 #(.WIDTH(WIDTH)) mul00230017(.x(x_17), .z(tmp00_17_23));
	booth__006 #(.WIDTH(WIDTH)) mul00230018(.x(x_18), .z(tmp00_18_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230019(.x(x_19), .z(tmp00_19_23));
	booth__010 #(.WIDTH(WIDTH)) mul00230020(.x(x_20), .z(tmp00_20_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230021(.x(x_21), .z(tmp00_21_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230022(.x(x_22), .z(tmp00_22_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230023(.x(x_23), .z(tmp00_23_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230024(.x(x_24), .z(tmp00_24_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230025(.x(x_25), .z(tmp00_25_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230026(.x(x_26), .z(tmp00_26_23));
	booth__006 #(.WIDTH(WIDTH)) mul00230027(.x(x_27), .z(tmp00_27_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230028(.x(x_28), .z(tmp00_28_23));
	booth__002 #(.WIDTH(WIDTH)) mul00230029(.x(x_29), .z(tmp00_29_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230030(.x(x_30), .z(tmp00_30_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230031(.x(x_31), .z(tmp00_31_23));
	booth_0006 #(.WIDTH(WIDTH)) mul00230032(.x(x_32), .z(tmp00_32_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230033(.x(x_33), .z(tmp00_33_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230034(.x(x_34), .z(tmp00_34_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230035(.x(x_35), .z(tmp00_35_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230036(.x(x_36), .z(tmp00_36_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230037(.x(x_37), .z(tmp00_37_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230038(.x(x_38), .z(tmp00_38_23));
	booth__002 #(.WIDTH(WIDTH)) mul00230039(.x(x_39), .z(tmp00_39_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230040(.x(x_40), .z(tmp00_40_23));
	booth__002 #(.WIDTH(WIDTH)) mul00230041(.x(x_41), .z(tmp00_41_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230042(.x(x_42), .z(tmp00_42_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230043(.x(x_43), .z(tmp00_43_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230044(.x(x_44), .z(tmp00_44_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230045(.x(x_45), .z(tmp00_45_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230046(.x(x_46), .z(tmp00_46_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230047(.x(x_47), .z(tmp00_47_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230048(.x(x_48), .z(tmp00_48_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230049(.x(x_49), .z(tmp00_49_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230050(.x(x_50), .z(tmp00_50_23));
	booth_0006 #(.WIDTH(WIDTH)) mul00230051(.x(x_51), .z(tmp00_51_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230052(.x(x_52), .z(tmp00_52_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230053(.x(x_53), .z(tmp00_53_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230054(.x(x_54), .z(tmp00_54_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230055(.x(x_55), .z(tmp00_55_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230056(.x(x_56), .z(tmp00_56_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230057(.x(x_57), .z(tmp00_57_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230058(.x(x_58), .z(tmp00_58_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230059(.x(x_59), .z(tmp00_59_23));
	booth__010 #(.WIDTH(WIDTH)) mul00230060(.x(x_60), .z(tmp00_60_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230061(.x(x_61), .z(tmp00_61_23));
	booth__006 #(.WIDTH(WIDTH)) mul00230062(.x(x_62), .z(tmp00_62_23));
	booth__006 #(.WIDTH(WIDTH)) mul00230063(.x(x_63), .z(tmp00_63_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230064(.x(x_64), .z(tmp00_64_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230065(.x(x_65), .z(tmp00_65_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230066(.x(x_66), .z(tmp00_66_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230067(.x(x_67), .z(tmp00_67_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230068(.x(x_68), .z(tmp00_68_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230069(.x(x_69), .z(tmp00_69_23));
	booth__006 #(.WIDTH(WIDTH)) mul00230070(.x(x_70), .z(tmp00_70_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230071(.x(x_71), .z(tmp00_71_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230072(.x(x_72), .z(tmp00_72_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230073(.x(x_73), .z(tmp00_73_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230074(.x(x_74), .z(tmp00_74_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230075(.x(x_75), .z(tmp00_75_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230076(.x(x_76), .z(tmp00_76_23));
	booth__006 #(.WIDTH(WIDTH)) mul00230077(.x(x_77), .z(tmp00_77_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230078(.x(x_78), .z(tmp00_78_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230079(.x(x_79), .z(tmp00_79_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230080(.x(x_80), .z(tmp00_80_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230081(.x(x_81), .z(tmp00_81_23));
	booth_0010 #(.WIDTH(WIDTH)) mul00230082(.x(x_82), .z(tmp00_82_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230083(.x(x_83), .z(tmp00_83_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230084(.x(x_84), .z(tmp00_84_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230085(.x(x_85), .z(tmp00_85_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230086(.x(x_86), .z(tmp00_86_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230087(.x(x_87), .z(tmp00_87_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230088(.x(x_88), .z(tmp00_88_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230089(.x(x_89), .z(tmp00_89_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230090(.x(x_90), .z(tmp00_90_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230091(.x(x_91), .z(tmp00_91_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230092(.x(x_92), .z(tmp00_92_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230093(.x(x_93), .z(tmp00_93_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230094(.x(x_94), .z(tmp00_94_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230095(.x(x_95), .z(tmp00_95_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230096(.x(x_96), .z(tmp00_96_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230097(.x(x_97), .z(tmp00_97_23));
	booth_0010 #(.WIDTH(WIDTH)) mul00230098(.x(x_98), .z(tmp00_98_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230099(.x(x_99), .z(tmp00_99_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230100(.x(x_100), .z(tmp00_100_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230101(.x(x_101), .z(tmp00_101_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230102(.x(x_102), .z(tmp00_102_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230103(.x(x_103), .z(tmp00_103_23));
	booth__012 #(.WIDTH(WIDTH)) mul00230104(.x(x_104), .z(tmp00_104_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230105(.x(x_105), .z(tmp00_105_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230106(.x(x_106), .z(tmp00_106_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230107(.x(x_107), .z(tmp00_107_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230108(.x(x_108), .z(tmp00_108_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230109(.x(x_109), .z(tmp00_109_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230110(.x(x_110), .z(tmp00_110_23));
	booth_0008 #(.WIDTH(WIDTH)) mul00230111(.x(x_111), .z(tmp00_111_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230112(.x(x_112), .z(tmp00_112_23));
	booth_0010 #(.WIDTH(WIDTH)) mul00230113(.x(x_113), .z(tmp00_113_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230114(.x(x_114), .z(tmp00_114_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230115(.x(x_115), .z(tmp00_115_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230116(.x(x_116), .z(tmp00_116_23));
	booth_0004 #(.WIDTH(WIDTH)) mul00230117(.x(x_117), .z(tmp00_117_23));
	booth_0002 #(.WIDTH(WIDTH)) mul00230118(.x(x_118), .z(tmp00_118_23));
	booth_0006 #(.WIDTH(WIDTH)) mul00230119(.x(x_119), .z(tmp00_119_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230120(.x(x_120), .z(tmp00_120_23));
	booth__012 #(.WIDTH(WIDTH)) mul00230121(.x(x_121), .z(tmp00_121_23));
	booth_0012 #(.WIDTH(WIDTH)) mul00230122(.x(x_122), .z(tmp00_122_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230123(.x(x_123), .z(tmp00_123_23));
	booth__012 #(.WIDTH(WIDTH)) mul00230124(.x(x_124), .z(tmp00_124_23));
	booth__008 #(.WIDTH(WIDTH)) mul00230125(.x(x_125), .z(tmp00_125_23));
	booth_0000 #(.WIDTH(WIDTH)) mul00230126(.x(x_126), .z(tmp00_126_23));
	booth__004 #(.WIDTH(WIDTH)) mul00230127(.x(x_127), .z(tmp00_127_23));
	booth_0010 #(.WIDTH(WIDTH)) mul00240000(.x(x_0), .z(tmp00_0_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240001(.x(x_1), .z(tmp00_1_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240002(.x(x_2), .z(tmp00_2_24));
	booth_0004 #(.WIDTH(WIDTH)) mul00240003(.x(x_3), .z(tmp00_3_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240004(.x(x_4), .z(tmp00_4_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240005(.x(x_5), .z(tmp00_5_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240006(.x(x_6), .z(tmp00_6_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240007(.x(x_7), .z(tmp00_7_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240008(.x(x_8), .z(tmp00_8_24));
	booth__010 #(.WIDTH(WIDTH)) mul00240009(.x(x_9), .z(tmp00_9_24));
	booth_0002 #(.WIDTH(WIDTH)) mul00240010(.x(x_10), .z(tmp00_10_24));
	booth__002 #(.WIDTH(WIDTH)) mul00240011(.x(x_11), .z(tmp00_11_24));
	booth_0004 #(.WIDTH(WIDTH)) mul00240012(.x(x_12), .z(tmp00_12_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240013(.x(x_13), .z(tmp00_13_24));
	booth_0010 #(.WIDTH(WIDTH)) mul00240014(.x(x_14), .z(tmp00_14_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240015(.x(x_15), .z(tmp00_15_24));
	booth_0002 #(.WIDTH(WIDTH)) mul00240016(.x(x_16), .z(tmp00_16_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240017(.x(x_17), .z(tmp00_17_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240018(.x(x_18), .z(tmp00_18_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240019(.x(x_19), .z(tmp00_19_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240020(.x(x_20), .z(tmp00_20_24));
	booth_0006 #(.WIDTH(WIDTH)) mul00240021(.x(x_21), .z(tmp00_21_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240022(.x(x_22), .z(tmp00_22_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240023(.x(x_23), .z(tmp00_23_24));
	booth__012 #(.WIDTH(WIDTH)) mul00240024(.x(x_24), .z(tmp00_24_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240025(.x(x_25), .z(tmp00_25_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240026(.x(x_26), .z(tmp00_26_24));
	booth__002 #(.WIDTH(WIDTH)) mul00240027(.x(x_27), .z(tmp00_27_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240028(.x(x_28), .z(tmp00_28_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240029(.x(x_29), .z(tmp00_29_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240030(.x(x_30), .z(tmp00_30_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240031(.x(x_31), .z(tmp00_31_24));
	booth_0010 #(.WIDTH(WIDTH)) mul00240032(.x(x_32), .z(tmp00_32_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240033(.x(x_33), .z(tmp00_33_24));
	booth__002 #(.WIDTH(WIDTH)) mul00240034(.x(x_34), .z(tmp00_34_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240035(.x(x_35), .z(tmp00_35_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240036(.x(x_36), .z(tmp00_36_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240037(.x(x_37), .z(tmp00_37_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240038(.x(x_38), .z(tmp00_38_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240039(.x(x_39), .z(tmp00_39_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240040(.x(x_40), .z(tmp00_40_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240041(.x(x_41), .z(tmp00_41_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240042(.x(x_42), .z(tmp00_42_24));
	booth__010 #(.WIDTH(WIDTH)) mul00240043(.x(x_43), .z(tmp00_43_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240044(.x(x_44), .z(tmp00_44_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240045(.x(x_45), .z(tmp00_45_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240046(.x(x_46), .z(tmp00_46_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240047(.x(x_47), .z(tmp00_47_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240048(.x(x_48), .z(tmp00_48_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240049(.x(x_49), .z(tmp00_49_24));
	booth_0010 #(.WIDTH(WIDTH)) mul00240050(.x(x_50), .z(tmp00_50_24));
	booth__006 #(.WIDTH(WIDTH)) mul00240051(.x(x_51), .z(tmp00_51_24));
	booth__006 #(.WIDTH(WIDTH)) mul00240052(.x(x_52), .z(tmp00_52_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240053(.x(x_53), .z(tmp00_53_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240054(.x(x_54), .z(tmp00_54_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240055(.x(x_55), .z(tmp00_55_24));
	booth__016 #(.WIDTH(WIDTH)) mul00240056(.x(x_56), .z(tmp00_56_24));
	booth__006 #(.WIDTH(WIDTH)) mul00240057(.x(x_57), .z(tmp00_57_24));
	booth_0012 #(.WIDTH(WIDTH)) mul00240058(.x(x_58), .z(tmp00_58_24));
	booth_0002 #(.WIDTH(WIDTH)) mul00240059(.x(x_59), .z(tmp00_59_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240060(.x(x_60), .z(tmp00_60_24));
	booth_0004 #(.WIDTH(WIDTH)) mul00240061(.x(x_61), .z(tmp00_61_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240062(.x(x_62), .z(tmp00_62_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240063(.x(x_63), .z(tmp00_63_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240064(.x(x_64), .z(tmp00_64_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240065(.x(x_65), .z(tmp00_65_24));
	booth__010 #(.WIDTH(WIDTH)) mul00240066(.x(x_66), .z(tmp00_66_24));
	booth_0012 #(.WIDTH(WIDTH)) mul00240067(.x(x_67), .z(tmp00_67_24));
	booth__016 #(.WIDTH(WIDTH)) mul00240068(.x(x_68), .z(tmp00_68_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240069(.x(x_69), .z(tmp00_69_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240070(.x(x_70), .z(tmp00_70_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240071(.x(x_71), .z(tmp00_71_24));
	booth__010 #(.WIDTH(WIDTH)) mul00240072(.x(x_72), .z(tmp00_72_24));
	booth_0006 #(.WIDTH(WIDTH)) mul00240073(.x(x_73), .z(tmp00_73_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240074(.x(x_74), .z(tmp00_74_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240075(.x(x_75), .z(tmp00_75_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240076(.x(x_76), .z(tmp00_76_24));
	booth_0002 #(.WIDTH(WIDTH)) mul00240077(.x(x_77), .z(tmp00_77_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240078(.x(x_78), .z(tmp00_78_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240079(.x(x_79), .z(tmp00_79_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240080(.x(x_80), .z(tmp00_80_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240081(.x(x_81), .z(tmp00_81_24));
	booth_0012 #(.WIDTH(WIDTH)) mul00240082(.x(x_82), .z(tmp00_82_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240083(.x(x_83), .z(tmp00_83_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240084(.x(x_84), .z(tmp00_84_24));
	booth__014 #(.WIDTH(WIDTH)) mul00240085(.x(x_85), .z(tmp00_85_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240086(.x(x_86), .z(tmp00_86_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240087(.x(x_87), .z(tmp00_87_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240088(.x(x_88), .z(tmp00_88_24));
	booth__008 #(.WIDTH(WIDTH)) mul00240089(.x(x_89), .z(tmp00_89_24));
	booth__012 #(.WIDTH(WIDTH)) mul00240090(.x(x_90), .z(tmp00_90_24));
	booth_0004 #(.WIDTH(WIDTH)) mul00240091(.x(x_91), .z(tmp00_91_24));
	booth_0014 #(.WIDTH(WIDTH)) mul00240092(.x(x_92), .z(tmp00_92_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240093(.x(x_93), .z(tmp00_93_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240094(.x(x_94), .z(tmp00_94_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240095(.x(x_95), .z(tmp00_95_24));
	booth_0002 #(.WIDTH(WIDTH)) mul00240096(.x(x_96), .z(tmp00_96_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240097(.x(x_97), .z(tmp00_97_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240098(.x(x_98), .z(tmp00_98_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240099(.x(x_99), .z(tmp00_99_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240100(.x(x_100), .z(tmp00_100_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240101(.x(x_101), .z(tmp00_101_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240102(.x(x_102), .z(tmp00_102_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240103(.x(x_103), .z(tmp00_103_24));
	booth_0004 #(.WIDTH(WIDTH)) mul00240104(.x(x_104), .z(tmp00_104_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240105(.x(x_105), .z(tmp00_105_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240106(.x(x_106), .z(tmp00_106_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240107(.x(x_107), .z(tmp00_107_24));
	booth__006 #(.WIDTH(WIDTH)) mul00240108(.x(x_108), .z(tmp00_108_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240109(.x(x_109), .z(tmp00_109_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240110(.x(x_110), .z(tmp00_110_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240111(.x(x_111), .z(tmp00_111_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240112(.x(x_112), .z(tmp00_112_24));
	booth_0012 #(.WIDTH(WIDTH)) mul00240113(.x(x_113), .z(tmp00_113_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240114(.x(x_114), .z(tmp00_114_24));
	booth__004 #(.WIDTH(WIDTH)) mul00240115(.x(x_115), .z(tmp00_115_24));
	booth__006 #(.WIDTH(WIDTH)) mul00240116(.x(x_116), .z(tmp00_116_24));
	booth__012 #(.WIDTH(WIDTH)) mul00240117(.x(x_117), .z(tmp00_117_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240118(.x(x_118), .z(tmp00_118_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00240119(.x(x_119), .z(tmp00_119_24));
	booth__016 #(.WIDTH(WIDTH)) mul00240120(.x(x_120), .z(tmp00_120_24));
	booth_0016 #(.WIDTH(WIDTH)) mul00240121(.x(x_121), .z(tmp00_121_24));
	booth_0004 #(.WIDTH(WIDTH)) mul00240122(.x(x_122), .z(tmp00_122_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240123(.x(x_123), .z(tmp00_123_24));
	booth_0008 #(.WIDTH(WIDTH)) mul00240124(.x(x_124), .z(tmp00_124_24));
	booth__010 #(.WIDTH(WIDTH)) mul00240125(.x(x_125), .z(tmp00_125_24));
	booth_0002 #(.WIDTH(WIDTH)) mul00240126(.x(x_126), .z(tmp00_126_24));
	booth_0014 #(.WIDTH(WIDTH)) mul00240127(.x(x_127), .z(tmp00_127_24));
	booth_0000 #(.WIDTH(WIDTH)) mul00250000(.x(x_0), .z(tmp00_0_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250001(.x(x_1), .z(tmp00_1_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250002(.x(x_2), .z(tmp00_2_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250003(.x(x_3), .z(tmp00_3_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250004(.x(x_4), .z(tmp00_4_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250005(.x(x_5), .z(tmp00_5_25));
	booth__010 #(.WIDTH(WIDTH)) mul00250006(.x(x_6), .z(tmp00_6_25));
	booth__006 #(.WIDTH(WIDTH)) mul00250007(.x(x_7), .z(tmp00_7_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250008(.x(x_8), .z(tmp00_8_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250009(.x(x_9), .z(tmp00_9_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250010(.x(x_10), .z(tmp00_10_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250011(.x(x_11), .z(tmp00_11_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250012(.x(x_12), .z(tmp00_12_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250013(.x(x_13), .z(tmp00_13_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250014(.x(x_14), .z(tmp00_14_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250015(.x(x_15), .z(tmp00_15_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250016(.x(x_16), .z(tmp00_16_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250017(.x(x_17), .z(tmp00_17_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250018(.x(x_18), .z(tmp00_18_25));
	booth_0006 #(.WIDTH(WIDTH)) mul00250019(.x(x_19), .z(tmp00_19_25));
	booth__002 #(.WIDTH(WIDTH)) mul00250020(.x(x_20), .z(tmp00_20_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250021(.x(x_21), .z(tmp00_21_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250022(.x(x_22), .z(tmp00_22_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250023(.x(x_23), .z(tmp00_23_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250024(.x(x_24), .z(tmp00_24_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250025(.x(x_25), .z(tmp00_25_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250026(.x(x_26), .z(tmp00_26_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250027(.x(x_27), .z(tmp00_27_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250028(.x(x_28), .z(tmp00_28_25));
	booth__006 #(.WIDTH(WIDTH)) mul00250029(.x(x_29), .z(tmp00_29_25));
	booth_0006 #(.WIDTH(WIDTH)) mul00250030(.x(x_30), .z(tmp00_30_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250031(.x(x_31), .z(tmp00_31_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250032(.x(x_32), .z(tmp00_32_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250033(.x(x_33), .z(tmp00_33_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250034(.x(x_34), .z(tmp00_34_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250035(.x(x_35), .z(tmp00_35_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250036(.x(x_36), .z(tmp00_36_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250037(.x(x_37), .z(tmp00_37_25));
	booth__006 #(.WIDTH(WIDTH)) mul00250038(.x(x_38), .z(tmp00_38_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250039(.x(x_39), .z(tmp00_39_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250040(.x(x_40), .z(tmp00_40_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250041(.x(x_41), .z(tmp00_41_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250042(.x(x_42), .z(tmp00_42_25));
	booth_0010 #(.WIDTH(WIDTH)) mul00250043(.x(x_43), .z(tmp00_43_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250044(.x(x_44), .z(tmp00_44_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250045(.x(x_45), .z(tmp00_45_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250046(.x(x_46), .z(tmp00_46_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250047(.x(x_47), .z(tmp00_47_25));
	booth__010 #(.WIDTH(WIDTH)) mul00250048(.x(x_48), .z(tmp00_48_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250049(.x(x_49), .z(tmp00_49_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250050(.x(x_50), .z(tmp00_50_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250051(.x(x_51), .z(tmp00_51_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250052(.x(x_52), .z(tmp00_52_25));
	booth__006 #(.WIDTH(WIDTH)) mul00250053(.x(x_53), .z(tmp00_53_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250054(.x(x_54), .z(tmp00_54_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250055(.x(x_55), .z(tmp00_55_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250056(.x(x_56), .z(tmp00_56_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250057(.x(x_57), .z(tmp00_57_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250058(.x(x_58), .z(tmp00_58_25));
	booth__006 #(.WIDTH(WIDTH)) mul00250059(.x(x_59), .z(tmp00_59_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250060(.x(x_60), .z(tmp00_60_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250061(.x(x_61), .z(tmp00_61_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250062(.x(x_62), .z(tmp00_62_25));
	booth__010 #(.WIDTH(WIDTH)) mul00250063(.x(x_63), .z(tmp00_63_25));
	booth__010 #(.WIDTH(WIDTH)) mul00250064(.x(x_64), .z(tmp00_64_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250065(.x(x_65), .z(tmp00_65_25));
	booth__006 #(.WIDTH(WIDTH)) mul00250066(.x(x_66), .z(tmp00_66_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250067(.x(x_67), .z(tmp00_67_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250068(.x(x_68), .z(tmp00_68_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250069(.x(x_69), .z(tmp00_69_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250070(.x(x_70), .z(tmp00_70_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250071(.x(x_71), .z(tmp00_71_25));
	booth__010 #(.WIDTH(WIDTH)) mul00250072(.x(x_72), .z(tmp00_72_25));
	booth_0006 #(.WIDTH(WIDTH)) mul00250073(.x(x_73), .z(tmp00_73_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250074(.x(x_74), .z(tmp00_74_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250075(.x(x_75), .z(tmp00_75_25));
	booth_0010 #(.WIDTH(WIDTH)) mul00250076(.x(x_76), .z(tmp00_76_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250077(.x(x_77), .z(tmp00_77_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250078(.x(x_78), .z(tmp00_78_25));
	booth_0012 #(.WIDTH(WIDTH)) mul00250079(.x(x_79), .z(tmp00_79_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250080(.x(x_80), .z(tmp00_80_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250081(.x(x_81), .z(tmp00_81_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250082(.x(x_82), .z(tmp00_82_25));
	booth_0012 #(.WIDTH(WIDTH)) mul00250083(.x(x_83), .z(tmp00_83_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250084(.x(x_84), .z(tmp00_84_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250085(.x(x_85), .z(tmp00_85_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250086(.x(x_86), .z(tmp00_86_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250087(.x(x_87), .z(tmp00_87_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250088(.x(x_88), .z(tmp00_88_25));
	booth__002 #(.WIDTH(WIDTH)) mul00250089(.x(x_89), .z(tmp00_89_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250090(.x(x_90), .z(tmp00_90_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250091(.x(x_91), .z(tmp00_91_25));
	booth_0006 #(.WIDTH(WIDTH)) mul00250092(.x(x_92), .z(tmp00_92_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250093(.x(x_93), .z(tmp00_93_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250094(.x(x_94), .z(tmp00_94_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250095(.x(x_95), .z(tmp00_95_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250096(.x(x_96), .z(tmp00_96_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250097(.x(x_97), .z(tmp00_97_25));
	booth_0002 #(.WIDTH(WIDTH)) mul00250098(.x(x_98), .z(tmp00_98_25));
	booth__002 #(.WIDTH(WIDTH)) mul00250099(.x(x_99), .z(tmp00_99_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250100(.x(x_100), .z(tmp00_100_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250101(.x(x_101), .z(tmp00_101_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250102(.x(x_102), .z(tmp00_102_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250103(.x(x_103), .z(tmp00_103_25));
	booth__010 #(.WIDTH(WIDTH)) mul00250104(.x(x_104), .z(tmp00_104_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250105(.x(x_105), .z(tmp00_105_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250106(.x(x_106), .z(tmp00_106_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250107(.x(x_107), .z(tmp00_107_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250108(.x(x_108), .z(tmp00_108_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250109(.x(x_109), .z(tmp00_109_25));
	booth__008 #(.WIDTH(WIDTH)) mul00250110(.x(x_110), .z(tmp00_110_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250111(.x(x_111), .z(tmp00_111_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250112(.x(x_112), .z(tmp00_112_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250113(.x(x_113), .z(tmp00_113_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250114(.x(x_114), .z(tmp00_114_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250115(.x(x_115), .z(tmp00_115_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250116(.x(x_116), .z(tmp00_116_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250117(.x(x_117), .z(tmp00_117_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250118(.x(x_118), .z(tmp00_118_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250119(.x(x_119), .z(tmp00_119_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00250120(.x(x_120), .z(tmp00_120_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250121(.x(x_121), .z(tmp00_121_25));
	booth__002 #(.WIDTH(WIDTH)) mul00250122(.x(x_122), .z(tmp00_122_25));
	booth_0008 #(.WIDTH(WIDTH)) mul00250123(.x(x_123), .z(tmp00_123_25));
	booth_0004 #(.WIDTH(WIDTH)) mul00250124(.x(x_124), .z(tmp00_124_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250125(.x(x_125), .z(tmp00_125_25));
	booth__004 #(.WIDTH(WIDTH)) mul00250126(.x(x_126), .z(tmp00_126_25));
	booth__002 #(.WIDTH(WIDTH)) mul00250127(.x(x_127), .z(tmp00_127_25));
	booth_0000 #(.WIDTH(WIDTH)) mul00260000(.x(x_0), .z(tmp00_0_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260001(.x(x_1), .z(tmp00_1_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260002(.x(x_2), .z(tmp00_2_26));
	booth__010 #(.WIDTH(WIDTH)) mul00260003(.x(x_3), .z(tmp00_3_26));
	booth__008 #(.WIDTH(WIDTH)) mul00260004(.x(x_4), .z(tmp00_4_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260005(.x(x_5), .z(tmp00_5_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260006(.x(x_6), .z(tmp00_6_26));
	booth_0012 #(.WIDTH(WIDTH)) mul00260007(.x(x_7), .z(tmp00_7_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260008(.x(x_8), .z(tmp00_8_26));
	booth__008 #(.WIDTH(WIDTH)) mul00260009(.x(x_9), .z(tmp00_9_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260010(.x(x_10), .z(tmp00_10_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260011(.x(x_11), .z(tmp00_11_26));
	booth__010 #(.WIDTH(WIDTH)) mul00260012(.x(x_12), .z(tmp00_12_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260013(.x(x_13), .z(tmp00_13_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260014(.x(x_14), .z(tmp00_14_26));
	booth_0010 #(.WIDTH(WIDTH)) mul00260015(.x(x_15), .z(tmp00_15_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260016(.x(x_16), .z(tmp00_16_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260017(.x(x_17), .z(tmp00_17_26));
	booth__010 #(.WIDTH(WIDTH)) mul00260018(.x(x_18), .z(tmp00_18_26));
	booth_0006 #(.WIDTH(WIDTH)) mul00260019(.x(x_19), .z(tmp00_19_26));
	booth__008 #(.WIDTH(WIDTH)) mul00260020(.x(x_20), .z(tmp00_20_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260021(.x(x_21), .z(tmp00_21_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260022(.x(x_22), .z(tmp00_22_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260023(.x(x_23), .z(tmp00_23_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260024(.x(x_24), .z(tmp00_24_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260025(.x(x_25), .z(tmp00_25_26));
	booth_0006 #(.WIDTH(WIDTH)) mul00260026(.x(x_26), .z(tmp00_26_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260027(.x(x_27), .z(tmp00_27_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260028(.x(x_28), .z(tmp00_28_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260029(.x(x_29), .z(tmp00_29_26));
	booth__006 #(.WIDTH(WIDTH)) mul00260030(.x(x_30), .z(tmp00_30_26));
	booth__006 #(.WIDTH(WIDTH)) mul00260031(.x(x_31), .z(tmp00_31_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260032(.x(x_32), .z(tmp00_32_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260033(.x(x_33), .z(tmp00_33_26));
	booth_0012 #(.WIDTH(WIDTH)) mul00260034(.x(x_34), .z(tmp00_34_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260035(.x(x_35), .z(tmp00_35_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260036(.x(x_36), .z(tmp00_36_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260037(.x(x_37), .z(tmp00_37_26));
	booth__010 #(.WIDTH(WIDTH)) mul00260038(.x(x_38), .z(tmp00_38_26));
	booth_0016 #(.WIDTH(WIDTH)) mul00260039(.x(x_39), .z(tmp00_39_26));
	booth_0016 #(.WIDTH(WIDTH)) mul00260040(.x(x_40), .z(tmp00_40_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260041(.x(x_41), .z(tmp00_41_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260042(.x(x_42), .z(tmp00_42_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260043(.x(x_43), .z(tmp00_43_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260044(.x(x_44), .z(tmp00_44_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260045(.x(x_45), .z(tmp00_45_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260046(.x(x_46), .z(tmp00_46_26));
	booth_0002 #(.WIDTH(WIDTH)) mul00260047(.x(x_47), .z(tmp00_47_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260048(.x(x_48), .z(tmp00_48_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260049(.x(x_49), .z(tmp00_49_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260050(.x(x_50), .z(tmp00_50_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260051(.x(x_51), .z(tmp00_51_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260052(.x(x_52), .z(tmp00_52_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260053(.x(x_53), .z(tmp00_53_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260054(.x(x_54), .z(tmp00_54_26));
	booth__010 #(.WIDTH(WIDTH)) mul00260055(.x(x_55), .z(tmp00_55_26));
	booth_0012 #(.WIDTH(WIDTH)) mul00260056(.x(x_56), .z(tmp00_56_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260057(.x(x_57), .z(tmp00_57_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260058(.x(x_58), .z(tmp00_58_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260059(.x(x_59), .z(tmp00_59_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260060(.x(x_60), .z(tmp00_60_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260061(.x(x_61), .z(tmp00_61_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260062(.x(x_62), .z(tmp00_62_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260063(.x(x_63), .z(tmp00_63_26));
	booth__012 #(.WIDTH(WIDTH)) mul00260064(.x(x_64), .z(tmp00_64_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260065(.x(x_65), .z(tmp00_65_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260066(.x(x_66), .z(tmp00_66_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260067(.x(x_67), .z(tmp00_67_26));
	booth_0002 #(.WIDTH(WIDTH)) mul00260068(.x(x_68), .z(tmp00_68_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260069(.x(x_69), .z(tmp00_69_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260070(.x(x_70), .z(tmp00_70_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260071(.x(x_71), .z(tmp00_71_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260072(.x(x_72), .z(tmp00_72_26));
	booth__008 #(.WIDTH(WIDTH)) mul00260073(.x(x_73), .z(tmp00_73_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260074(.x(x_74), .z(tmp00_74_26));
	booth__012 #(.WIDTH(WIDTH)) mul00260075(.x(x_75), .z(tmp00_75_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260076(.x(x_76), .z(tmp00_76_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260077(.x(x_77), .z(tmp00_77_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260078(.x(x_78), .z(tmp00_78_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260079(.x(x_79), .z(tmp00_79_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260080(.x(x_80), .z(tmp00_80_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260081(.x(x_81), .z(tmp00_81_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260082(.x(x_82), .z(tmp00_82_26));
	booth_0010 #(.WIDTH(WIDTH)) mul00260083(.x(x_83), .z(tmp00_83_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260084(.x(x_84), .z(tmp00_84_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260085(.x(x_85), .z(tmp00_85_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260086(.x(x_86), .z(tmp00_86_26));
	booth_0014 #(.WIDTH(WIDTH)) mul00260087(.x(x_87), .z(tmp00_87_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260088(.x(x_88), .z(tmp00_88_26));
	booth_0006 #(.WIDTH(WIDTH)) mul00260089(.x(x_89), .z(tmp00_89_26));
	booth_0002 #(.WIDTH(WIDTH)) mul00260090(.x(x_90), .z(tmp00_90_26));
	booth_0012 #(.WIDTH(WIDTH)) mul00260091(.x(x_91), .z(tmp00_91_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260092(.x(x_92), .z(tmp00_92_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260093(.x(x_93), .z(tmp00_93_26));
	booth__008 #(.WIDTH(WIDTH)) mul00260094(.x(x_94), .z(tmp00_94_26));
	booth__010 #(.WIDTH(WIDTH)) mul00260095(.x(x_95), .z(tmp00_95_26));
	booth_0002 #(.WIDTH(WIDTH)) mul00260096(.x(x_96), .z(tmp00_96_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260097(.x(x_97), .z(tmp00_97_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260098(.x(x_98), .z(tmp00_98_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260099(.x(x_99), .z(tmp00_99_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260100(.x(x_100), .z(tmp00_100_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260101(.x(x_101), .z(tmp00_101_26));
	booth__006 #(.WIDTH(WIDTH)) mul00260102(.x(x_102), .z(tmp00_102_26));
	booth_0012 #(.WIDTH(WIDTH)) mul00260103(.x(x_103), .z(tmp00_103_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260104(.x(x_104), .z(tmp00_104_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260105(.x(x_105), .z(tmp00_105_26));
	booth_0004 #(.WIDTH(WIDTH)) mul00260106(.x(x_106), .z(tmp00_106_26));
	booth__008 #(.WIDTH(WIDTH)) mul00260107(.x(x_107), .z(tmp00_107_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260108(.x(x_108), .z(tmp00_108_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260109(.x(x_109), .z(tmp00_109_26));
	booth__008 #(.WIDTH(WIDTH)) mul00260110(.x(x_110), .z(tmp00_110_26));
	booth__008 #(.WIDTH(WIDTH)) mul00260111(.x(x_111), .z(tmp00_111_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260112(.x(x_112), .z(tmp00_112_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260113(.x(x_113), .z(tmp00_113_26));
	booth_0008 #(.WIDTH(WIDTH)) mul00260114(.x(x_114), .z(tmp00_114_26));
	booth__002 #(.WIDTH(WIDTH)) mul00260115(.x(x_115), .z(tmp00_115_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260116(.x(x_116), .z(tmp00_116_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260117(.x(x_117), .z(tmp00_117_26));
	booth__012 #(.WIDTH(WIDTH)) mul00260118(.x(x_118), .z(tmp00_118_26));
	booth__016 #(.WIDTH(WIDTH)) mul00260119(.x(x_119), .z(tmp00_119_26));
	booth_0012 #(.WIDTH(WIDTH)) mul00260120(.x(x_120), .z(tmp00_120_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260121(.x(x_121), .z(tmp00_121_26));
	booth_0002 #(.WIDTH(WIDTH)) mul00260122(.x(x_122), .z(tmp00_122_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260123(.x(x_123), .z(tmp00_123_26));
	booth_0016 #(.WIDTH(WIDTH)) mul00260124(.x(x_124), .z(tmp00_124_26));
	booth__004 #(.WIDTH(WIDTH)) mul00260125(.x(x_125), .z(tmp00_125_26));
	booth__012 #(.WIDTH(WIDTH)) mul00260126(.x(x_126), .z(tmp00_126_26));
	booth_0000 #(.WIDTH(WIDTH)) mul00260127(.x(x_127), .z(tmp00_127_26));
	booth__008 #(.WIDTH(WIDTH)) mul00270000(.x(x_0), .z(tmp00_0_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270001(.x(x_1), .z(tmp00_1_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270002(.x(x_2), .z(tmp00_2_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270003(.x(x_3), .z(tmp00_3_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270004(.x(x_4), .z(tmp00_4_27));
	booth_0012 #(.WIDTH(WIDTH)) mul00270005(.x(x_5), .z(tmp00_5_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270006(.x(x_6), .z(tmp00_6_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270007(.x(x_7), .z(tmp00_7_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270008(.x(x_8), .z(tmp00_8_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270009(.x(x_9), .z(tmp00_9_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270010(.x(x_10), .z(tmp00_10_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270011(.x(x_11), .z(tmp00_11_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270012(.x(x_12), .z(tmp00_12_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270013(.x(x_13), .z(tmp00_13_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270014(.x(x_14), .z(tmp00_14_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270015(.x(x_15), .z(tmp00_15_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270016(.x(x_16), .z(tmp00_16_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270017(.x(x_17), .z(tmp00_17_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270018(.x(x_18), .z(tmp00_18_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270019(.x(x_19), .z(tmp00_19_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270020(.x(x_20), .z(tmp00_20_27));
	booth__002 #(.WIDTH(WIDTH)) mul00270021(.x(x_21), .z(tmp00_21_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270022(.x(x_22), .z(tmp00_22_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270023(.x(x_23), .z(tmp00_23_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270024(.x(x_24), .z(tmp00_24_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270025(.x(x_25), .z(tmp00_25_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270026(.x(x_26), .z(tmp00_26_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270027(.x(x_27), .z(tmp00_27_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270028(.x(x_28), .z(tmp00_28_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270029(.x(x_29), .z(tmp00_29_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270030(.x(x_30), .z(tmp00_30_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270031(.x(x_31), .z(tmp00_31_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270032(.x(x_32), .z(tmp00_32_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270033(.x(x_33), .z(tmp00_33_27));
	booth__012 #(.WIDTH(WIDTH)) mul00270034(.x(x_34), .z(tmp00_34_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270035(.x(x_35), .z(tmp00_35_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270036(.x(x_36), .z(tmp00_36_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270037(.x(x_37), .z(tmp00_37_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270038(.x(x_38), .z(tmp00_38_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270039(.x(x_39), .z(tmp00_39_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270040(.x(x_40), .z(tmp00_40_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270041(.x(x_41), .z(tmp00_41_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270042(.x(x_42), .z(tmp00_42_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270043(.x(x_43), .z(tmp00_43_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270044(.x(x_44), .z(tmp00_44_27));
	booth_0012 #(.WIDTH(WIDTH)) mul00270045(.x(x_45), .z(tmp00_45_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270046(.x(x_46), .z(tmp00_46_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270047(.x(x_47), .z(tmp00_47_27));
	booth_0002 #(.WIDTH(WIDTH)) mul00270048(.x(x_48), .z(tmp00_48_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270049(.x(x_49), .z(tmp00_49_27));
	booth__006 #(.WIDTH(WIDTH)) mul00270050(.x(x_50), .z(tmp00_50_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270051(.x(x_51), .z(tmp00_51_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270052(.x(x_52), .z(tmp00_52_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270053(.x(x_53), .z(tmp00_53_27));
	booth_0002 #(.WIDTH(WIDTH)) mul00270054(.x(x_54), .z(tmp00_54_27));
	booth__012 #(.WIDTH(WIDTH)) mul00270055(.x(x_55), .z(tmp00_55_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270056(.x(x_56), .z(tmp00_56_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270057(.x(x_57), .z(tmp00_57_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270058(.x(x_58), .z(tmp00_58_27));
	booth_0006 #(.WIDTH(WIDTH)) mul00270059(.x(x_59), .z(tmp00_59_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270060(.x(x_60), .z(tmp00_60_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270061(.x(x_61), .z(tmp00_61_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270062(.x(x_62), .z(tmp00_62_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270063(.x(x_63), .z(tmp00_63_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270064(.x(x_64), .z(tmp00_64_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270065(.x(x_65), .z(tmp00_65_27));
	booth_0006 #(.WIDTH(WIDTH)) mul00270066(.x(x_66), .z(tmp00_66_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270067(.x(x_67), .z(tmp00_67_27));
	booth__006 #(.WIDTH(WIDTH)) mul00270068(.x(x_68), .z(tmp00_68_27));
	booth__002 #(.WIDTH(WIDTH)) mul00270069(.x(x_69), .z(tmp00_69_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270070(.x(x_70), .z(tmp00_70_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270071(.x(x_71), .z(tmp00_71_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270072(.x(x_72), .z(tmp00_72_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270073(.x(x_73), .z(tmp00_73_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270074(.x(x_74), .z(tmp00_74_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270075(.x(x_75), .z(tmp00_75_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270076(.x(x_76), .z(tmp00_76_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270077(.x(x_77), .z(tmp00_77_27));
	booth__006 #(.WIDTH(WIDTH)) mul00270078(.x(x_78), .z(tmp00_78_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270079(.x(x_79), .z(tmp00_79_27));
	booth__012 #(.WIDTH(WIDTH)) mul00270080(.x(x_80), .z(tmp00_80_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270081(.x(x_81), .z(tmp00_81_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270082(.x(x_82), .z(tmp00_82_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270083(.x(x_83), .z(tmp00_83_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270084(.x(x_84), .z(tmp00_84_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270085(.x(x_85), .z(tmp00_85_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270086(.x(x_86), .z(tmp00_86_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270087(.x(x_87), .z(tmp00_87_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270088(.x(x_88), .z(tmp00_88_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270089(.x(x_89), .z(tmp00_89_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270090(.x(x_90), .z(tmp00_90_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270091(.x(x_91), .z(tmp00_91_27));
	booth_0002 #(.WIDTH(WIDTH)) mul00270092(.x(x_92), .z(tmp00_92_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270093(.x(x_93), .z(tmp00_93_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270094(.x(x_94), .z(tmp00_94_27));
	booth__002 #(.WIDTH(WIDTH)) mul00270095(.x(x_95), .z(tmp00_95_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270096(.x(x_96), .z(tmp00_96_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270097(.x(x_97), .z(tmp00_97_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270098(.x(x_98), .z(tmp00_98_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270099(.x(x_99), .z(tmp00_99_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270100(.x(x_100), .z(tmp00_100_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270101(.x(x_101), .z(tmp00_101_27));
	booth__006 #(.WIDTH(WIDTH)) mul00270102(.x(x_102), .z(tmp00_102_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270103(.x(x_103), .z(tmp00_103_27));
	booth__002 #(.WIDTH(WIDTH)) mul00270104(.x(x_104), .z(tmp00_104_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270105(.x(x_105), .z(tmp00_105_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270106(.x(x_106), .z(tmp00_106_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00270107(.x(x_107), .z(tmp00_107_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270108(.x(x_108), .z(tmp00_108_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270109(.x(x_109), .z(tmp00_109_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270110(.x(x_110), .z(tmp00_110_27));
	booth_0008 #(.WIDTH(WIDTH)) mul00270111(.x(x_111), .z(tmp00_111_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270112(.x(x_112), .z(tmp00_112_27));
	booth__008 #(.WIDTH(WIDTH)) mul00270113(.x(x_113), .z(tmp00_113_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270114(.x(x_114), .z(tmp00_114_27));
	booth__002 #(.WIDTH(WIDTH)) mul00270115(.x(x_115), .z(tmp00_115_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270116(.x(x_116), .z(tmp00_116_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270117(.x(x_117), .z(tmp00_117_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270118(.x(x_118), .z(tmp00_118_27));
	booth_0000 #(.WIDTH(WIDTH)) mul00270119(.x(x_119), .z(tmp00_119_27));
	booth__010 #(.WIDTH(WIDTH)) mul00270120(.x(x_120), .z(tmp00_120_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270121(.x(x_121), .z(tmp00_121_27));
	booth__002 #(.WIDTH(WIDTH)) mul00270122(.x(x_122), .z(tmp00_122_27));
	booth__004 #(.WIDTH(WIDTH)) mul00270123(.x(x_123), .z(tmp00_123_27));
	booth__002 #(.WIDTH(WIDTH)) mul00270124(.x(x_124), .z(tmp00_124_27));
	booth_0004 #(.WIDTH(WIDTH)) mul00270125(.x(x_125), .z(tmp00_125_27));
	booth__006 #(.WIDTH(WIDTH)) mul00270126(.x(x_126), .z(tmp00_126_27));
	booth_0006 #(.WIDTH(WIDTH)) mul00270127(.x(x_127), .z(tmp00_127_27));
	booth_0010 #(.WIDTH(WIDTH)) mul00280000(.x(x_0), .z(tmp00_0_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280001(.x(x_1), .z(tmp00_1_28));
	booth_0002 #(.WIDTH(WIDTH)) mul00280002(.x(x_2), .z(tmp00_2_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280003(.x(x_3), .z(tmp00_3_28));
	booth_0016 #(.WIDTH(WIDTH)) mul00280004(.x(x_4), .z(tmp00_4_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280005(.x(x_5), .z(tmp00_5_28));
	booth_0014 #(.WIDTH(WIDTH)) mul00280006(.x(x_6), .z(tmp00_6_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280007(.x(x_7), .z(tmp00_7_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280008(.x(x_8), .z(tmp00_8_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280009(.x(x_9), .z(tmp00_9_28));
	booth__006 #(.WIDTH(WIDTH)) mul00280010(.x(x_10), .z(tmp00_10_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280011(.x(x_11), .z(tmp00_11_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280012(.x(x_12), .z(tmp00_12_28));
	booth_0012 #(.WIDTH(WIDTH)) mul00280013(.x(x_13), .z(tmp00_13_28));
	booth__006 #(.WIDTH(WIDTH)) mul00280014(.x(x_14), .z(tmp00_14_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280015(.x(x_15), .z(tmp00_15_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280016(.x(x_16), .z(tmp00_16_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280017(.x(x_17), .z(tmp00_17_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280018(.x(x_18), .z(tmp00_18_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280019(.x(x_19), .z(tmp00_19_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280020(.x(x_20), .z(tmp00_20_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280021(.x(x_21), .z(tmp00_21_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280022(.x(x_22), .z(tmp00_22_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280023(.x(x_23), .z(tmp00_23_28));
	booth__010 #(.WIDTH(WIDTH)) mul00280024(.x(x_24), .z(tmp00_24_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280025(.x(x_25), .z(tmp00_25_28));
	booth_0006 #(.WIDTH(WIDTH)) mul00280026(.x(x_26), .z(tmp00_26_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280027(.x(x_27), .z(tmp00_27_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280028(.x(x_28), .z(tmp00_28_28));
	booth__002 #(.WIDTH(WIDTH)) mul00280029(.x(x_29), .z(tmp00_29_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280030(.x(x_30), .z(tmp00_30_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280031(.x(x_31), .z(tmp00_31_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280032(.x(x_32), .z(tmp00_32_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280033(.x(x_33), .z(tmp00_33_28));
	booth__012 #(.WIDTH(WIDTH)) mul00280034(.x(x_34), .z(tmp00_34_28));
	booth_0012 #(.WIDTH(WIDTH)) mul00280035(.x(x_35), .z(tmp00_35_28));
	booth_0006 #(.WIDTH(WIDTH)) mul00280036(.x(x_36), .z(tmp00_36_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280037(.x(x_37), .z(tmp00_37_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280038(.x(x_38), .z(tmp00_38_28));
	booth__002 #(.WIDTH(WIDTH)) mul00280039(.x(x_39), .z(tmp00_39_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280040(.x(x_40), .z(tmp00_40_28));
	booth__006 #(.WIDTH(WIDTH)) mul00280041(.x(x_41), .z(tmp00_41_28));
	booth_0010 #(.WIDTH(WIDTH)) mul00280042(.x(x_42), .z(tmp00_42_28));
	booth_0010 #(.WIDTH(WIDTH)) mul00280043(.x(x_43), .z(tmp00_43_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280044(.x(x_44), .z(tmp00_44_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280045(.x(x_45), .z(tmp00_45_28));
	booth_0012 #(.WIDTH(WIDTH)) mul00280046(.x(x_46), .z(tmp00_46_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280047(.x(x_47), .z(tmp00_47_28));
	booth__012 #(.WIDTH(WIDTH)) mul00280048(.x(x_48), .z(tmp00_48_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280049(.x(x_49), .z(tmp00_49_28));
	booth__010 #(.WIDTH(WIDTH)) mul00280050(.x(x_50), .z(tmp00_50_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280051(.x(x_51), .z(tmp00_51_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280052(.x(x_52), .z(tmp00_52_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280053(.x(x_53), .z(tmp00_53_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280054(.x(x_54), .z(tmp00_54_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280055(.x(x_55), .z(tmp00_55_28));
	booth_0002 #(.WIDTH(WIDTH)) mul00280056(.x(x_56), .z(tmp00_56_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280057(.x(x_57), .z(tmp00_57_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280058(.x(x_58), .z(tmp00_58_28));
	booth__012 #(.WIDTH(WIDTH)) mul00280059(.x(x_59), .z(tmp00_59_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280060(.x(x_60), .z(tmp00_60_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280061(.x(x_61), .z(tmp00_61_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280062(.x(x_62), .z(tmp00_62_28));
	booth_0002 #(.WIDTH(WIDTH)) mul00280063(.x(x_63), .z(tmp00_63_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280064(.x(x_64), .z(tmp00_64_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280065(.x(x_65), .z(tmp00_65_28));
	booth_0012 #(.WIDTH(WIDTH)) mul00280066(.x(x_66), .z(tmp00_66_28));
	booth__002 #(.WIDTH(WIDTH)) mul00280067(.x(x_67), .z(tmp00_67_28));
	booth_0006 #(.WIDTH(WIDTH)) mul00280068(.x(x_68), .z(tmp00_68_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280069(.x(x_69), .z(tmp00_69_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280070(.x(x_70), .z(tmp00_70_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280071(.x(x_71), .z(tmp00_71_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280072(.x(x_72), .z(tmp00_72_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280073(.x(x_73), .z(tmp00_73_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280074(.x(x_74), .z(tmp00_74_28));
	booth__006 #(.WIDTH(WIDTH)) mul00280075(.x(x_75), .z(tmp00_75_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280076(.x(x_76), .z(tmp00_76_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280077(.x(x_77), .z(tmp00_77_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280078(.x(x_78), .z(tmp00_78_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280079(.x(x_79), .z(tmp00_79_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280080(.x(x_80), .z(tmp00_80_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280081(.x(x_81), .z(tmp00_81_28));
	booth__002 #(.WIDTH(WIDTH)) mul00280082(.x(x_82), .z(tmp00_82_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280083(.x(x_83), .z(tmp00_83_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280084(.x(x_84), .z(tmp00_84_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280085(.x(x_85), .z(tmp00_85_28));
	booth__010 #(.WIDTH(WIDTH)) mul00280086(.x(x_86), .z(tmp00_86_28));
	booth_0014 #(.WIDTH(WIDTH)) mul00280087(.x(x_87), .z(tmp00_87_28));
	booth_0012 #(.WIDTH(WIDTH)) mul00280088(.x(x_88), .z(tmp00_88_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280089(.x(x_89), .z(tmp00_89_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280090(.x(x_90), .z(tmp00_90_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280091(.x(x_91), .z(tmp00_91_28));
	booth__006 #(.WIDTH(WIDTH)) mul00280092(.x(x_92), .z(tmp00_92_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280093(.x(x_93), .z(tmp00_93_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280094(.x(x_94), .z(tmp00_94_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280095(.x(x_95), .z(tmp00_95_28));
	booth_0016 #(.WIDTH(WIDTH)) mul00280096(.x(x_96), .z(tmp00_96_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280097(.x(x_97), .z(tmp00_97_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280098(.x(x_98), .z(tmp00_98_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280099(.x(x_99), .z(tmp00_99_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280100(.x(x_100), .z(tmp00_100_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280101(.x(x_101), .z(tmp00_101_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280102(.x(x_102), .z(tmp00_102_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280103(.x(x_103), .z(tmp00_103_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280104(.x(x_104), .z(tmp00_104_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280105(.x(x_105), .z(tmp00_105_28));
	booth__010 #(.WIDTH(WIDTH)) mul00280106(.x(x_106), .z(tmp00_106_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280107(.x(x_107), .z(tmp00_107_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280108(.x(x_108), .z(tmp00_108_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280109(.x(x_109), .z(tmp00_109_28));
	booth_0008 #(.WIDTH(WIDTH)) mul00280110(.x(x_110), .z(tmp00_110_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280111(.x(x_111), .z(tmp00_111_28));
	booth__002 #(.WIDTH(WIDTH)) mul00280112(.x(x_112), .z(tmp00_112_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280113(.x(x_113), .z(tmp00_113_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280114(.x(x_114), .z(tmp00_114_28));
	booth__006 #(.WIDTH(WIDTH)) mul00280115(.x(x_115), .z(tmp00_115_28));
	booth__004 #(.WIDTH(WIDTH)) mul00280116(.x(x_116), .z(tmp00_116_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280117(.x(x_117), .z(tmp00_117_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280118(.x(x_118), .z(tmp00_118_28));
	booth_0012 #(.WIDTH(WIDTH)) mul00280119(.x(x_119), .z(tmp00_119_28));
	booth_0004 #(.WIDTH(WIDTH)) mul00280120(.x(x_120), .z(tmp00_120_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280121(.x(x_121), .z(tmp00_121_28));
	booth__010 #(.WIDTH(WIDTH)) mul00280122(.x(x_122), .z(tmp00_122_28));
	booth__008 #(.WIDTH(WIDTH)) mul00280123(.x(x_123), .z(tmp00_123_28));
	booth_0006 #(.WIDTH(WIDTH)) mul00280124(.x(x_124), .z(tmp00_124_28));
	booth_0006 #(.WIDTH(WIDTH)) mul00280125(.x(x_125), .z(tmp00_125_28));
	booth__012 #(.WIDTH(WIDTH)) mul00280126(.x(x_126), .z(tmp00_126_28));
	booth_0000 #(.WIDTH(WIDTH)) mul00280127(.x(x_127), .z(tmp00_127_28));
	booth__002 #(.WIDTH(WIDTH)) mul00290000(.x(x_0), .z(tmp00_0_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290001(.x(x_1), .z(tmp00_1_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290002(.x(x_2), .z(tmp00_2_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290003(.x(x_3), .z(tmp00_3_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290004(.x(x_4), .z(tmp00_4_29));
	booth__006 #(.WIDTH(WIDTH)) mul00290005(.x(x_5), .z(tmp00_5_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290006(.x(x_6), .z(tmp00_6_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290007(.x(x_7), .z(tmp00_7_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290008(.x(x_8), .z(tmp00_8_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290009(.x(x_9), .z(tmp00_9_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290010(.x(x_10), .z(tmp00_10_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290011(.x(x_11), .z(tmp00_11_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290012(.x(x_12), .z(tmp00_12_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290013(.x(x_13), .z(tmp00_13_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290014(.x(x_14), .z(tmp00_14_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290015(.x(x_15), .z(tmp00_15_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290016(.x(x_16), .z(tmp00_16_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290017(.x(x_17), .z(tmp00_17_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290018(.x(x_18), .z(tmp00_18_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290019(.x(x_19), .z(tmp00_19_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290020(.x(x_20), .z(tmp00_20_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290021(.x(x_21), .z(tmp00_21_29));
	booth__012 #(.WIDTH(WIDTH)) mul00290022(.x(x_22), .z(tmp00_22_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290023(.x(x_23), .z(tmp00_23_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290024(.x(x_24), .z(tmp00_24_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290025(.x(x_25), .z(tmp00_25_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290026(.x(x_26), .z(tmp00_26_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290027(.x(x_27), .z(tmp00_27_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290028(.x(x_28), .z(tmp00_28_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290029(.x(x_29), .z(tmp00_29_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290030(.x(x_30), .z(tmp00_30_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290031(.x(x_31), .z(tmp00_31_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290032(.x(x_32), .z(tmp00_32_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290033(.x(x_33), .z(tmp00_33_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290034(.x(x_34), .z(tmp00_34_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290035(.x(x_35), .z(tmp00_35_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290036(.x(x_36), .z(tmp00_36_29));
	booth__006 #(.WIDTH(WIDTH)) mul00290037(.x(x_37), .z(tmp00_37_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290038(.x(x_38), .z(tmp00_38_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290039(.x(x_39), .z(tmp00_39_29));
	booth_0002 #(.WIDTH(WIDTH)) mul00290040(.x(x_40), .z(tmp00_40_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290041(.x(x_41), .z(tmp00_41_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290042(.x(x_42), .z(tmp00_42_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290043(.x(x_43), .z(tmp00_43_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290044(.x(x_44), .z(tmp00_44_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290045(.x(x_45), .z(tmp00_45_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290046(.x(x_46), .z(tmp00_46_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290047(.x(x_47), .z(tmp00_47_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290048(.x(x_48), .z(tmp00_48_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290049(.x(x_49), .z(tmp00_49_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290050(.x(x_50), .z(tmp00_50_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290051(.x(x_51), .z(tmp00_51_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290052(.x(x_52), .z(tmp00_52_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290053(.x(x_53), .z(tmp00_53_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290054(.x(x_54), .z(tmp00_54_29));
	booth__002 #(.WIDTH(WIDTH)) mul00290055(.x(x_55), .z(tmp00_55_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290056(.x(x_56), .z(tmp00_56_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290057(.x(x_57), .z(tmp00_57_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290058(.x(x_58), .z(tmp00_58_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290059(.x(x_59), .z(tmp00_59_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290060(.x(x_60), .z(tmp00_60_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290061(.x(x_61), .z(tmp00_61_29));
	booth__006 #(.WIDTH(WIDTH)) mul00290062(.x(x_62), .z(tmp00_62_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290063(.x(x_63), .z(tmp00_63_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290064(.x(x_64), .z(tmp00_64_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290065(.x(x_65), .z(tmp00_65_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290066(.x(x_66), .z(tmp00_66_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290067(.x(x_67), .z(tmp00_67_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290068(.x(x_68), .z(tmp00_68_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290069(.x(x_69), .z(tmp00_69_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290070(.x(x_70), .z(tmp00_70_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290071(.x(x_71), .z(tmp00_71_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290072(.x(x_72), .z(tmp00_72_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290073(.x(x_73), .z(tmp00_73_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290074(.x(x_74), .z(tmp00_74_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290075(.x(x_75), .z(tmp00_75_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290076(.x(x_76), .z(tmp00_76_29));
	booth_0006 #(.WIDTH(WIDTH)) mul00290077(.x(x_77), .z(tmp00_77_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290078(.x(x_78), .z(tmp00_78_29));
	booth__006 #(.WIDTH(WIDTH)) mul00290079(.x(x_79), .z(tmp00_79_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290080(.x(x_80), .z(tmp00_80_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290081(.x(x_81), .z(tmp00_81_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290082(.x(x_82), .z(tmp00_82_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290083(.x(x_83), .z(tmp00_83_29));
	booth_0006 #(.WIDTH(WIDTH)) mul00290084(.x(x_84), .z(tmp00_84_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290085(.x(x_85), .z(tmp00_85_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290086(.x(x_86), .z(tmp00_86_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290087(.x(x_87), .z(tmp00_87_29));
	booth_0012 #(.WIDTH(WIDTH)) mul00290088(.x(x_88), .z(tmp00_88_29));
	booth__002 #(.WIDTH(WIDTH)) mul00290089(.x(x_89), .z(tmp00_89_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290090(.x(x_90), .z(tmp00_90_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290091(.x(x_91), .z(tmp00_91_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290092(.x(x_92), .z(tmp00_92_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290093(.x(x_93), .z(tmp00_93_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290094(.x(x_94), .z(tmp00_94_29));
	booth__002 #(.WIDTH(WIDTH)) mul00290095(.x(x_95), .z(tmp00_95_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290096(.x(x_96), .z(tmp00_96_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290097(.x(x_97), .z(tmp00_97_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290098(.x(x_98), .z(tmp00_98_29));
	booth_0002 #(.WIDTH(WIDTH)) mul00290099(.x(x_99), .z(tmp00_99_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290100(.x(x_100), .z(tmp00_100_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290101(.x(x_101), .z(tmp00_101_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290102(.x(x_102), .z(tmp00_102_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290103(.x(x_103), .z(tmp00_103_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290104(.x(x_104), .z(tmp00_104_29));
	booth_0006 #(.WIDTH(WIDTH)) mul00290105(.x(x_105), .z(tmp00_105_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290106(.x(x_106), .z(tmp00_106_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290107(.x(x_107), .z(tmp00_107_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290108(.x(x_108), .z(tmp00_108_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290109(.x(x_109), .z(tmp00_109_29));
	booth__010 #(.WIDTH(WIDTH)) mul00290110(.x(x_110), .z(tmp00_110_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290111(.x(x_111), .z(tmp00_111_29));
	booth_0006 #(.WIDTH(WIDTH)) mul00290112(.x(x_112), .z(tmp00_112_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00290113(.x(x_113), .z(tmp00_113_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290114(.x(x_114), .z(tmp00_114_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290115(.x(x_115), .z(tmp00_115_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290116(.x(x_116), .z(tmp00_116_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290117(.x(x_117), .z(tmp00_117_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290118(.x(x_118), .z(tmp00_118_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290119(.x(x_119), .z(tmp00_119_29));
	booth_0004 #(.WIDTH(WIDTH)) mul00290120(.x(x_120), .z(tmp00_120_29));
	booth_0000 #(.WIDTH(WIDTH)) mul00290121(.x(x_121), .z(tmp00_121_29));
	booth_0006 #(.WIDTH(WIDTH)) mul00290122(.x(x_122), .z(tmp00_122_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290123(.x(x_123), .z(tmp00_123_29));
	booth__008 #(.WIDTH(WIDTH)) mul00290124(.x(x_124), .z(tmp00_124_29));
	booth_0010 #(.WIDTH(WIDTH)) mul00290125(.x(x_125), .z(tmp00_125_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290126(.x(x_126), .z(tmp00_126_29));
	booth__004 #(.WIDTH(WIDTH)) mul00290127(.x(x_127), .z(tmp00_127_29));
	booth_0008 #(.WIDTH(WIDTH)) mul00300000(.x(x_0), .z(tmp00_0_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300001(.x(x_1), .z(tmp00_1_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300002(.x(x_2), .z(tmp00_2_30));
	booth__010 #(.WIDTH(WIDTH)) mul00300003(.x(x_3), .z(tmp00_3_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300004(.x(x_4), .z(tmp00_4_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300005(.x(x_5), .z(tmp00_5_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300006(.x(x_6), .z(tmp00_6_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300007(.x(x_7), .z(tmp00_7_30));
	booth__012 #(.WIDTH(WIDTH)) mul00300008(.x(x_8), .z(tmp00_8_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300009(.x(x_9), .z(tmp00_9_30));
	booth_0006 #(.WIDTH(WIDTH)) mul00300010(.x(x_10), .z(tmp00_10_30));
	booth_0010 #(.WIDTH(WIDTH)) mul00300011(.x(x_11), .z(tmp00_11_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300012(.x(x_12), .z(tmp00_12_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300013(.x(x_13), .z(tmp00_13_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300014(.x(x_14), .z(tmp00_14_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300015(.x(x_15), .z(tmp00_15_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300016(.x(x_16), .z(tmp00_16_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300017(.x(x_17), .z(tmp00_17_30));
	booth__004 #(.WIDTH(WIDTH)) mul00300018(.x(x_18), .z(tmp00_18_30));
	booth__012 #(.WIDTH(WIDTH)) mul00300019(.x(x_19), .z(tmp00_19_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300020(.x(x_20), .z(tmp00_20_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300021(.x(x_21), .z(tmp00_21_30));
	booth_0016 #(.WIDTH(WIDTH)) mul00300022(.x(x_22), .z(tmp00_22_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300023(.x(x_23), .z(tmp00_23_30));
	booth__002 #(.WIDTH(WIDTH)) mul00300024(.x(x_24), .z(tmp00_24_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300025(.x(x_25), .z(tmp00_25_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300026(.x(x_26), .z(tmp00_26_30));
	booth__004 #(.WIDTH(WIDTH)) mul00300027(.x(x_27), .z(tmp00_27_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300028(.x(x_28), .z(tmp00_28_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300029(.x(x_29), .z(tmp00_29_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300030(.x(x_30), .z(tmp00_30_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300031(.x(x_31), .z(tmp00_31_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300032(.x(x_32), .z(tmp00_32_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300033(.x(x_33), .z(tmp00_33_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300034(.x(x_34), .z(tmp00_34_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300035(.x(x_35), .z(tmp00_35_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300036(.x(x_36), .z(tmp00_36_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300037(.x(x_37), .z(tmp00_37_30));
	booth__016 #(.WIDTH(WIDTH)) mul00300038(.x(x_38), .z(tmp00_38_30));
	booth_0024 #(.WIDTH(WIDTH)) mul00300039(.x(x_39), .z(tmp00_39_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300040(.x(x_40), .z(tmp00_40_30));
	booth__012 #(.WIDTH(WIDTH)) mul00300041(.x(x_41), .z(tmp00_41_30));
	booth_0020 #(.WIDTH(WIDTH)) mul00300042(.x(x_42), .z(tmp00_42_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300043(.x(x_43), .z(tmp00_43_30));
	booth_0012 #(.WIDTH(WIDTH)) mul00300044(.x(x_44), .z(tmp00_44_30));
	booth_0006 #(.WIDTH(WIDTH)) mul00300045(.x(x_45), .z(tmp00_45_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300046(.x(x_46), .z(tmp00_46_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300047(.x(x_47), .z(tmp00_47_30));
	booth_0016 #(.WIDTH(WIDTH)) mul00300048(.x(x_48), .z(tmp00_48_30));
	booth__006 #(.WIDTH(WIDTH)) mul00300049(.x(x_49), .z(tmp00_49_30));
	booth__006 #(.WIDTH(WIDTH)) mul00300050(.x(x_50), .z(tmp00_50_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300051(.x(x_51), .z(tmp00_51_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300052(.x(x_52), .z(tmp00_52_30));
	booth_0012 #(.WIDTH(WIDTH)) mul00300053(.x(x_53), .z(tmp00_53_30));
	booth_0016 #(.WIDTH(WIDTH)) mul00300054(.x(x_54), .z(tmp00_54_30));
	booth__012 #(.WIDTH(WIDTH)) mul00300055(.x(x_55), .z(tmp00_55_30));
	booth_0016 #(.WIDTH(WIDTH)) mul00300056(.x(x_56), .z(tmp00_56_30));
	booth_0006 #(.WIDTH(WIDTH)) mul00300057(.x(x_57), .z(tmp00_57_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300058(.x(x_58), .z(tmp00_58_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300059(.x(x_59), .z(tmp00_59_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300060(.x(x_60), .z(tmp00_60_30));
	booth_0012 #(.WIDTH(WIDTH)) mul00300061(.x(x_61), .z(tmp00_61_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300062(.x(x_62), .z(tmp00_62_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300063(.x(x_63), .z(tmp00_63_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300064(.x(x_64), .z(tmp00_64_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300065(.x(x_65), .z(tmp00_65_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300066(.x(x_66), .z(tmp00_66_30));
	booth__004 #(.WIDTH(WIDTH)) mul00300067(.x(x_67), .z(tmp00_67_30));
	booth_0012 #(.WIDTH(WIDTH)) mul00300068(.x(x_68), .z(tmp00_68_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300069(.x(x_69), .z(tmp00_69_30));
	booth__004 #(.WIDTH(WIDTH)) mul00300070(.x(x_70), .z(tmp00_70_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300071(.x(x_71), .z(tmp00_71_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300072(.x(x_72), .z(tmp00_72_30));
	booth__006 #(.WIDTH(WIDTH)) mul00300073(.x(x_73), .z(tmp00_73_30));
	booth_0006 #(.WIDTH(WIDTH)) mul00300074(.x(x_74), .z(tmp00_74_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300075(.x(x_75), .z(tmp00_75_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300076(.x(x_76), .z(tmp00_76_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300077(.x(x_77), .z(tmp00_77_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300078(.x(x_78), .z(tmp00_78_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300079(.x(x_79), .z(tmp00_79_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300080(.x(x_80), .z(tmp00_80_30));
	booth_0010 #(.WIDTH(WIDTH)) mul00300081(.x(x_81), .z(tmp00_81_30));
	booth_0012 #(.WIDTH(WIDTH)) mul00300082(.x(x_82), .z(tmp00_82_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300083(.x(x_83), .z(tmp00_83_30));
	booth_0006 #(.WIDTH(WIDTH)) mul00300084(.x(x_84), .z(tmp00_84_30));
	booth_0014 #(.WIDTH(WIDTH)) mul00300085(.x(x_85), .z(tmp00_85_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300086(.x(x_86), .z(tmp00_86_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300087(.x(x_87), .z(tmp00_87_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300088(.x(x_88), .z(tmp00_88_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300089(.x(x_89), .z(tmp00_89_30));
	booth_0024 #(.WIDTH(WIDTH)) mul00300090(.x(x_90), .z(tmp00_90_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300091(.x(x_91), .z(tmp00_91_30));
	booth_0012 #(.WIDTH(WIDTH)) mul00300092(.x(x_92), .z(tmp00_92_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300093(.x(x_93), .z(tmp00_93_30));
	booth__012 #(.WIDTH(WIDTH)) mul00300094(.x(x_94), .z(tmp00_94_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300095(.x(x_95), .z(tmp00_95_30));
	booth__012 #(.WIDTH(WIDTH)) mul00300096(.x(x_96), .z(tmp00_96_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300097(.x(x_97), .z(tmp00_97_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300098(.x(x_98), .z(tmp00_98_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300099(.x(x_99), .z(tmp00_99_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300100(.x(x_100), .z(tmp00_100_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300101(.x(x_101), .z(tmp00_101_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300102(.x(x_102), .z(tmp00_102_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300103(.x(x_103), .z(tmp00_103_30));
	booth__004 #(.WIDTH(WIDTH)) mul00300104(.x(x_104), .z(tmp00_104_30));
	booth__004 #(.WIDTH(WIDTH)) mul00300105(.x(x_105), .z(tmp00_105_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300106(.x(x_106), .z(tmp00_106_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300107(.x(x_107), .z(tmp00_107_30));
	booth_0012 #(.WIDTH(WIDTH)) mul00300108(.x(x_108), .z(tmp00_108_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300109(.x(x_109), .z(tmp00_109_30));
	booth__014 #(.WIDTH(WIDTH)) mul00300110(.x(x_110), .z(tmp00_110_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300111(.x(x_111), .z(tmp00_111_30));
	booth_0006 #(.WIDTH(WIDTH)) mul00300112(.x(x_112), .z(tmp00_112_30));
	booth_0018 #(.WIDTH(WIDTH)) mul00300113(.x(x_113), .z(tmp00_113_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300114(.x(x_114), .z(tmp00_114_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300115(.x(x_115), .z(tmp00_115_30));
	booth__002 #(.WIDTH(WIDTH)) mul00300116(.x(x_116), .z(tmp00_116_30));
	booth__010 #(.WIDTH(WIDTH)) mul00300117(.x(x_117), .z(tmp00_117_30));
	booth_0000 #(.WIDTH(WIDTH)) mul00300118(.x(x_118), .z(tmp00_118_30));
	booth_0006 #(.WIDTH(WIDTH)) mul00300119(.x(x_119), .z(tmp00_119_30));
	booth_0018 #(.WIDTH(WIDTH)) mul00300120(.x(x_120), .z(tmp00_120_30));
	booth__014 #(.WIDTH(WIDTH)) mul00300121(.x(x_121), .z(tmp00_121_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300122(.x(x_122), .z(tmp00_122_30));
	booth__008 #(.WIDTH(WIDTH)) mul00300123(.x(x_123), .z(tmp00_123_30));
	booth__012 #(.WIDTH(WIDTH)) mul00300124(.x(x_124), .z(tmp00_124_30));
	booth_0004 #(.WIDTH(WIDTH)) mul00300125(.x(x_125), .z(tmp00_125_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00300126(.x(x_126), .z(tmp00_126_30));
	booth__004 #(.WIDTH(WIDTH)) mul00300127(.x(x_127), .z(tmp00_127_30));
	booth_0008 #(.WIDTH(WIDTH)) mul00310000(.x(x_0), .z(tmp00_0_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310001(.x(x_1), .z(tmp00_1_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310002(.x(x_2), .z(tmp00_2_31));
	booth__002 #(.WIDTH(WIDTH)) mul00310003(.x(x_3), .z(tmp00_3_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310004(.x(x_4), .z(tmp00_4_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310005(.x(x_5), .z(tmp00_5_31));
	booth_0006 #(.WIDTH(WIDTH)) mul00310006(.x(x_6), .z(tmp00_6_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310007(.x(x_7), .z(tmp00_7_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310008(.x(x_8), .z(tmp00_8_31));
	booth__010 #(.WIDTH(WIDTH)) mul00310009(.x(x_9), .z(tmp00_9_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310010(.x(x_10), .z(tmp00_10_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310011(.x(x_11), .z(tmp00_11_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310012(.x(x_12), .z(tmp00_12_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310013(.x(x_13), .z(tmp00_13_31));
	booth_0002 #(.WIDTH(WIDTH)) mul00310014(.x(x_14), .z(tmp00_14_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310015(.x(x_15), .z(tmp00_15_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310016(.x(x_16), .z(tmp00_16_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310017(.x(x_17), .z(tmp00_17_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310018(.x(x_18), .z(tmp00_18_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310019(.x(x_19), .z(tmp00_19_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310020(.x(x_20), .z(tmp00_20_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310021(.x(x_21), .z(tmp00_21_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310022(.x(x_22), .z(tmp00_22_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310023(.x(x_23), .z(tmp00_23_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310024(.x(x_24), .z(tmp00_24_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310025(.x(x_25), .z(tmp00_25_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310026(.x(x_26), .z(tmp00_26_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310027(.x(x_27), .z(tmp00_27_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310028(.x(x_28), .z(tmp00_28_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310029(.x(x_29), .z(tmp00_29_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310030(.x(x_30), .z(tmp00_30_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310031(.x(x_31), .z(tmp00_31_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310032(.x(x_32), .z(tmp00_32_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310033(.x(x_33), .z(tmp00_33_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310034(.x(x_34), .z(tmp00_34_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310035(.x(x_35), .z(tmp00_35_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310036(.x(x_36), .z(tmp00_36_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310037(.x(x_37), .z(tmp00_37_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310038(.x(x_38), .z(tmp00_38_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310039(.x(x_39), .z(tmp00_39_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310040(.x(x_40), .z(tmp00_40_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310041(.x(x_41), .z(tmp00_41_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310042(.x(x_42), .z(tmp00_42_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310043(.x(x_43), .z(tmp00_43_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310044(.x(x_44), .z(tmp00_44_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310045(.x(x_45), .z(tmp00_45_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310046(.x(x_46), .z(tmp00_46_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310047(.x(x_47), .z(tmp00_47_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310048(.x(x_48), .z(tmp00_48_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310049(.x(x_49), .z(tmp00_49_31));
	booth_0006 #(.WIDTH(WIDTH)) mul00310050(.x(x_50), .z(tmp00_50_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310051(.x(x_51), .z(tmp00_51_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310052(.x(x_52), .z(tmp00_52_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310053(.x(x_53), .z(tmp00_53_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310054(.x(x_54), .z(tmp00_54_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310055(.x(x_55), .z(tmp00_55_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310056(.x(x_56), .z(tmp00_56_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310057(.x(x_57), .z(tmp00_57_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310058(.x(x_58), .z(tmp00_58_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310059(.x(x_59), .z(tmp00_59_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310060(.x(x_60), .z(tmp00_60_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310061(.x(x_61), .z(tmp00_61_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310062(.x(x_62), .z(tmp00_62_31));
	booth__010 #(.WIDTH(WIDTH)) mul00310063(.x(x_63), .z(tmp00_63_31));
	booth_0002 #(.WIDTH(WIDTH)) mul00310064(.x(x_64), .z(tmp00_64_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310065(.x(x_65), .z(tmp00_65_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310066(.x(x_66), .z(tmp00_66_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310067(.x(x_67), .z(tmp00_67_31));
	booth__010 #(.WIDTH(WIDTH)) mul00310068(.x(x_68), .z(tmp00_68_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310069(.x(x_69), .z(tmp00_69_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310070(.x(x_70), .z(tmp00_70_31));
	booth_0010 #(.WIDTH(WIDTH)) mul00310071(.x(x_71), .z(tmp00_71_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310072(.x(x_72), .z(tmp00_72_31));
	booth__002 #(.WIDTH(WIDTH)) mul00310073(.x(x_73), .z(tmp00_73_31));
	booth__010 #(.WIDTH(WIDTH)) mul00310074(.x(x_74), .z(tmp00_74_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310075(.x(x_75), .z(tmp00_75_31));
	booth_0010 #(.WIDTH(WIDTH)) mul00310076(.x(x_76), .z(tmp00_76_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310077(.x(x_77), .z(tmp00_77_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310078(.x(x_78), .z(tmp00_78_31));
	booth__002 #(.WIDTH(WIDTH)) mul00310079(.x(x_79), .z(tmp00_79_31));
	booth__010 #(.WIDTH(WIDTH)) mul00310080(.x(x_80), .z(tmp00_80_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310081(.x(x_81), .z(tmp00_81_31));
	booth__012 #(.WIDTH(WIDTH)) mul00310082(.x(x_82), .z(tmp00_82_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310083(.x(x_83), .z(tmp00_83_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310084(.x(x_84), .z(tmp00_84_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310085(.x(x_85), .z(tmp00_85_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310086(.x(x_86), .z(tmp00_86_31));
	booth_0010 #(.WIDTH(WIDTH)) mul00310087(.x(x_87), .z(tmp00_87_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310088(.x(x_88), .z(tmp00_88_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310089(.x(x_89), .z(tmp00_89_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310090(.x(x_90), .z(tmp00_90_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310091(.x(x_91), .z(tmp00_91_31));
	booth__010 #(.WIDTH(WIDTH)) mul00310092(.x(x_92), .z(tmp00_92_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310093(.x(x_93), .z(tmp00_93_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310094(.x(x_94), .z(tmp00_94_31));
	booth__006 #(.WIDTH(WIDTH)) mul00310095(.x(x_95), .z(tmp00_95_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310096(.x(x_96), .z(tmp00_96_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310097(.x(x_97), .z(tmp00_97_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310098(.x(x_98), .z(tmp00_98_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310099(.x(x_99), .z(tmp00_99_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310100(.x(x_100), .z(tmp00_100_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310101(.x(x_101), .z(tmp00_101_31));
	booth__002 #(.WIDTH(WIDTH)) mul00310102(.x(x_102), .z(tmp00_102_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310103(.x(x_103), .z(tmp00_103_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310104(.x(x_104), .z(tmp00_104_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310105(.x(x_105), .z(tmp00_105_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310106(.x(x_106), .z(tmp00_106_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310107(.x(x_107), .z(tmp00_107_31));
	booth_0012 #(.WIDTH(WIDTH)) mul00310108(.x(x_108), .z(tmp00_108_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310109(.x(x_109), .z(tmp00_109_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310110(.x(x_110), .z(tmp00_110_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310111(.x(x_111), .z(tmp00_111_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310112(.x(x_112), .z(tmp00_112_31));
	booth__008 #(.WIDTH(WIDTH)) mul00310113(.x(x_113), .z(tmp00_113_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310114(.x(x_114), .z(tmp00_114_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310115(.x(x_115), .z(tmp00_115_31));
	booth_0010 #(.WIDTH(WIDTH)) mul00310116(.x(x_116), .z(tmp00_116_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310117(.x(x_117), .z(tmp00_117_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310118(.x(x_118), .z(tmp00_118_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310119(.x(x_119), .z(tmp00_119_31));
	booth_0004 #(.WIDTH(WIDTH)) mul00310120(.x(x_120), .z(tmp00_120_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310121(.x(x_121), .z(tmp00_121_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310122(.x(x_122), .z(tmp00_122_31));
	booth_0008 #(.WIDTH(WIDTH)) mul00310123(.x(x_123), .z(tmp00_123_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310124(.x(x_124), .z(tmp00_124_31));
	booth_0000 #(.WIDTH(WIDTH)) mul00310125(.x(x_125), .z(tmp00_125_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310126(.x(x_126), .z(tmp00_126_31));
	booth__004 #(.WIDTH(WIDTH)) mul00310127(.x(x_127), .z(tmp00_127_31));
	booth__010 #(.WIDTH(WIDTH)) mul00320000(.x(x_0), .z(tmp00_0_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320001(.x(x_1), .z(tmp00_1_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320002(.x(x_2), .z(tmp00_2_32));
	booth_0002 #(.WIDTH(WIDTH)) mul00320003(.x(x_3), .z(tmp00_3_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320004(.x(x_4), .z(tmp00_4_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320005(.x(x_5), .z(tmp00_5_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320006(.x(x_6), .z(tmp00_6_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320007(.x(x_7), .z(tmp00_7_32));
	booth__010 #(.WIDTH(WIDTH)) mul00320008(.x(x_8), .z(tmp00_8_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320009(.x(x_9), .z(tmp00_9_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320010(.x(x_10), .z(tmp00_10_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320011(.x(x_11), .z(tmp00_11_32));
	booth_0010 #(.WIDTH(WIDTH)) mul00320012(.x(x_12), .z(tmp00_12_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320013(.x(x_13), .z(tmp00_13_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320014(.x(x_14), .z(tmp00_14_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320015(.x(x_15), .z(tmp00_15_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320016(.x(x_16), .z(tmp00_16_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320017(.x(x_17), .z(tmp00_17_32));
	booth__002 #(.WIDTH(WIDTH)) mul00320018(.x(x_18), .z(tmp00_18_32));
	booth_0002 #(.WIDTH(WIDTH)) mul00320019(.x(x_19), .z(tmp00_19_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320020(.x(x_20), .z(tmp00_20_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320021(.x(x_21), .z(tmp00_21_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320022(.x(x_22), .z(tmp00_22_32));
	booth__006 #(.WIDTH(WIDTH)) mul00320023(.x(x_23), .z(tmp00_23_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320024(.x(x_24), .z(tmp00_24_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320025(.x(x_25), .z(tmp00_25_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320026(.x(x_26), .z(tmp00_26_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320027(.x(x_27), .z(tmp00_27_32));
	booth_0006 #(.WIDTH(WIDTH)) mul00320028(.x(x_28), .z(tmp00_28_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320029(.x(x_29), .z(tmp00_29_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320030(.x(x_30), .z(tmp00_30_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320031(.x(x_31), .z(tmp00_31_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320032(.x(x_32), .z(tmp00_32_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320033(.x(x_33), .z(tmp00_33_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320034(.x(x_34), .z(tmp00_34_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320035(.x(x_35), .z(tmp00_35_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320036(.x(x_36), .z(tmp00_36_32));
	booth__010 #(.WIDTH(WIDTH)) mul00320037(.x(x_37), .z(tmp00_37_32));
	booth__014 #(.WIDTH(WIDTH)) mul00320038(.x(x_38), .z(tmp00_38_32));
	booth_0016 #(.WIDTH(WIDTH)) mul00320039(.x(x_39), .z(tmp00_39_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320040(.x(x_40), .z(tmp00_40_32));
	booth__010 #(.WIDTH(WIDTH)) mul00320041(.x(x_41), .z(tmp00_41_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320042(.x(x_42), .z(tmp00_42_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320043(.x(x_43), .z(tmp00_43_32));
	booth_0010 #(.WIDTH(WIDTH)) mul00320044(.x(x_44), .z(tmp00_44_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320045(.x(x_45), .z(tmp00_45_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320046(.x(x_46), .z(tmp00_46_32));
	booth__002 #(.WIDTH(WIDTH)) mul00320047(.x(x_47), .z(tmp00_47_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320048(.x(x_48), .z(tmp00_48_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320049(.x(x_49), .z(tmp00_49_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320050(.x(x_50), .z(tmp00_50_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320051(.x(x_51), .z(tmp00_51_32));
	booth__010 #(.WIDTH(WIDTH)) mul00320052(.x(x_52), .z(tmp00_52_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320053(.x(x_53), .z(tmp00_53_32));
	booth_0012 #(.WIDTH(WIDTH)) mul00320054(.x(x_54), .z(tmp00_54_32));
	booth__002 #(.WIDTH(WIDTH)) mul00320055(.x(x_55), .z(tmp00_55_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320056(.x(x_56), .z(tmp00_56_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320057(.x(x_57), .z(tmp00_57_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320058(.x(x_58), .z(tmp00_58_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320059(.x(x_59), .z(tmp00_59_32));
	booth_0010 #(.WIDTH(WIDTH)) mul00320060(.x(x_60), .z(tmp00_60_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320061(.x(x_61), .z(tmp00_61_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320062(.x(x_62), .z(tmp00_62_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320063(.x(x_63), .z(tmp00_63_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320064(.x(x_64), .z(tmp00_64_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320065(.x(x_65), .z(tmp00_65_32));
	booth_0002 #(.WIDTH(WIDTH)) mul00320066(.x(x_66), .z(tmp00_66_32));
	booth__010 #(.WIDTH(WIDTH)) mul00320067(.x(x_67), .z(tmp00_67_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320068(.x(x_68), .z(tmp00_68_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320069(.x(x_69), .z(tmp00_69_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320070(.x(x_70), .z(tmp00_70_32));
	booth_0010 #(.WIDTH(WIDTH)) mul00320071(.x(x_71), .z(tmp00_71_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320072(.x(x_72), .z(tmp00_72_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320073(.x(x_73), .z(tmp00_73_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320074(.x(x_74), .z(tmp00_74_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320075(.x(x_75), .z(tmp00_75_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320076(.x(x_76), .z(tmp00_76_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320077(.x(x_77), .z(tmp00_77_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320078(.x(x_78), .z(tmp00_78_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320079(.x(x_79), .z(tmp00_79_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320080(.x(x_80), .z(tmp00_80_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320081(.x(x_81), .z(tmp00_81_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320082(.x(x_82), .z(tmp00_82_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320083(.x(x_83), .z(tmp00_83_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320084(.x(x_84), .z(tmp00_84_32));
	booth_0010 #(.WIDTH(WIDTH)) mul00320085(.x(x_85), .z(tmp00_85_32));
	booth__010 #(.WIDTH(WIDTH)) mul00320086(.x(x_86), .z(tmp00_86_32));
	booth_0012 #(.WIDTH(WIDTH)) mul00320087(.x(x_87), .z(tmp00_87_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320088(.x(x_88), .z(tmp00_88_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320089(.x(x_89), .z(tmp00_89_32));
	booth_0006 #(.WIDTH(WIDTH)) mul00320090(.x(x_90), .z(tmp00_90_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320091(.x(x_91), .z(tmp00_91_32));
	booth_0006 #(.WIDTH(WIDTH)) mul00320092(.x(x_92), .z(tmp00_92_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320093(.x(x_93), .z(tmp00_93_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320094(.x(x_94), .z(tmp00_94_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320095(.x(x_95), .z(tmp00_95_32));
	booth_0012 #(.WIDTH(WIDTH)) mul00320096(.x(x_96), .z(tmp00_96_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320097(.x(x_97), .z(tmp00_97_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320098(.x(x_98), .z(tmp00_98_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320099(.x(x_99), .z(tmp00_99_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320100(.x(x_100), .z(tmp00_100_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320101(.x(x_101), .z(tmp00_101_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320102(.x(x_102), .z(tmp00_102_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320103(.x(x_103), .z(tmp00_103_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320104(.x(x_104), .z(tmp00_104_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320105(.x(x_105), .z(tmp00_105_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320106(.x(x_106), .z(tmp00_106_32));
	booth_0010 #(.WIDTH(WIDTH)) mul00320107(.x(x_107), .z(tmp00_107_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320108(.x(x_108), .z(tmp00_108_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320109(.x(x_109), .z(tmp00_109_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320110(.x(x_110), .z(tmp00_110_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320111(.x(x_111), .z(tmp00_111_32));
	booth__002 #(.WIDTH(WIDTH)) mul00320112(.x(x_112), .z(tmp00_112_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320113(.x(x_113), .z(tmp00_113_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320114(.x(x_114), .z(tmp00_114_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320115(.x(x_115), .z(tmp00_115_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320116(.x(x_116), .z(tmp00_116_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320117(.x(x_117), .z(tmp00_117_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00320118(.x(x_118), .z(tmp00_118_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320119(.x(x_119), .z(tmp00_119_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320120(.x(x_120), .z(tmp00_120_32));
	booth__004 #(.WIDTH(WIDTH)) mul00320121(.x(x_121), .z(tmp00_121_32));
	booth__008 #(.WIDTH(WIDTH)) mul00320122(.x(x_122), .z(tmp00_122_32));
	booth_0000 #(.WIDTH(WIDTH)) mul00320123(.x(x_123), .z(tmp00_123_32));
	booth_0010 #(.WIDTH(WIDTH)) mul00320124(.x(x_124), .z(tmp00_124_32));
	booth__002 #(.WIDTH(WIDTH)) mul00320125(.x(x_125), .z(tmp00_125_32));
	booth_0008 #(.WIDTH(WIDTH)) mul00320126(.x(x_126), .z(tmp00_126_32));
	booth_0002 #(.WIDTH(WIDTH)) mul00320127(.x(x_127), .z(tmp00_127_32));
	booth_0004 #(.WIDTH(WIDTH)) mul00330000(.x(x_0), .z(tmp00_0_33));
	booth__002 #(.WIDTH(WIDTH)) mul00330001(.x(x_1), .z(tmp00_1_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330002(.x(x_2), .z(tmp00_2_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330003(.x(x_3), .z(tmp00_3_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330004(.x(x_4), .z(tmp00_4_33));
	booth_0010 #(.WIDTH(WIDTH)) mul00330005(.x(x_5), .z(tmp00_5_33));
	booth__004 #(.WIDTH(WIDTH)) mul00330006(.x(x_6), .z(tmp00_6_33));
	booth__004 #(.WIDTH(WIDTH)) mul00330007(.x(x_7), .z(tmp00_7_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330008(.x(x_8), .z(tmp00_8_33));
	booth_0002 #(.WIDTH(WIDTH)) mul00330009(.x(x_9), .z(tmp00_9_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330010(.x(x_10), .z(tmp00_10_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330011(.x(x_11), .z(tmp00_11_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330012(.x(x_12), .z(tmp00_12_33));
	booth_0016 #(.WIDTH(WIDTH)) mul00330013(.x(x_13), .z(tmp00_13_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330014(.x(x_14), .z(tmp00_14_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330015(.x(x_15), .z(tmp00_15_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330016(.x(x_16), .z(tmp00_16_33));
	booth_0012 #(.WIDTH(WIDTH)) mul00330017(.x(x_17), .z(tmp00_17_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330018(.x(x_18), .z(tmp00_18_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330019(.x(x_19), .z(tmp00_19_33));
	booth_0016 #(.WIDTH(WIDTH)) mul00330020(.x(x_20), .z(tmp00_20_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330021(.x(x_21), .z(tmp00_21_33));
	booth_0010 #(.WIDTH(WIDTH)) mul00330022(.x(x_22), .z(tmp00_22_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330023(.x(x_23), .z(tmp00_23_33));
	booth_0010 #(.WIDTH(WIDTH)) mul00330024(.x(x_24), .z(tmp00_24_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330025(.x(x_25), .z(tmp00_25_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330026(.x(x_26), .z(tmp00_26_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330027(.x(x_27), .z(tmp00_27_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330028(.x(x_28), .z(tmp00_28_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330029(.x(x_29), .z(tmp00_29_33));
	booth_0012 #(.WIDTH(WIDTH)) mul00330030(.x(x_30), .z(tmp00_30_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330031(.x(x_31), .z(tmp00_31_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330032(.x(x_32), .z(tmp00_32_33));
	booth__010 #(.WIDTH(WIDTH)) mul00330033(.x(x_33), .z(tmp00_33_33));
	booth__006 #(.WIDTH(WIDTH)) mul00330034(.x(x_34), .z(tmp00_34_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330035(.x(x_35), .z(tmp00_35_33));
	booth__002 #(.WIDTH(WIDTH)) mul00330036(.x(x_36), .z(tmp00_36_33));
	booth__012 #(.WIDTH(WIDTH)) mul00330037(.x(x_37), .z(tmp00_37_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330038(.x(x_38), .z(tmp00_38_33));
	booth_0024 #(.WIDTH(WIDTH)) mul00330039(.x(x_39), .z(tmp00_39_33));
	booth__010 #(.WIDTH(WIDTH)) mul00330040(.x(x_40), .z(tmp00_40_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330041(.x(x_41), .z(tmp00_41_33));
	booth__010 #(.WIDTH(WIDTH)) mul00330042(.x(x_42), .z(tmp00_42_33));
	booth__006 #(.WIDTH(WIDTH)) mul00330043(.x(x_43), .z(tmp00_43_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330044(.x(x_44), .z(tmp00_44_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330045(.x(x_45), .z(tmp00_45_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330046(.x(x_46), .z(tmp00_46_33));
	booth__016 #(.WIDTH(WIDTH)) mul00330047(.x(x_47), .z(tmp00_47_33));
	booth_0010 #(.WIDTH(WIDTH)) mul00330048(.x(x_48), .z(tmp00_48_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330049(.x(x_49), .z(tmp00_49_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330050(.x(x_50), .z(tmp00_50_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330051(.x(x_51), .z(tmp00_51_33));
	booth__006 #(.WIDTH(WIDTH)) mul00330052(.x(x_52), .z(tmp00_52_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330053(.x(x_53), .z(tmp00_53_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330054(.x(x_54), .z(tmp00_54_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330055(.x(x_55), .z(tmp00_55_33));
	booth__004 #(.WIDTH(WIDTH)) mul00330056(.x(x_56), .z(tmp00_56_33));
	booth_0006 #(.WIDTH(WIDTH)) mul00330057(.x(x_57), .z(tmp00_57_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330058(.x(x_58), .z(tmp00_58_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330059(.x(x_59), .z(tmp00_59_33));
	booth__004 #(.WIDTH(WIDTH)) mul00330060(.x(x_60), .z(tmp00_60_33));
	booth__004 #(.WIDTH(WIDTH)) mul00330061(.x(x_61), .z(tmp00_61_33));
	booth__006 #(.WIDTH(WIDTH)) mul00330062(.x(x_62), .z(tmp00_62_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330063(.x(x_63), .z(tmp00_63_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330064(.x(x_64), .z(tmp00_64_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330065(.x(x_65), .z(tmp00_65_33));
	booth__004 #(.WIDTH(WIDTH)) mul00330066(.x(x_66), .z(tmp00_66_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330067(.x(x_67), .z(tmp00_67_33));
	booth_0016 #(.WIDTH(WIDTH)) mul00330068(.x(x_68), .z(tmp00_68_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330069(.x(x_69), .z(tmp00_69_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330070(.x(x_70), .z(tmp00_70_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330071(.x(x_71), .z(tmp00_71_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330072(.x(x_72), .z(tmp00_72_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330073(.x(x_73), .z(tmp00_73_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330074(.x(x_74), .z(tmp00_74_33));
	booth_0016 #(.WIDTH(WIDTH)) mul00330075(.x(x_75), .z(tmp00_75_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330076(.x(x_76), .z(tmp00_76_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330077(.x(x_77), .z(tmp00_77_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330078(.x(x_78), .z(tmp00_78_33));
	booth_0010 #(.WIDTH(WIDTH)) mul00330079(.x(x_79), .z(tmp00_79_33));
	booth__012 #(.WIDTH(WIDTH)) mul00330080(.x(x_80), .z(tmp00_80_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330081(.x(x_81), .z(tmp00_81_33));
	booth__012 #(.WIDTH(WIDTH)) mul00330082(.x(x_82), .z(tmp00_82_33));
	booth__006 #(.WIDTH(WIDTH)) mul00330083(.x(x_83), .z(tmp00_83_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330084(.x(x_84), .z(tmp00_84_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330085(.x(x_85), .z(tmp00_85_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330086(.x(x_86), .z(tmp00_86_33));
	booth_0012 #(.WIDTH(WIDTH)) mul00330087(.x(x_87), .z(tmp00_87_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330088(.x(x_88), .z(tmp00_88_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330089(.x(x_89), .z(tmp00_89_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330090(.x(x_90), .z(tmp00_90_33));
	booth_0010 #(.WIDTH(WIDTH)) mul00330091(.x(x_91), .z(tmp00_91_33));
	booth_0010 #(.WIDTH(WIDTH)) mul00330092(.x(x_92), .z(tmp00_92_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330093(.x(x_93), .z(tmp00_93_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330094(.x(x_94), .z(tmp00_94_33));
	booth__010 #(.WIDTH(WIDTH)) mul00330095(.x(x_95), .z(tmp00_95_33));
	booth_0016 #(.WIDTH(WIDTH)) mul00330096(.x(x_96), .z(tmp00_96_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330097(.x(x_97), .z(tmp00_97_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330098(.x(x_98), .z(tmp00_98_33));
	booth_0002 #(.WIDTH(WIDTH)) mul00330099(.x(x_99), .z(tmp00_99_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330100(.x(x_100), .z(tmp00_100_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330101(.x(x_101), .z(tmp00_101_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330102(.x(x_102), .z(tmp00_102_33));
	booth__010 #(.WIDTH(WIDTH)) mul00330103(.x(x_103), .z(tmp00_103_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330104(.x(x_104), .z(tmp00_104_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330105(.x(x_105), .z(tmp00_105_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330106(.x(x_106), .z(tmp00_106_33));
	booth__002 #(.WIDTH(WIDTH)) mul00330107(.x(x_107), .z(tmp00_107_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330108(.x(x_108), .z(tmp00_108_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330109(.x(x_109), .z(tmp00_109_33));
	booth_0014 #(.WIDTH(WIDTH)) mul00330110(.x(x_110), .z(tmp00_110_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330111(.x(x_111), .z(tmp00_111_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330112(.x(x_112), .z(tmp00_112_33));
	booth__012 #(.WIDTH(WIDTH)) mul00330113(.x(x_113), .z(tmp00_113_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330114(.x(x_114), .z(tmp00_114_33));
	booth__016 #(.WIDTH(WIDTH)) mul00330115(.x(x_115), .z(tmp00_115_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330116(.x(x_116), .z(tmp00_116_33));
	booth__004 #(.WIDTH(WIDTH)) mul00330117(.x(x_117), .z(tmp00_117_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330118(.x(x_118), .z(tmp00_118_33));
	booth__010 #(.WIDTH(WIDTH)) mul00330119(.x(x_119), .z(tmp00_119_33));
	booth_0016 #(.WIDTH(WIDTH)) mul00330120(.x(x_120), .z(tmp00_120_33));
	booth__016 #(.WIDTH(WIDTH)) mul00330121(.x(x_121), .z(tmp00_121_33));
	booth_0008 #(.WIDTH(WIDTH)) mul00330122(.x(x_122), .z(tmp00_122_33));
	booth__012 #(.WIDTH(WIDTH)) mul00330123(.x(x_123), .z(tmp00_123_33));
	booth_0000 #(.WIDTH(WIDTH)) mul00330124(.x(x_124), .z(tmp00_124_33));
	booth_0004 #(.WIDTH(WIDTH)) mul00330125(.x(x_125), .z(tmp00_125_33));
	booth__008 #(.WIDTH(WIDTH)) mul00330126(.x(x_126), .z(tmp00_126_33));
	booth_0014 #(.WIDTH(WIDTH)) mul00330127(.x(x_127), .z(tmp00_127_33));
	booth_0002 #(.WIDTH(WIDTH)) mul00340000(.x(x_0), .z(tmp00_0_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340001(.x(x_1), .z(tmp00_1_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340002(.x(x_2), .z(tmp00_2_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340003(.x(x_3), .z(tmp00_3_34));
	booth__006 #(.WIDTH(WIDTH)) mul00340004(.x(x_4), .z(tmp00_4_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340005(.x(x_5), .z(tmp00_5_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340006(.x(x_6), .z(tmp00_6_34));
	booth__010 #(.WIDTH(WIDTH)) mul00340007(.x(x_7), .z(tmp00_7_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340008(.x(x_8), .z(tmp00_8_34));
	booth__002 #(.WIDTH(WIDTH)) mul00340009(.x(x_9), .z(tmp00_9_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340010(.x(x_10), .z(tmp00_10_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340011(.x(x_11), .z(tmp00_11_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340012(.x(x_12), .z(tmp00_12_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340013(.x(x_13), .z(tmp00_13_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340014(.x(x_14), .z(tmp00_14_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340015(.x(x_15), .z(tmp00_15_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340016(.x(x_16), .z(tmp00_16_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340017(.x(x_17), .z(tmp00_17_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340018(.x(x_18), .z(tmp00_18_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340019(.x(x_19), .z(tmp00_19_34));
	booth_0002 #(.WIDTH(WIDTH)) mul00340020(.x(x_20), .z(tmp00_20_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340021(.x(x_21), .z(tmp00_21_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340022(.x(x_22), .z(tmp00_22_34));
	booth_0002 #(.WIDTH(WIDTH)) mul00340023(.x(x_23), .z(tmp00_23_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340024(.x(x_24), .z(tmp00_24_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340025(.x(x_25), .z(tmp00_25_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340026(.x(x_26), .z(tmp00_26_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340027(.x(x_27), .z(tmp00_27_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340028(.x(x_28), .z(tmp00_28_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340029(.x(x_29), .z(tmp00_29_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340030(.x(x_30), .z(tmp00_30_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340031(.x(x_31), .z(tmp00_31_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340032(.x(x_32), .z(tmp00_32_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340033(.x(x_33), .z(tmp00_33_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340034(.x(x_34), .z(tmp00_34_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340035(.x(x_35), .z(tmp00_35_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340036(.x(x_36), .z(tmp00_36_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340037(.x(x_37), .z(tmp00_37_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340038(.x(x_38), .z(tmp00_38_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340039(.x(x_39), .z(tmp00_39_34));
	booth__012 #(.WIDTH(WIDTH)) mul00340040(.x(x_40), .z(tmp00_40_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340041(.x(x_41), .z(tmp00_41_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340042(.x(x_42), .z(tmp00_42_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340043(.x(x_43), .z(tmp00_43_34));
	booth__012 #(.WIDTH(WIDTH)) mul00340044(.x(x_44), .z(tmp00_44_34));
	booth_0002 #(.WIDTH(WIDTH)) mul00340045(.x(x_45), .z(tmp00_45_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340046(.x(x_46), .z(tmp00_46_34));
	booth__014 #(.WIDTH(WIDTH)) mul00340047(.x(x_47), .z(tmp00_47_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340048(.x(x_48), .z(tmp00_48_34));
	booth__012 #(.WIDTH(WIDTH)) mul00340049(.x(x_49), .z(tmp00_49_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340050(.x(x_50), .z(tmp00_50_34));
	booth_0006 #(.WIDTH(WIDTH)) mul00340051(.x(x_51), .z(tmp00_51_34));
	booth_0012 #(.WIDTH(WIDTH)) mul00340052(.x(x_52), .z(tmp00_52_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340053(.x(x_53), .z(tmp00_53_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340054(.x(x_54), .z(tmp00_54_34));
	booth_0014 #(.WIDTH(WIDTH)) mul00340055(.x(x_55), .z(tmp00_55_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340056(.x(x_56), .z(tmp00_56_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340057(.x(x_57), .z(tmp00_57_34));
	booth__002 #(.WIDTH(WIDTH)) mul00340058(.x(x_58), .z(tmp00_58_34));
	booth_0018 #(.WIDTH(WIDTH)) mul00340059(.x(x_59), .z(tmp00_59_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340060(.x(x_60), .z(tmp00_60_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340061(.x(x_61), .z(tmp00_61_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340062(.x(x_62), .z(tmp00_62_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340063(.x(x_63), .z(tmp00_63_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340064(.x(x_64), .z(tmp00_64_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340065(.x(x_65), .z(tmp00_65_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340066(.x(x_66), .z(tmp00_66_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340067(.x(x_67), .z(tmp00_67_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340068(.x(x_68), .z(tmp00_68_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340069(.x(x_69), .z(tmp00_69_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340070(.x(x_70), .z(tmp00_70_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340071(.x(x_71), .z(tmp00_71_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340072(.x(x_72), .z(tmp00_72_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340073(.x(x_73), .z(tmp00_73_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340074(.x(x_74), .z(tmp00_74_34));
	booth_0014 #(.WIDTH(WIDTH)) mul00340075(.x(x_75), .z(tmp00_75_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340076(.x(x_76), .z(tmp00_76_34));
	booth__010 #(.WIDTH(WIDTH)) mul00340077(.x(x_77), .z(tmp00_77_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340078(.x(x_78), .z(tmp00_78_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340079(.x(x_79), .z(tmp00_79_34));
	booth__016 #(.WIDTH(WIDTH)) mul00340080(.x(x_80), .z(tmp00_80_34));
	booth_0012 #(.WIDTH(WIDTH)) mul00340081(.x(x_81), .z(tmp00_81_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340082(.x(x_82), .z(tmp00_82_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340083(.x(x_83), .z(tmp00_83_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340084(.x(x_84), .z(tmp00_84_34));
	booth_0016 #(.WIDTH(WIDTH)) mul00340085(.x(x_85), .z(tmp00_85_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340086(.x(x_86), .z(tmp00_86_34));
	booth__012 #(.WIDTH(WIDTH)) mul00340087(.x(x_87), .z(tmp00_87_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340088(.x(x_88), .z(tmp00_88_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340089(.x(x_89), .z(tmp00_89_34));
	booth__012 #(.WIDTH(WIDTH)) mul00340090(.x(x_90), .z(tmp00_90_34));
	booth_0012 #(.WIDTH(WIDTH)) mul00340091(.x(x_91), .z(tmp00_91_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340092(.x(x_92), .z(tmp00_92_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340093(.x(x_93), .z(tmp00_93_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340094(.x(x_94), .z(tmp00_94_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340095(.x(x_95), .z(tmp00_95_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340096(.x(x_96), .z(tmp00_96_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340097(.x(x_97), .z(tmp00_97_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340098(.x(x_98), .z(tmp00_98_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340099(.x(x_99), .z(tmp00_99_34));
	booth__016 #(.WIDTH(WIDTH)) mul00340100(.x(x_100), .z(tmp00_100_34));
	booth__002 #(.WIDTH(WIDTH)) mul00340101(.x(x_101), .z(tmp00_101_34));
	booth__004 #(.WIDTH(WIDTH)) mul00340102(.x(x_102), .z(tmp00_102_34));
	booth__002 #(.WIDTH(WIDTH)) mul00340103(.x(x_103), .z(tmp00_103_34));
	booth__010 #(.WIDTH(WIDTH)) mul00340104(.x(x_104), .z(tmp00_104_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340105(.x(x_105), .z(tmp00_105_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340106(.x(x_106), .z(tmp00_106_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340107(.x(x_107), .z(tmp00_107_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340108(.x(x_108), .z(tmp00_108_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340109(.x(x_109), .z(tmp00_109_34));
	booth_0016 #(.WIDTH(WIDTH)) mul00340110(.x(x_110), .z(tmp00_110_34));
	booth__002 #(.WIDTH(WIDTH)) mul00340111(.x(x_111), .z(tmp00_111_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340112(.x(x_112), .z(tmp00_112_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340113(.x(x_113), .z(tmp00_113_34));
	booth__008 #(.WIDTH(WIDTH)) mul00340114(.x(x_114), .z(tmp00_114_34));
	booth_0016 #(.WIDTH(WIDTH)) mul00340115(.x(x_115), .z(tmp00_115_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340116(.x(x_116), .z(tmp00_116_34));
	booth_0010 #(.WIDTH(WIDTH)) mul00340117(.x(x_117), .z(tmp00_117_34));
	booth_0002 #(.WIDTH(WIDTH)) mul00340118(.x(x_118), .z(tmp00_118_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340119(.x(x_119), .z(tmp00_119_34));
	booth_0016 #(.WIDTH(WIDTH)) mul00340120(.x(x_120), .z(tmp00_120_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340121(.x(x_121), .z(tmp00_121_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340122(.x(x_122), .z(tmp00_122_34));
	booth_0004 #(.WIDTH(WIDTH)) mul00340123(.x(x_123), .z(tmp00_123_34));
	booth_0000 #(.WIDTH(WIDTH)) mul00340124(.x(x_124), .z(tmp00_124_34));
	booth_0002 #(.WIDTH(WIDTH)) mul00340125(.x(x_125), .z(tmp00_125_34));
	booth_0012 #(.WIDTH(WIDTH)) mul00340126(.x(x_126), .z(tmp00_126_34));
	booth_0008 #(.WIDTH(WIDTH)) mul00340127(.x(x_127), .z(tmp00_127_34));
	booth__006 #(.WIDTH(WIDTH)) mul00350000(.x(x_0), .z(tmp00_0_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350001(.x(x_1), .z(tmp00_1_35));
	booth_0010 #(.WIDTH(WIDTH)) mul00350002(.x(x_2), .z(tmp00_2_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350003(.x(x_3), .z(tmp00_3_35));
	booth__020 #(.WIDTH(WIDTH)) mul00350004(.x(x_4), .z(tmp00_4_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350005(.x(x_5), .z(tmp00_5_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350006(.x(x_6), .z(tmp00_6_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350007(.x(x_7), .z(tmp00_7_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350008(.x(x_8), .z(tmp00_8_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350009(.x(x_9), .z(tmp00_9_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350010(.x(x_10), .z(tmp00_10_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350011(.x(x_11), .z(tmp00_11_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350012(.x(x_12), .z(tmp00_12_35));
	booth__002 #(.WIDTH(WIDTH)) mul00350013(.x(x_13), .z(tmp00_13_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350014(.x(x_14), .z(tmp00_14_35));
	booth__002 #(.WIDTH(WIDTH)) mul00350015(.x(x_15), .z(tmp00_15_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350016(.x(x_16), .z(tmp00_16_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350017(.x(x_17), .z(tmp00_17_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350018(.x(x_18), .z(tmp00_18_35));
	booth_0002 #(.WIDTH(WIDTH)) mul00350019(.x(x_19), .z(tmp00_19_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350020(.x(x_20), .z(tmp00_20_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350021(.x(x_21), .z(tmp00_21_35));
	booth_0018 #(.WIDTH(WIDTH)) mul00350022(.x(x_22), .z(tmp00_22_35));
	booth__006 #(.WIDTH(WIDTH)) mul00350023(.x(x_23), .z(tmp00_23_35));
	booth_0014 #(.WIDTH(WIDTH)) mul00350024(.x(x_24), .z(tmp00_24_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350025(.x(x_25), .z(tmp00_25_35));
	booth__012 #(.WIDTH(WIDTH)) mul00350026(.x(x_26), .z(tmp00_26_35));
	booth_0002 #(.WIDTH(WIDTH)) mul00350027(.x(x_27), .z(tmp00_27_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350028(.x(x_28), .z(tmp00_28_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350029(.x(x_29), .z(tmp00_29_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350030(.x(x_30), .z(tmp00_30_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350031(.x(x_31), .z(tmp00_31_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350032(.x(x_32), .z(tmp00_32_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350033(.x(x_33), .z(tmp00_33_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350034(.x(x_34), .z(tmp00_34_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350035(.x(x_35), .z(tmp00_35_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350036(.x(x_36), .z(tmp00_36_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350037(.x(x_37), .z(tmp00_37_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350038(.x(x_38), .z(tmp00_38_35));
	booth_0002 #(.WIDTH(WIDTH)) mul00350039(.x(x_39), .z(tmp00_39_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350040(.x(x_40), .z(tmp00_40_35));
	booth_0014 #(.WIDTH(WIDTH)) mul00350041(.x(x_41), .z(tmp00_41_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350042(.x(x_42), .z(tmp00_42_35));
	booth_0012 #(.WIDTH(WIDTH)) mul00350043(.x(x_43), .z(tmp00_43_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350044(.x(x_44), .z(tmp00_44_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350045(.x(x_45), .z(tmp00_45_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350046(.x(x_46), .z(tmp00_46_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350047(.x(x_47), .z(tmp00_47_35));
	booth__002 #(.WIDTH(WIDTH)) mul00350048(.x(x_48), .z(tmp00_48_35));
	booth_0006 #(.WIDTH(WIDTH)) mul00350049(.x(x_49), .z(tmp00_49_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350050(.x(x_50), .z(tmp00_50_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350051(.x(x_51), .z(tmp00_51_35));
	booth_0018 #(.WIDTH(WIDTH)) mul00350052(.x(x_52), .z(tmp00_52_35));
	booth__010 #(.WIDTH(WIDTH)) mul00350053(.x(x_53), .z(tmp00_53_35));
	booth_0006 #(.WIDTH(WIDTH)) mul00350054(.x(x_54), .z(tmp00_54_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350055(.x(x_55), .z(tmp00_55_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350056(.x(x_56), .z(tmp00_56_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350057(.x(x_57), .z(tmp00_57_35));
	booth_0002 #(.WIDTH(WIDTH)) mul00350058(.x(x_58), .z(tmp00_58_35));
	booth_0028 #(.WIDTH(WIDTH)) mul00350059(.x(x_59), .z(tmp00_59_35));
	booth__006 #(.WIDTH(WIDTH)) mul00350060(.x(x_60), .z(tmp00_60_35));
	booth__006 #(.WIDTH(WIDTH)) mul00350061(.x(x_61), .z(tmp00_61_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350062(.x(x_62), .z(tmp00_62_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350063(.x(x_63), .z(tmp00_63_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350064(.x(x_64), .z(tmp00_64_35));
	booth_0002 #(.WIDTH(WIDTH)) mul00350065(.x(x_65), .z(tmp00_65_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350066(.x(x_66), .z(tmp00_66_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350067(.x(x_67), .z(tmp00_67_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350068(.x(x_68), .z(tmp00_68_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350069(.x(x_69), .z(tmp00_69_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350070(.x(x_70), .z(tmp00_70_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350071(.x(x_71), .z(tmp00_71_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350072(.x(x_72), .z(tmp00_72_35));
	booth__002 #(.WIDTH(WIDTH)) mul00350073(.x(x_73), .z(tmp00_73_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350074(.x(x_74), .z(tmp00_74_35));
	booth_0006 #(.WIDTH(WIDTH)) mul00350075(.x(x_75), .z(tmp00_75_35));
	booth__002 #(.WIDTH(WIDTH)) mul00350076(.x(x_76), .z(tmp00_76_35));
	booth_0012 #(.WIDTH(WIDTH)) mul00350077(.x(x_77), .z(tmp00_77_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350078(.x(x_78), .z(tmp00_78_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350079(.x(x_79), .z(tmp00_79_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350080(.x(x_80), .z(tmp00_80_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350081(.x(x_81), .z(tmp00_81_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350082(.x(x_82), .z(tmp00_82_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350083(.x(x_83), .z(tmp00_83_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350084(.x(x_84), .z(tmp00_84_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350085(.x(x_85), .z(tmp00_85_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350086(.x(x_86), .z(tmp00_86_35));
	booth__016 #(.WIDTH(WIDTH)) mul00350087(.x(x_87), .z(tmp00_87_35));
	booth__016 #(.WIDTH(WIDTH)) mul00350088(.x(x_88), .z(tmp00_88_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350089(.x(x_89), .z(tmp00_89_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350090(.x(x_90), .z(tmp00_90_35));
	booth_0016 #(.WIDTH(WIDTH)) mul00350091(.x(x_91), .z(tmp00_91_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350092(.x(x_92), .z(tmp00_92_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350093(.x(x_93), .z(tmp00_93_35));
	booth_0006 #(.WIDTH(WIDTH)) mul00350094(.x(x_94), .z(tmp00_94_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350095(.x(x_95), .z(tmp00_95_35));
	booth__014 #(.WIDTH(WIDTH)) mul00350096(.x(x_96), .z(tmp00_96_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350097(.x(x_97), .z(tmp00_97_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350098(.x(x_98), .z(tmp00_98_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350099(.x(x_99), .z(tmp00_99_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350100(.x(x_100), .z(tmp00_100_35));
	booth__002 #(.WIDTH(WIDTH)) mul00350101(.x(x_101), .z(tmp00_101_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350102(.x(x_102), .z(tmp00_102_35));
	booth_0006 #(.WIDTH(WIDTH)) mul00350103(.x(x_103), .z(tmp00_103_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350104(.x(x_104), .z(tmp00_104_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350105(.x(x_105), .z(tmp00_105_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350106(.x(x_106), .z(tmp00_106_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350107(.x(x_107), .z(tmp00_107_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350108(.x(x_108), .z(tmp00_108_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350109(.x(x_109), .z(tmp00_109_35));
	booth__016 #(.WIDTH(WIDTH)) mul00350110(.x(x_110), .z(tmp00_110_35));
	booth__010 #(.WIDTH(WIDTH)) mul00350111(.x(x_111), .z(tmp00_111_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350112(.x(x_112), .z(tmp00_112_35));
	booth_0020 #(.WIDTH(WIDTH)) mul00350113(.x(x_113), .z(tmp00_113_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350114(.x(x_114), .z(tmp00_114_35));
	booth_0020 #(.WIDTH(WIDTH)) mul00350115(.x(x_115), .z(tmp00_115_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350116(.x(x_116), .z(tmp00_116_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350117(.x(x_117), .z(tmp00_117_35));
	booth_0008 #(.WIDTH(WIDTH)) mul00350118(.x(x_118), .z(tmp00_118_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350119(.x(x_119), .z(tmp00_119_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350120(.x(x_120), .z(tmp00_120_35));
	booth_0012 #(.WIDTH(WIDTH)) mul00350121(.x(x_121), .z(tmp00_121_35));
	booth__008 #(.WIDTH(WIDTH)) mul00350122(.x(x_122), .z(tmp00_122_35));
	booth__004 #(.WIDTH(WIDTH)) mul00350123(.x(x_123), .z(tmp00_123_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350124(.x(x_124), .z(tmp00_124_35));
	booth_0004 #(.WIDTH(WIDTH)) mul00350125(.x(x_125), .z(tmp00_125_35));
	booth_0016 #(.WIDTH(WIDTH)) mul00350126(.x(x_126), .z(tmp00_126_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00350127(.x(x_127), .z(tmp00_127_35));
	booth_0000 #(.WIDTH(WIDTH)) mul00360000(.x(x_0), .z(tmp00_0_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360001(.x(x_1), .z(tmp00_1_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360002(.x(x_2), .z(tmp00_2_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360003(.x(x_3), .z(tmp00_3_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360004(.x(x_4), .z(tmp00_4_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360005(.x(x_5), .z(tmp00_5_36));
	booth_0006 #(.WIDTH(WIDTH)) mul00360006(.x(x_6), .z(tmp00_6_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360007(.x(x_7), .z(tmp00_7_36));
	booth__010 #(.WIDTH(WIDTH)) mul00360008(.x(x_8), .z(tmp00_8_36));
	booth_0002 #(.WIDTH(WIDTH)) mul00360009(.x(x_9), .z(tmp00_9_36));
	booth__012 #(.WIDTH(WIDTH)) mul00360010(.x(x_10), .z(tmp00_10_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360011(.x(x_11), .z(tmp00_11_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360012(.x(x_12), .z(tmp00_12_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360013(.x(x_13), .z(tmp00_13_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360014(.x(x_14), .z(tmp00_14_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360015(.x(x_15), .z(tmp00_15_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360016(.x(x_16), .z(tmp00_16_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360017(.x(x_17), .z(tmp00_17_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360018(.x(x_18), .z(tmp00_18_36));
	booth_0002 #(.WIDTH(WIDTH)) mul00360019(.x(x_19), .z(tmp00_19_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360020(.x(x_20), .z(tmp00_20_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360021(.x(x_21), .z(tmp00_21_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360022(.x(x_22), .z(tmp00_22_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360023(.x(x_23), .z(tmp00_23_36));
	booth_0012 #(.WIDTH(WIDTH)) mul00360024(.x(x_24), .z(tmp00_24_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360025(.x(x_25), .z(tmp00_25_36));
	booth_0012 #(.WIDTH(WIDTH)) mul00360026(.x(x_26), .z(tmp00_26_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360027(.x(x_27), .z(tmp00_27_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360028(.x(x_28), .z(tmp00_28_36));
	booth_0010 #(.WIDTH(WIDTH)) mul00360029(.x(x_29), .z(tmp00_29_36));
	booth__012 #(.WIDTH(WIDTH)) mul00360030(.x(x_30), .z(tmp00_30_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360031(.x(x_31), .z(tmp00_31_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360032(.x(x_32), .z(tmp00_32_36));
	booth_0006 #(.WIDTH(WIDTH)) mul00360033(.x(x_33), .z(tmp00_33_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360034(.x(x_34), .z(tmp00_34_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360035(.x(x_35), .z(tmp00_35_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360036(.x(x_36), .z(tmp00_36_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360037(.x(x_37), .z(tmp00_37_36));
	booth_0010 #(.WIDTH(WIDTH)) mul00360038(.x(x_38), .z(tmp00_38_36));
	booth__012 #(.WIDTH(WIDTH)) mul00360039(.x(x_39), .z(tmp00_39_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360040(.x(x_40), .z(tmp00_40_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360041(.x(x_41), .z(tmp00_41_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360042(.x(x_42), .z(tmp00_42_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360043(.x(x_43), .z(tmp00_43_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360044(.x(x_44), .z(tmp00_44_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360045(.x(x_45), .z(tmp00_45_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360046(.x(x_46), .z(tmp00_46_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360047(.x(x_47), .z(tmp00_47_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360048(.x(x_48), .z(tmp00_48_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360049(.x(x_49), .z(tmp00_49_36));
	booth__006 #(.WIDTH(WIDTH)) mul00360050(.x(x_50), .z(tmp00_50_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360051(.x(x_51), .z(tmp00_51_36));
	booth_0012 #(.WIDTH(WIDTH)) mul00360052(.x(x_52), .z(tmp00_52_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360053(.x(x_53), .z(tmp00_53_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360054(.x(x_54), .z(tmp00_54_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360055(.x(x_55), .z(tmp00_55_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360056(.x(x_56), .z(tmp00_56_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360057(.x(x_57), .z(tmp00_57_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360058(.x(x_58), .z(tmp00_58_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360059(.x(x_59), .z(tmp00_59_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360060(.x(x_60), .z(tmp00_60_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360061(.x(x_61), .z(tmp00_61_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360062(.x(x_62), .z(tmp00_62_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360063(.x(x_63), .z(tmp00_63_36));
	booth__002 #(.WIDTH(WIDTH)) mul00360064(.x(x_64), .z(tmp00_64_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360065(.x(x_65), .z(tmp00_65_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360066(.x(x_66), .z(tmp00_66_36));
	booth__006 #(.WIDTH(WIDTH)) mul00360067(.x(x_67), .z(tmp00_67_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360068(.x(x_68), .z(tmp00_68_36));
	booth_0002 #(.WIDTH(WIDTH)) mul00360069(.x(x_69), .z(tmp00_69_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360070(.x(x_70), .z(tmp00_70_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360071(.x(x_71), .z(tmp00_71_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360072(.x(x_72), .z(tmp00_72_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360073(.x(x_73), .z(tmp00_73_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360074(.x(x_74), .z(tmp00_74_36));
	booth__002 #(.WIDTH(WIDTH)) mul00360075(.x(x_75), .z(tmp00_75_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360076(.x(x_76), .z(tmp00_76_36));
	booth_0006 #(.WIDTH(WIDTH)) mul00360077(.x(x_77), .z(tmp00_77_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360078(.x(x_78), .z(tmp00_78_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360079(.x(x_79), .z(tmp00_79_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360080(.x(x_80), .z(tmp00_80_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360081(.x(x_81), .z(tmp00_81_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360082(.x(x_82), .z(tmp00_82_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360083(.x(x_83), .z(tmp00_83_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360084(.x(x_84), .z(tmp00_84_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360085(.x(x_85), .z(tmp00_85_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360086(.x(x_86), .z(tmp00_86_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360087(.x(x_87), .z(tmp00_87_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360088(.x(x_88), .z(tmp00_88_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360089(.x(x_89), .z(tmp00_89_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360090(.x(x_90), .z(tmp00_90_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360091(.x(x_91), .z(tmp00_91_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360092(.x(x_92), .z(tmp00_92_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360093(.x(x_93), .z(tmp00_93_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360094(.x(x_94), .z(tmp00_94_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360095(.x(x_95), .z(tmp00_95_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360096(.x(x_96), .z(tmp00_96_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360097(.x(x_97), .z(tmp00_97_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360098(.x(x_98), .z(tmp00_98_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360099(.x(x_99), .z(tmp00_99_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360100(.x(x_100), .z(tmp00_100_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360101(.x(x_101), .z(tmp00_101_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360102(.x(x_102), .z(tmp00_102_36));
	booth__008 #(.WIDTH(WIDTH)) mul00360103(.x(x_103), .z(tmp00_103_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360104(.x(x_104), .z(tmp00_104_36));
	booth__006 #(.WIDTH(WIDTH)) mul00360105(.x(x_105), .z(tmp00_105_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360106(.x(x_106), .z(tmp00_106_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360107(.x(x_107), .z(tmp00_107_36));
	booth__010 #(.WIDTH(WIDTH)) mul00360108(.x(x_108), .z(tmp00_108_36));
	booth_0006 #(.WIDTH(WIDTH)) mul00360109(.x(x_109), .z(tmp00_109_36));
	booth_0010 #(.WIDTH(WIDTH)) mul00360110(.x(x_110), .z(tmp00_110_36));
	booth_0004 #(.WIDTH(WIDTH)) mul00360111(.x(x_111), .z(tmp00_111_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360112(.x(x_112), .z(tmp00_112_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360113(.x(x_113), .z(tmp00_113_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360114(.x(x_114), .z(tmp00_114_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360115(.x(x_115), .z(tmp00_115_36));
	booth_0010 #(.WIDTH(WIDTH)) mul00360116(.x(x_116), .z(tmp00_116_36));
	booth__002 #(.WIDTH(WIDTH)) mul00360117(.x(x_117), .z(tmp00_117_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360118(.x(x_118), .z(tmp00_118_36));
	booth_0006 #(.WIDTH(WIDTH)) mul00360119(.x(x_119), .z(tmp00_119_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360120(.x(x_120), .z(tmp00_120_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360121(.x(x_121), .z(tmp00_121_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360122(.x(x_122), .z(tmp00_122_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360123(.x(x_123), .z(tmp00_123_36));
	booth_0008 #(.WIDTH(WIDTH)) mul00360124(.x(x_124), .z(tmp00_124_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360125(.x(x_125), .z(tmp00_125_36));
	booth__004 #(.WIDTH(WIDTH)) mul00360126(.x(x_126), .z(tmp00_126_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00360127(.x(x_127), .z(tmp00_127_36));
	booth_0000 #(.WIDTH(WIDTH)) mul00370000(.x(x_0), .z(tmp00_0_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370001(.x(x_1), .z(tmp00_1_37));
	booth__010 #(.WIDTH(WIDTH)) mul00370002(.x(x_2), .z(tmp00_2_37));
	booth_0010 #(.WIDTH(WIDTH)) mul00370003(.x(x_3), .z(tmp00_3_37));
	booth_0012 #(.WIDTH(WIDTH)) mul00370004(.x(x_4), .z(tmp00_4_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370005(.x(x_5), .z(tmp00_5_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370006(.x(x_6), .z(tmp00_6_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370007(.x(x_7), .z(tmp00_7_37));
	booth_0010 #(.WIDTH(WIDTH)) mul00370008(.x(x_8), .z(tmp00_8_37));
	booth_0010 #(.WIDTH(WIDTH)) mul00370009(.x(x_9), .z(tmp00_9_37));
	booth__010 #(.WIDTH(WIDTH)) mul00370010(.x(x_10), .z(tmp00_10_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370011(.x(x_11), .z(tmp00_11_37));
	booth_0006 #(.WIDTH(WIDTH)) mul00370012(.x(x_12), .z(tmp00_12_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370013(.x(x_13), .z(tmp00_13_37));
	booth_0004 #(.WIDTH(WIDTH)) mul00370014(.x(x_14), .z(tmp00_14_37));
	booth__010 #(.WIDTH(WIDTH)) mul00370015(.x(x_15), .z(tmp00_15_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370016(.x(x_16), .z(tmp00_16_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370017(.x(x_17), .z(tmp00_17_37));
	booth_0010 #(.WIDTH(WIDTH)) mul00370018(.x(x_18), .z(tmp00_18_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370019(.x(x_19), .z(tmp00_19_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370020(.x(x_20), .z(tmp00_20_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370021(.x(x_21), .z(tmp00_21_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370022(.x(x_22), .z(tmp00_22_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370023(.x(x_23), .z(tmp00_23_37));
	booth_0002 #(.WIDTH(WIDTH)) mul00370024(.x(x_24), .z(tmp00_24_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370025(.x(x_25), .z(tmp00_25_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370026(.x(x_26), .z(tmp00_26_37));
	booth_0002 #(.WIDTH(WIDTH)) mul00370027(.x(x_27), .z(tmp00_27_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370028(.x(x_28), .z(tmp00_28_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370029(.x(x_29), .z(tmp00_29_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370030(.x(x_30), .z(tmp00_30_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370031(.x(x_31), .z(tmp00_31_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370032(.x(x_32), .z(tmp00_32_37));
	booth__012 #(.WIDTH(WIDTH)) mul00370033(.x(x_33), .z(tmp00_33_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370034(.x(x_34), .z(tmp00_34_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370035(.x(x_35), .z(tmp00_35_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370036(.x(x_36), .z(tmp00_36_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370037(.x(x_37), .z(tmp00_37_37));
	booth_0006 #(.WIDTH(WIDTH)) mul00370038(.x(x_38), .z(tmp00_38_37));
	booth_0010 #(.WIDTH(WIDTH)) mul00370039(.x(x_39), .z(tmp00_39_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370040(.x(x_40), .z(tmp00_40_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370041(.x(x_41), .z(tmp00_41_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370042(.x(x_42), .z(tmp00_42_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370043(.x(x_43), .z(tmp00_43_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370044(.x(x_44), .z(tmp00_44_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370045(.x(x_45), .z(tmp00_45_37));
	booth_0014 #(.WIDTH(WIDTH)) mul00370046(.x(x_46), .z(tmp00_46_37));
	booth__014 #(.WIDTH(WIDTH)) mul00370047(.x(x_47), .z(tmp00_47_37));
	booth__006 #(.WIDTH(WIDTH)) mul00370048(.x(x_48), .z(tmp00_48_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370049(.x(x_49), .z(tmp00_49_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370050(.x(x_50), .z(tmp00_50_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370051(.x(x_51), .z(tmp00_51_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370052(.x(x_52), .z(tmp00_52_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370053(.x(x_53), .z(tmp00_53_37));
	booth__010 #(.WIDTH(WIDTH)) mul00370054(.x(x_54), .z(tmp00_54_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370055(.x(x_55), .z(tmp00_55_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370056(.x(x_56), .z(tmp00_56_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370057(.x(x_57), .z(tmp00_57_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370058(.x(x_58), .z(tmp00_58_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370059(.x(x_59), .z(tmp00_59_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370060(.x(x_60), .z(tmp00_60_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370061(.x(x_61), .z(tmp00_61_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370062(.x(x_62), .z(tmp00_62_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370063(.x(x_63), .z(tmp00_63_37));
	booth_0010 #(.WIDTH(WIDTH)) mul00370064(.x(x_64), .z(tmp00_64_37));
	booth_0004 #(.WIDTH(WIDTH)) mul00370065(.x(x_65), .z(tmp00_65_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370066(.x(x_66), .z(tmp00_66_37));
	booth__010 #(.WIDTH(WIDTH)) mul00370067(.x(x_67), .z(tmp00_67_37));
	booth_0012 #(.WIDTH(WIDTH)) mul00370068(.x(x_68), .z(tmp00_68_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370069(.x(x_69), .z(tmp00_69_37));
	booth_0004 #(.WIDTH(WIDTH)) mul00370070(.x(x_70), .z(tmp00_70_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370071(.x(x_71), .z(tmp00_71_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370072(.x(x_72), .z(tmp00_72_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370073(.x(x_73), .z(tmp00_73_37));
	booth_0004 #(.WIDTH(WIDTH)) mul00370074(.x(x_74), .z(tmp00_74_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370075(.x(x_75), .z(tmp00_75_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370076(.x(x_76), .z(tmp00_76_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370077(.x(x_77), .z(tmp00_77_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370078(.x(x_78), .z(tmp00_78_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370079(.x(x_79), .z(tmp00_79_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370080(.x(x_80), .z(tmp00_80_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370081(.x(x_81), .z(tmp00_81_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370082(.x(x_82), .z(tmp00_82_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370083(.x(x_83), .z(tmp00_83_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370084(.x(x_84), .z(tmp00_84_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370085(.x(x_85), .z(tmp00_85_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370086(.x(x_86), .z(tmp00_86_37));
	booth_0002 #(.WIDTH(WIDTH)) mul00370087(.x(x_87), .z(tmp00_87_37));
	booth_0012 #(.WIDTH(WIDTH)) mul00370088(.x(x_88), .z(tmp00_88_37));
	booth__002 #(.WIDTH(WIDTH)) mul00370089(.x(x_89), .z(tmp00_89_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370090(.x(x_90), .z(tmp00_90_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370091(.x(x_91), .z(tmp00_91_37));
	booth_0002 #(.WIDTH(WIDTH)) mul00370092(.x(x_92), .z(tmp00_92_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370093(.x(x_93), .z(tmp00_93_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370094(.x(x_94), .z(tmp00_94_37));
	booth__008 #(.WIDTH(WIDTH)) mul00370095(.x(x_95), .z(tmp00_95_37));
	booth_0010 #(.WIDTH(WIDTH)) mul00370096(.x(x_96), .z(tmp00_96_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370097(.x(x_97), .z(tmp00_97_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370098(.x(x_98), .z(tmp00_98_37));
	booth_0006 #(.WIDTH(WIDTH)) mul00370099(.x(x_99), .z(tmp00_99_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370100(.x(x_100), .z(tmp00_100_37));
	booth__002 #(.WIDTH(WIDTH)) mul00370101(.x(x_101), .z(tmp00_101_37));
	booth_0012 #(.WIDTH(WIDTH)) mul00370102(.x(x_102), .z(tmp00_102_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370103(.x(x_103), .z(tmp00_103_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370104(.x(x_104), .z(tmp00_104_37));
	booth__002 #(.WIDTH(WIDTH)) mul00370105(.x(x_105), .z(tmp00_105_37));
	booth_0010 #(.WIDTH(WIDTH)) mul00370106(.x(x_106), .z(tmp00_106_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370107(.x(x_107), .z(tmp00_107_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370108(.x(x_108), .z(tmp00_108_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370109(.x(x_109), .z(tmp00_109_37));
	booth_0006 #(.WIDTH(WIDTH)) mul00370110(.x(x_110), .z(tmp00_110_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370111(.x(x_111), .z(tmp00_111_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370112(.x(x_112), .z(tmp00_112_37));
	booth__012 #(.WIDTH(WIDTH)) mul00370113(.x(x_113), .z(tmp00_113_37));
	booth__016 #(.WIDTH(WIDTH)) mul00370114(.x(x_114), .z(tmp00_114_37));
	booth__014 #(.WIDTH(WIDTH)) mul00370115(.x(x_115), .z(tmp00_115_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370116(.x(x_116), .z(tmp00_116_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370117(.x(x_117), .z(tmp00_117_37));
	booth_0012 #(.WIDTH(WIDTH)) mul00370118(.x(x_118), .z(tmp00_118_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370119(.x(x_119), .z(tmp00_119_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370120(.x(x_120), .z(tmp00_120_37));
	booth__016 #(.WIDTH(WIDTH)) mul00370121(.x(x_121), .z(tmp00_121_37));
	booth__006 #(.WIDTH(WIDTH)) mul00370122(.x(x_122), .z(tmp00_122_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370123(.x(x_123), .z(tmp00_123_37));
	booth__004 #(.WIDTH(WIDTH)) mul00370124(.x(x_124), .z(tmp00_124_37));
	booth__012 #(.WIDTH(WIDTH)) mul00370125(.x(x_125), .z(tmp00_125_37));
	booth_0008 #(.WIDTH(WIDTH)) mul00370126(.x(x_126), .z(tmp00_126_37));
	booth_0000 #(.WIDTH(WIDTH)) mul00370127(.x(x_127), .z(tmp00_127_37));
	booth__008 #(.WIDTH(WIDTH)) mul00380000(.x(x_0), .z(tmp00_0_38));
	booth__002 #(.WIDTH(WIDTH)) mul00380001(.x(x_1), .z(tmp00_1_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380002(.x(x_2), .z(tmp00_2_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380003(.x(x_3), .z(tmp00_3_38));
	booth__006 #(.WIDTH(WIDTH)) mul00380004(.x(x_4), .z(tmp00_4_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380005(.x(x_5), .z(tmp00_5_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380006(.x(x_6), .z(tmp00_6_38));
	booth__006 #(.WIDTH(WIDTH)) mul00380007(.x(x_7), .z(tmp00_7_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380008(.x(x_8), .z(tmp00_8_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380009(.x(x_9), .z(tmp00_9_38));
	booth_0002 #(.WIDTH(WIDTH)) mul00380010(.x(x_10), .z(tmp00_10_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380011(.x(x_11), .z(tmp00_11_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380012(.x(x_12), .z(tmp00_12_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380013(.x(x_13), .z(tmp00_13_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380014(.x(x_14), .z(tmp00_14_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380015(.x(x_15), .z(tmp00_15_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380016(.x(x_16), .z(tmp00_16_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380017(.x(x_17), .z(tmp00_17_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380018(.x(x_18), .z(tmp00_18_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380019(.x(x_19), .z(tmp00_19_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380020(.x(x_20), .z(tmp00_20_38));
	booth__006 #(.WIDTH(WIDTH)) mul00380021(.x(x_21), .z(tmp00_21_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380022(.x(x_22), .z(tmp00_22_38));
	booth_0010 #(.WIDTH(WIDTH)) mul00380023(.x(x_23), .z(tmp00_23_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380024(.x(x_24), .z(tmp00_24_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380025(.x(x_25), .z(tmp00_25_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380026(.x(x_26), .z(tmp00_26_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380027(.x(x_27), .z(tmp00_27_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380028(.x(x_28), .z(tmp00_28_38));
	booth_0006 #(.WIDTH(WIDTH)) mul00380029(.x(x_29), .z(tmp00_29_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380030(.x(x_30), .z(tmp00_30_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380031(.x(x_31), .z(tmp00_31_38));
	booth__006 #(.WIDTH(WIDTH)) mul00380032(.x(x_32), .z(tmp00_32_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380033(.x(x_33), .z(tmp00_33_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380034(.x(x_34), .z(tmp00_34_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380035(.x(x_35), .z(tmp00_35_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380036(.x(x_36), .z(tmp00_36_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380037(.x(x_37), .z(tmp00_37_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380038(.x(x_38), .z(tmp00_38_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380039(.x(x_39), .z(tmp00_39_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380040(.x(x_40), .z(tmp00_40_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380041(.x(x_41), .z(tmp00_41_38));
	booth_0006 #(.WIDTH(WIDTH)) mul00380042(.x(x_42), .z(tmp00_42_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380043(.x(x_43), .z(tmp00_43_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380044(.x(x_44), .z(tmp00_44_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380045(.x(x_45), .z(tmp00_45_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380046(.x(x_46), .z(tmp00_46_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380047(.x(x_47), .z(tmp00_47_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380048(.x(x_48), .z(tmp00_48_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380049(.x(x_49), .z(tmp00_49_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380050(.x(x_50), .z(tmp00_50_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380051(.x(x_51), .z(tmp00_51_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380052(.x(x_52), .z(tmp00_52_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380053(.x(x_53), .z(tmp00_53_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380054(.x(x_54), .z(tmp00_54_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380055(.x(x_55), .z(tmp00_55_38));
	booth__010 #(.WIDTH(WIDTH)) mul00380056(.x(x_56), .z(tmp00_56_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380057(.x(x_57), .z(tmp00_57_38));
	booth__002 #(.WIDTH(WIDTH)) mul00380058(.x(x_58), .z(tmp00_58_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380059(.x(x_59), .z(tmp00_59_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380060(.x(x_60), .z(tmp00_60_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380061(.x(x_61), .z(tmp00_61_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380062(.x(x_62), .z(tmp00_62_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380063(.x(x_63), .z(tmp00_63_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380064(.x(x_64), .z(tmp00_64_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380065(.x(x_65), .z(tmp00_65_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380066(.x(x_66), .z(tmp00_66_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380067(.x(x_67), .z(tmp00_67_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380068(.x(x_68), .z(tmp00_68_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380069(.x(x_69), .z(tmp00_69_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380070(.x(x_70), .z(tmp00_70_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380071(.x(x_71), .z(tmp00_71_38));
	booth_0006 #(.WIDTH(WIDTH)) mul00380072(.x(x_72), .z(tmp00_72_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380073(.x(x_73), .z(tmp00_73_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380074(.x(x_74), .z(tmp00_74_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380075(.x(x_75), .z(tmp00_75_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380076(.x(x_76), .z(tmp00_76_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380077(.x(x_77), .z(tmp00_77_38));
	booth_0002 #(.WIDTH(WIDTH)) mul00380078(.x(x_78), .z(tmp00_78_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380079(.x(x_79), .z(tmp00_79_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380080(.x(x_80), .z(tmp00_80_38));
	booth__006 #(.WIDTH(WIDTH)) mul00380081(.x(x_81), .z(tmp00_81_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380082(.x(x_82), .z(tmp00_82_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380083(.x(x_83), .z(tmp00_83_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380084(.x(x_84), .z(tmp00_84_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380085(.x(x_85), .z(tmp00_85_38));
	booth__010 #(.WIDTH(WIDTH)) mul00380086(.x(x_86), .z(tmp00_86_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380087(.x(x_87), .z(tmp00_87_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380088(.x(x_88), .z(tmp00_88_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380089(.x(x_89), .z(tmp00_89_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380090(.x(x_90), .z(tmp00_90_38));
	booth__002 #(.WIDTH(WIDTH)) mul00380091(.x(x_91), .z(tmp00_91_38));
	booth_0002 #(.WIDTH(WIDTH)) mul00380092(.x(x_92), .z(tmp00_92_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380093(.x(x_93), .z(tmp00_93_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380094(.x(x_94), .z(tmp00_94_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380095(.x(x_95), .z(tmp00_95_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380096(.x(x_96), .z(tmp00_96_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380097(.x(x_97), .z(tmp00_97_38));
	booth_0006 #(.WIDTH(WIDTH)) mul00380098(.x(x_98), .z(tmp00_98_38));
	booth_0010 #(.WIDTH(WIDTH)) mul00380099(.x(x_99), .z(tmp00_99_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380100(.x(x_100), .z(tmp00_100_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380101(.x(x_101), .z(tmp00_101_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380102(.x(x_102), .z(tmp00_102_38));
	booth__002 #(.WIDTH(WIDTH)) mul00380103(.x(x_103), .z(tmp00_103_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380104(.x(x_104), .z(tmp00_104_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380105(.x(x_105), .z(tmp00_105_38));
	booth__006 #(.WIDTH(WIDTH)) mul00380106(.x(x_106), .z(tmp00_106_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380107(.x(x_107), .z(tmp00_107_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380108(.x(x_108), .z(tmp00_108_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380109(.x(x_109), .z(tmp00_109_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380110(.x(x_110), .z(tmp00_110_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380111(.x(x_111), .z(tmp00_111_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380112(.x(x_112), .z(tmp00_112_38));
	booth__004 #(.WIDTH(WIDTH)) mul00380113(.x(x_113), .z(tmp00_113_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380114(.x(x_114), .z(tmp00_114_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380115(.x(x_115), .z(tmp00_115_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380116(.x(x_116), .z(tmp00_116_38));
	booth_0006 #(.WIDTH(WIDTH)) mul00380117(.x(x_117), .z(tmp00_117_38));
	booth__010 #(.WIDTH(WIDTH)) mul00380118(.x(x_118), .z(tmp00_118_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380119(.x(x_119), .z(tmp00_119_38));
	booth_0008 #(.WIDTH(WIDTH)) mul00380120(.x(x_120), .z(tmp00_120_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380121(.x(x_121), .z(tmp00_121_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380122(.x(x_122), .z(tmp00_122_38));
	booth_0004 #(.WIDTH(WIDTH)) mul00380123(.x(x_123), .z(tmp00_123_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380124(.x(x_124), .z(tmp00_124_38));
	booth__008 #(.WIDTH(WIDTH)) mul00380125(.x(x_125), .z(tmp00_125_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380126(.x(x_126), .z(tmp00_126_38));
	booth_0000 #(.WIDTH(WIDTH)) mul00380127(.x(x_127), .z(tmp00_127_38));
	booth__004 #(.WIDTH(WIDTH)) mul00390000(.x(x_0), .z(tmp00_0_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390001(.x(x_1), .z(tmp00_1_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390002(.x(x_2), .z(tmp00_2_39));
	booth__010 #(.WIDTH(WIDTH)) mul00390003(.x(x_3), .z(tmp00_3_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390004(.x(x_4), .z(tmp00_4_39));
	booth_0006 #(.WIDTH(WIDTH)) mul00390005(.x(x_5), .z(tmp00_5_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390006(.x(x_6), .z(tmp00_6_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390007(.x(x_7), .z(tmp00_7_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390008(.x(x_8), .z(tmp00_8_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390009(.x(x_9), .z(tmp00_9_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390010(.x(x_10), .z(tmp00_10_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390011(.x(x_11), .z(tmp00_11_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390012(.x(x_12), .z(tmp00_12_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390013(.x(x_13), .z(tmp00_13_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390014(.x(x_14), .z(tmp00_14_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390015(.x(x_15), .z(tmp00_15_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390016(.x(x_16), .z(tmp00_16_39));
	booth__010 #(.WIDTH(WIDTH)) mul00390017(.x(x_17), .z(tmp00_17_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390018(.x(x_18), .z(tmp00_18_39));
	booth__010 #(.WIDTH(WIDTH)) mul00390019(.x(x_19), .z(tmp00_19_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390020(.x(x_20), .z(tmp00_20_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390021(.x(x_21), .z(tmp00_21_39));
	booth_0012 #(.WIDTH(WIDTH)) mul00390022(.x(x_22), .z(tmp00_22_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390023(.x(x_23), .z(tmp00_23_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390024(.x(x_24), .z(tmp00_24_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390025(.x(x_25), .z(tmp00_25_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390026(.x(x_26), .z(tmp00_26_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390027(.x(x_27), .z(tmp00_27_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390028(.x(x_28), .z(tmp00_28_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390029(.x(x_29), .z(tmp00_29_39));
	booth_0006 #(.WIDTH(WIDTH)) mul00390030(.x(x_30), .z(tmp00_30_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390031(.x(x_31), .z(tmp00_31_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390032(.x(x_32), .z(tmp00_32_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390033(.x(x_33), .z(tmp00_33_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390034(.x(x_34), .z(tmp00_34_39));
	booth__012 #(.WIDTH(WIDTH)) mul00390035(.x(x_35), .z(tmp00_35_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390036(.x(x_36), .z(tmp00_36_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390037(.x(x_37), .z(tmp00_37_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390038(.x(x_38), .z(tmp00_38_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390039(.x(x_39), .z(tmp00_39_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390040(.x(x_40), .z(tmp00_40_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390041(.x(x_41), .z(tmp00_41_39));
	booth_0006 #(.WIDTH(WIDTH)) mul00390042(.x(x_42), .z(tmp00_42_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390043(.x(x_43), .z(tmp00_43_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390044(.x(x_44), .z(tmp00_44_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390045(.x(x_45), .z(tmp00_45_39));
	booth_0012 #(.WIDTH(WIDTH)) mul00390046(.x(x_46), .z(tmp00_46_39));
	booth__010 #(.WIDTH(WIDTH)) mul00390047(.x(x_47), .z(tmp00_47_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390048(.x(x_48), .z(tmp00_48_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390049(.x(x_49), .z(tmp00_49_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390050(.x(x_50), .z(tmp00_50_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390051(.x(x_51), .z(tmp00_51_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390052(.x(x_52), .z(tmp00_52_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390053(.x(x_53), .z(tmp00_53_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390054(.x(x_54), .z(tmp00_54_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390055(.x(x_55), .z(tmp00_55_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390056(.x(x_56), .z(tmp00_56_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390057(.x(x_57), .z(tmp00_57_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390058(.x(x_58), .z(tmp00_58_39));
	booth_0006 #(.WIDTH(WIDTH)) mul00390059(.x(x_59), .z(tmp00_59_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390060(.x(x_60), .z(tmp00_60_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390061(.x(x_61), .z(tmp00_61_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390062(.x(x_62), .z(tmp00_62_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390063(.x(x_63), .z(tmp00_63_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390064(.x(x_64), .z(tmp00_64_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390065(.x(x_65), .z(tmp00_65_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390066(.x(x_66), .z(tmp00_66_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390067(.x(x_67), .z(tmp00_67_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390068(.x(x_68), .z(tmp00_68_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390069(.x(x_69), .z(tmp00_69_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390070(.x(x_70), .z(tmp00_70_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390071(.x(x_71), .z(tmp00_71_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390072(.x(x_72), .z(tmp00_72_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390073(.x(x_73), .z(tmp00_73_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390074(.x(x_74), .z(tmp00_74_39));
	booth__010 #(.WIDTH(WIDTH)) mul00390075(.x(x_75), .z(tmp00_75_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390076(.x(x_76), .z(tmp00_76_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390077(.x(x_77), .z(tmp00_77_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390078(.x(x_78), .z(tmp00_78_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390079(.x(x_79), .z(tmp00_79_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390080(.x(x_80), .z(tmp00_80_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390081(.x(x_81), .z(tmp00_81_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390082(.x(x_82), .z(tmp00_82_39));
	booth__010 #(.WIDTH(WIDTH)) mul00390083(.x(x_83), .z(tmp00_83_39));
	booth_0012 #(.WIDTH(WIDTH)) mul00390084(.x(x_84), .z(tmp00_84_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390085(.x(x_85), .z(tmp00_85_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390086(.x(x_86), .z(tmp00_86_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390087(.x(x_87), .z(tmp00_87_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390088(.x(x_88), .z(tmp00_88_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390089(.x(x_89), .z(tmp00_89_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390090(.x(x_90), .z(tmp00_90_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390091(.x(x_91), .z(tmp00_91_39));
	booth_0012 #(.WIDTH(WIDTH)) mul00390092(.x(x_92), .z(tmp00_92_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390093(.x(x_93), .z(tmp00_93_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390094(.x(x_94), .z(tmp00_94_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390095(.x(x_95), .z(tmp00_95_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390096(.x(x_96), .z(tmp00_96_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390097(.x(x_97), .z(tmp00_97_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390098(.x(x_98), .z(tmp00_98_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390099(.x(x_99), .z(tmp00_99_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390100(.x(x_100), .z(tmp00_100_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390101(.x(x_101), .z(tmp00_101_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390102(.x(x_102), .z(tmp00_102_39));
	booth_0006 #(.WIDTH(WIDTH)) mul00390103(.x(x_103), .z(tmp00_103_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390104(.x(x_104), .z(tmp00_104_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390105(.x(x_105), .z(tmp00_105_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390106(.x(x_106), .z(tmp00_106_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390107(.x(x_107), .z(tmp00_107_39));
	booth__006 #(.WIDTH(WIDTH)) mul00390108(.x(x_108), .z(tmp00_108_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390109(.x(x_109), .z(tmp00_109_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390110(.x(x_110), .z(tmp00_110_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390111(.x(x_111), .z(tmp00_111_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390112(.x(x_112), .z(tmp00_112_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390113(.x(x_113), .z(tmp00_113_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390114(.x(x_114), .z(tmp00_114_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390115(.x(x_115), .z(tmp00_115_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390116(.x(x_116), .z(tmp00_116_39));
	booth_0006 #(.WIDTH(WIDTH)) mul00390117(.x(x_117), .z(tmp00_117_39));
	booth_0000 #(.WIDTH(WIDTH)) mul00390118(.x(x_118), .z(tmp00_118_39));
	booth_0004 #(.WIDTH(WIDTH)) mul00390119(.x(x_119), .z(tmp00_119_39));
	booth__002 #(.WIDTH(WIDTH)) mul00390120(.x(x_120), .z(tmp00_120_39));
	booth_0002 #(.WIDTH(WIDTH)) mul00390121(.x(x_121), .z(tmp00_121_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390122(.x(x_122), .z(tmp00_122_39));
	booth__004 #(.WIDTH(WIDTH)) mul00390123(.x(x_123), .z(tmp00_123_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390124(.x(x_124), .z(tmp00_124_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390125(.x(x_125), .z(tmp00_125_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00390126(.x(x_126), .z(tmp00_126_39));
	booth__008 #(.WIDTH(WIDTH)) mul00390127(.x(x_127), .z(tmp00_127_39));
	booth_0008 #(.WIDTH(WIDTH)) mul00400000(.x(x_0), .z(tmp00_0_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400001(.x(x_1), .z(tmp00_1_40));
	booth_0010 #(.WIDTH(WIDTH)) mul00400002(.x(x_2), .z(tmp00_2_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400003(.x(x_3), .z(tmp00_3_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400004(.x(x_4), .z(tmp00_4_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400005(.x(x_5), .z(tmp00_5_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400006(.x(x_6), .z(tmp00_6_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400007(.x(x_7), .z(tmp00_7_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400008(.x(x_8), .z(tmp00_8_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400009(.x(x_9), .z(tmp00_9_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400010(.x(x_10), .z(tmp00_10_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400011(.x(x_11), .z(tmp00_11_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400012(.x(x_12), .z(tmp00_12_40));
	booth_0010 #(.WIDTH(WIDTH)) mul00400013(.x(x_13), .z(tmp00_13_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400014(.x(x_14), .z(tmp00_14_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400015(.x(x_15), .z(tmp00_15_40));
	booth_0002 #(.WIDTH(WIDTH)) mul00400016(.x(x_16), .z(tmp00_16_40));
	booth__006 #(.WIDTH(WIDTH)) mul00400017(.x(x_17), .z(tmp00_17_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400018(.x(x_18), .z(tmp00_18_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400019(.x(x_19), .z(tmp00_19_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400020(.x(x_20), .z(tmp00_20_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400021(.x(x_21), .z(tmp00_21_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400022(.x(x_22), .z(tmp00_22_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400023(.x(x_23), .z(tmp00_23_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400024(.x(x_24), .z(tmp00_24_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400025(.x(x_25), .z(tmp00_25_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400026(.x(x_26), .z(tmp00_26_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400027(.x(x_27), .z(tmp00_27_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400028(.x(x_28), .z(tmp00_28_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400029(.x(x_29), .z(tmp00_29_40));
	booth_0006 #(.WIDTH(WIDTH)) mul00400030(.x(x_30), .z(tmp00_30_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400031(.x(x_31), .z(tmp00_31_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400032(.x(x_32), .z(tmp00_32_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400033(.x(x_33), .z(tmp00_33_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400034(.x(x_34), .z(tmp00_34_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400035(.x(x_35), .z(tmp00_35_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400036(.x(x_36), .z(tmp00_36_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400037(.x(x_37), .z(tmp00_37_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400038(.x(x_38), .z(tmp00_38_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400039(.x(x_39), .z(tmp00_39_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400040(.x(x_40), .z(tmp00_40_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400041(.x(x_41), .z(tmp00_41_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400042(.x(x_42), .z(tmp00_42_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400043(.x(x_43), .z(tmp00_43_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400044(.x(x_44), .z(tmp00_44_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400045(.x(x_45), .z(tmp00_45_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400046(.x(x_46), .z(tmp00_46_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400047(.x(x_47), .z(tmp00_47_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400048(.x(x_48), .z(tmp00_48_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400049(.x(x_49), .z(tmp00_49_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400050(.x(x_50), .z(tmp00_50_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400051(.x(x_51), .z(tmp00_51_40));
	booth_0010 #(.WIDTH(WIDTH)) mul00400052(.x(x_52), .z(tmp00_52_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400053(.x(x_53), .z(tmp00_53_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400054(.x(x_54), .z(tmp00_54_40));
	booth_0006 #(.WIDTH(WIDTH)) mul00400055(.x(x_55), .z(tmp00_55_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400056(.x(x_56), .z(tmp00_56_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400057(.x(x_57), .z(tmp00_57_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400058(.x(x_58), .z(tmp00_58_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400059(.x(x_59), .z(tmp00_59_40));
	booth__006 #(.WIDTH(WIDTH)) mul00400060(.x(x_60), .z(tmp00_60_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400061(.x(x_61), .z(tmp00_61_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400062(.x(x_62), .z(tmp00_62_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400063(.x(x_63), .z(tmp00_63_40));
	booth_0006 #(.WIDTH(WIDTH)) mul00400064(.x(x_64), .z(tmp00_64_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400065(.x(x_65), .z(tmp00_65_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400066(.x(x_66), .z(tmp00_66_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400067(.x(x_67), .z(tmp00_67_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400068(.x(x_68), .z(tmp00_68_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400069(.x(x_69), .z(tmp00_69_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400070(.x(x_70), .z(tmp00_70_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400071(.x(x_71), .z(tmp00_71_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400072(.x(x_72), .z(tmp00_72_40));
	booth_0006 #(.WIDTH(WIDTH)) mul00400073(.x(x_73), .z(tmp00_73_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400074(.x(x_74), .z(tmp00_74_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400075(.x(x_75), .z(tmp00_75_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400076(.x(x_76), .z(tmp00_76_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400077(.x(x_77), .z(tmp00_77_40));
	booth_0010 #(.WIDTH(WIDTH)) mul00400078(.x(x_78), .z(tmp00_78_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400079(.x(x_79), .z(tmp00_79_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400080(.x(x_80), .z(tmp00_80_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400081(.x(x_81), .z(tmp00_81_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400082(.x(x_82), .z(tmp00_82_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400083(.x(x_83), .z(tmp00_83_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400084(.x(x_84), .z(tmp00_84_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400085(.x(x_85), .z(tmp00_85_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400086(.x(x_86), .z(tmp00_86_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400087(.x(x_87), .z(tmp00_87_40));
	booth_0008 #(.WIDTH(WIDTH)) mul00400088(.x(x_88), .z(tmp00_88_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400089(.x(x_89), .z(tmp00_89_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400090(.x(x_90), .z(tmp00_90_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400091(.x(x_91), .z(tmp00_91_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400092(.x(x_92), .z(tmp00_92_40));
	booth_0012 #(.WIDTH(WIDTH)) mul00400093(.x(x_93), .z(tmp00_93_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400094(.x(x_94), .z(tmp00_94_40));
	booth_0002 #(.WIDTH(WIDTH)) mul00400095(.x(x_95), .z(tmp00_95_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400096(.x(x_96), .z(tmp00_96_40));
	booth_0006 #(.WIDTH(WIDTH)) mul00400097(.x(x_97), .z(tmp00_97_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400098(.x(x_98), .z(tmp00_98_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400099(.x(x_99), .z(tmp00_99_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400100(.x(x_100), .z(tmp00_100_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400101(.x(x_101), .z(tmp00_101_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400102(.x(x_102), .z(tmp00_102_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400103(.x(x_103), .z(tmp00_103_40));
	booth_0006 #(.WIDTH(WIDTH)) mul00400104(.x(x_104), .z(tmp00_104_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400105(.x(x_105), .z(tmp00_105_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400106(.x(x_106), .z(tmp00_106_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400107(.x(x_107), .z(tmp00_107_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400108(.x(x_108), .z(tmp00_108_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400109(.x(x_109), .z(tmp00_109_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400110(.x(x_110), .z(tmp00_110_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400111(.x(x_111), .z(tmp00_111_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400112(.x(x_112), .z(tmp00_112_40));
	booth_0012 #(.WIDTH(WIDTH)) mul00400113(.x(x_113), .z(tmp00_113_40));
	booth__006 #(.WIDTH(WIDTH)) mul00400114(.x(x_114), .z(tmp00_114_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400115(.x(x_115), .z(tmp00_115_40));
	booth__012 #(.WIDTH(WIDTH)) mul00400116(.x(x_116), .z(tmp00_116_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400117(.x(x_117), .z(tmp00_117_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400118(.x(x_118), .z(tmp00_118_40));
	booth_0010 #(.WIDTH(WIDTH)) mul00400119(.x(x_119), .z(tmp00_119_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400120(.x(x_120), .z(tmp00_120_40));
	booth_0000 #(.WIDTH(WIDTH)) mul00400121(.x(x_121), .z(tmp00_121_40));
	booth__004 #(.WIDTH(WIDTH)) mul00400122(.x(x_122), .z(tmp00_122_40));
	booth__010 #(.WIDTH(WIDTH)) mul00400123(.x(x_123), .z(tmp00_123_40));
	booth_0004 #(.WIDTH(WIDTH)) mul00400124(.x(x_124), .z(tmp00_124_40));
	booth_0010 #(.WIDTH(WIDTH)) mul00400125(.x(x_125), .z(tmp00_125_40));
	booth__002 #(.WIDTH(WIDTH)) mul00400126(.x(x_126), .z(tmp00_126_40));
	booth__008 #(.WIDTH(WIDTH)) mul00400127(.x(x_127), .z(tmp00_127_40));
	booth__008 #(.WIDTH(WIDTH)) mul00410000(.x(x_0), .z(tmp00_0_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410001(.x(x_1), .z(tmp00_1_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410002(.x(x_2), .z(tmp00_2_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410003(.x(x_3), .z(tmp00_3_41));
	booth_0016 #(.WIDTH(WIDTH)) mul00410004(.x(x_4), .z(tmp00_4_41));
	booth_0006 #(.WIDTH(WIDTH)) mul00410005(.x(x_5), .z(tmp00_5_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410006(.x(x_6), .z(tmp00_6_41));
	booth_0012 #(.WIDTH(WIDTH)) mul00410007(.x(x_7), .z(tmp00_7_41));
	booth__006 #(.WIDTH(WIDTH)) mul00410008(.x(x_8), .z(tmp00_8_41));
	booth__006 #(.WIDTH(WIDTH)) mul00410009(.x(x_9), .z(tmp00_9_41));
	booth__010 #(.WIDTH(WIDTH)) mul00410010(.x(x_10), .z(tmp00_10_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410011(.x(x_11), .z(tmp00_11_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410012(.x(x_12), .z(tmp00_12_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410013(.x(x_13), .z(tmp00_13_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410014(.x(x_14), .z(tmp00_14_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410015(.x(x_15), .z(tmp00_15_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410016(.x(x_16), .z(tmp00_16_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410017(.x(x_17), .z(tmp00_17_41));
	booth__006 #(.WIDTH(WIDTH)) mul00410018(.x(x_18), .z(tmp00_18_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410019(.x(x_19), .z(tmp00_19_41));
	booth_0006 #(.WIDTH(WIDTH)) mul00410020(.x(x_20), .z(tmp00_20_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410021(.x(x_21), .z(tmp00_21_41));
	booth__016 #(.WIDTH(WIDTH)) mul00410022(.x(x_22), .z(tmp00_22_41));
	booth_0012 #(.WIDTH(WIDTH)) mul00410023(.x(x_23), .z(tmp00_23_41));
	booth__002 #(.WIDTH(WIDTH)) mul00410024(.x(x_24), .z(tmp00_24_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410025(.x(x_25), .z(tmp00_25_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410026(.x(x_26), .z(tmp00_26_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410027(.x(x_27), .z(tmp00_27_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410028(.x(x_28), .z(tmp00_28_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410029(.x(x_29), .z(tmp00_29_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410030(.x(x_30), .z(tmp00_30_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410031(.x(x_31), .z(tmp00_31_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410032(.x(x_32), .z(tmp00_32_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410033(.x(x_33), .z(tmp00_33_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410034(.x(x_34), .z(tmp00_34_41));
	booth__006 #(.WIDTH(WIDTH)) mul00410035(.x(x_35), .z(tmp00_35_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410036(.x(x_36), .z(tmp00_36_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410037(.x(x_37), .z(tmp00_37_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410038(.x(x_38), .z(tmp00_38_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410039(.x(x_39), .z(tmp00_39_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410040(.x(x_40), .z(tmp00_40_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410041(.x(x_41), .z(tmp00_41_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410042(.x(x_42), .z(tmp00_42_41));
	booth_0016 #(.WIDTH(WIDTH)) mul00410043(.x(x_43), .z(tmp00_43_41));
	booth__016 #(.WIDTH(WIDTH)) mul00410044(.x(x_44), .z(tmp00_44_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410045(.x(x_45), .z(tmp00_45_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410046(.x(x_46), .z(tmp00_46_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410047(.x(x_47), .z(tmp00_47_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410048(.x(x_48), .z(tmp00_48_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410049(.x(x_49), .z(tmp00_49_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410050(.x(x_50), .z(tmp00_50_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410051(.x(x_51), .z(tmp00_51_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410052(.x(x_52), .z(tmp00_52_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410053(.x(x_53), .z(tmp00_53_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410054(.x(x_54), .z(tmp00_54_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410055(.x(x_55), .z(tmp00_55_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410056(.x(x_56), .z(tmp00_56_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410057(.x(x_57), .z(tmp00_57_41));
	booth__006 #(.WIDTH(WIDTH)) mul00410058(.x(x_58), .z(tmp00_58_41));
	booth__002 #(.WIDTH(WIDTH)) mul00410059(.x(x_59), .z(tmp00_59_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410060(.x(x_60), .z(tmp00_60_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410061(.x(x_61), .z(tmp00_61_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410062(.x(x_62), .z(tmp00_62_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410063(.x(x_63), .z(tmp00_63_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410064(.x(x_64), .z(tmp00_64_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410065(.x(x_65), .z(tmp00_65_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410066(.x(x_66), .z(tmp00_66_41));
	booth__006 #(.WIDTH(WIDTH)) mul00410067(.x(x_67), .z(tmp00_67_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410068(.x(x_68), .z(tmp00_68_41));
	booth_0016 #(.WIDTH(WIDTH)) mul00410069(.x(x_69), .z(tmp00_69_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410070(.x(x_70), .z(tmp00_70_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410071(.x(x_71), .z(tmp00_71_41));
	booth_0010 #(.WIDTH(WIDTH)) mul00410072(.x(x_72), .z(tmp00_72_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410073(.x(x_73), .z(tmp00_73_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410074(.x(x_74), .z(tmp00_74_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410075(.x(x_75), .z(tmp00_75_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410076(.x(x_76), .z(tmp00_76_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410077(.x(x_77), .z(tmp00_77_41));
	booth__002 #(.WIDTH(WIDTH)) mul00410078(.x(x_78), .z(tmp00_78_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410079(.x(x_79), .z(tmp00_79_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410080(.x(x_80), .z(tmp00_80_41));
	booth_0002 #(.WIDTH(WIDTH)) mul00410081(.x(x_81), .z(tmp00_81_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410082(.x(x_82), .z(tmp00_82_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410083(.x(x_83), .z(tmp00_83_41));
	booth_0002 #(.WIDTH(WIDTH)) mul00410084(.x(x_84), .z(tmp00_84_41));
	booth__006 #(.WIDTH(WIDTH)) mul00410085(.x(x_85), .z(tmp00_85_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410086(.x(x_86), .z(tmp00_86_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410087(.x(x_87), .z(tmp00_87_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410088(.x(x_88), .z(tmp00_88_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410089(.x(x_89), .z(tmp00_89_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410090(.x(x_90), .z(tmp00_90_41));
	booth_0012 #(.WIDTH(WIDTH)) mul00410091(.x(x_91), .z(tmp00_91_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410092(.x(x_92), .z(tmp00_92_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410093(.x(x_93), .z(tmp00_93_41));
	booth_0010 #(.WIDTH(WIDTH)) mul00410094(.x(x_94), .z(tmp00_94_41));
	booth_0006 #(.WIDTH(WIDTH)) mul00410095(.x(x_95), .z(tmp00_95_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410096(.x(x_96), .z(tmp00_96_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410097(.x(x_97), .z(tmp00_97_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410098(.x(x_98), .z(tmp00_98_41));
	booth__012 #(.WIDTH(WIDTH)) mul00410099(.x(x_99), .z(tmp00_99_41));
	booth__014 #(.WIDTH(WIDTH)) mul00410100(.x(x_100), .z(tmp00_100_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410101(.x(x_101), .z(tmp00_101_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410102(.x(x_102), .z(tmp00_102_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410103(.x(x_103), .z(tmp00_103_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410104(.x(x_104), .z(tmp00_104_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410105(.x(x_105), .z(tmp00_105_41));
	booth_0000 #(.WIDTH(WIDTH)) mul00410106(.x(x_106), .z(tmp00_106_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410107(.x(x_107), .z(tmp00_107_41));
	booth__004 #(.WIDTH(WIDTH)) mul00410108(.x(x_108), .z(tmp00_108_41));
	booth_0002 #(.WIDTH(WIDTH)) mul00410109(.x(x_109), .z(tmp00_109_41));
	booth_0014 #(.WIDTH(WIDTH)) mul00410110(.x(x_110), .z(tmp00_110_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410111(.x(x_111), .z(tmp00_111_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410112(.x(x_112), .z(tmp00_112_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410113(.x(x_113), .z(tmp00_113_41));
	booth__006 #(.WIDTH(WIDTH)) mul00410114(.x(x_114), .z(tmp00_114_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410115(.x(x_115), .z(tmp00_115_41));
	booth_0010 #(.WIDTH(WIDTH)) mul00410116(.x(x_116), .z(tmp00_116_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410117(.x(x_117), .z(tmp00_117_41));
	booth__012 #(.WIDTH(WIDTH)) mul00410118(.x(x_118), .z(tmp00_118_41));
	booth__010 #(.WIDTH(WIDTH)) mul00410119(.x(x_119), .z(tmp00_119_41));
	booth_0012 #(.WIDTH(WIDTH)) mul00410120(.x(x_120), .z(tmp00_120_41));
	booth_0012 #(.WIDTH(WIDTH)) mul00410121(.x(x_121), .z(tmp00_121_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410122(.x(x_122), .z(tmp00_122_41));
	booth_0006 #(.WIDTH(WIDTH)) mul00410123(.x(x_123), .z(tmp00_123_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410124(.x(x_124), .z(tmp00_124_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00410125(.x(x_125), .z(tmp00_125_41));
	booth__008 #(.WIDTH(WIDTH)) mul00410126(.x(x_126), .z(tmp00_126_41));
	booth_0004 #(.WIDTH(WIDTH)) mul00410127(.x(x_127), .z(tmp00_127_41));
	booth_0008 #(.WIDTH(WIDTH)) mul00420000(.x(x_0), .z(tmp00_0_42));
	booth__006 #(.WIDTH(WIDTH)) mul00420001(.x(x_1), .z(tmp00_1_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420002(.x(x_2), .z(tmp00_2_42));
	booth__002 #(.WIDTH(WIDTH)) mul00420003(.x(x_3), .z(tmp00_3_42));
	booth_0020 #(.WIDTH(WIDTH)) mul00420004(.x(x_4), .z(tmp00_4_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420005(.x(x_5), .z(tmp00_5_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420006(.x(x_6), .z(tmp00_6_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420007(.x(x_7), .z(tmp00_7_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420008(.x(x_8), .z(tmp00_8_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420009(.x(x_9), .z(tmp00_9_42));
	booth__002 #(.WIDTH(WIDTH)) mul00420010(.x(x_10), .z(tmp00_10_42));
	booth__002 #(.WIDTH(WIDTH)) mul00420011(.x(x_11), .z(tmp00_11_42));
	booth__006 #(.WIDTH(WIDTH)) mul00420012(.x(x_12), .z(tmp00_12_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420013(.x(x_13), .z(tmp00_13_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420014(.x(x_14), .z(tmp00_14_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420015(.x(x_15), .z(tmp00_15_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420016(.x(x_16), .z(tmp00_16_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420017(.x(x_17), .z(tmp00_17_42));
	booth__012 #(.WIDTH(WIDTH)) mul00420018(.x(x_18), .z(tmp00_18_42));
	booth__012 #(.WIDTH(WIDTH)) mul00420019(.x(x_19), .z(tmp00_19_42));
	booth_0012 #(.WIDTH(WIDTH)) mul00420020(.x(x_20), .z(tmp00_20_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420021(.x(x_21), .z(tmp00_21_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420022(.x(x_22), .z(tmp00_22_42));
	booth_0006 #(.WIDTH(WIDTH)) mul00420023(.x(x_23), .z(tmp00_23_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420024(.x(x_24), .z(tmp00_24_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420025(.x(x_25), .z(tmp00_25_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420026(.x(x_26), .z(tmp00_26_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420027(.x(x_27), .z(tmp00_27_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420028(.x(x_28), .z(tmp00_28_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420029(.x(x_29), .z(tmp00_29_42));
	booth__016 #(.WIDTH(WIDTH)) mul00420030(.x(x_30), .z(tmp00_30_42));
	booth_0010 #(.WIDTH(WIDTH)) mul00420031(.x(x_31), .z(tmp00_31_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420032(.x(x_32), .z(tmp00_32_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420033(.x(x_33), .z(tmp00_33_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420034(.x(x_34), .z(tmp00_34_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420035(.x(x_35), .z(tmp00_35_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420036(.x(x_36), .z(tmp00_36_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420037(.x(x_37), .z(tmp00_37_42));
	booth_0012 #(.WIDTH(WIDTH)) mul00420038(.x(x_38), .z(tmp00_38_42));
	booth__016 #(.WIDTH(WIDTH)) mul00420039(.x(x_39), .z(tmp00_39_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420040(.x(x_40), .z(tmp00_40_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420041(.x(x_41), .z(tmp00_41_42));
	booth_0016 #(.WIDTH(WIDTH)) mul00420042(.x(x_42), .z(tmp00_42_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420043(.x(x_43), .z(tmp00_43_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420044(.x(x_44), .z(tmp00_44_42));
	booth_0006 #(.WIDTH(WIDTH)) mul00420045(.x(x_45), .z(tmp00_45_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420046(.x(x_46), .z(tmp00_46_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420047(.x(x_47), .z(tmp00_47_42));
	booth__002 #(.WIDTH(WIDTH)) mul00420048(.x(x_48), .z(tmp00_48_42));
	booth__002 #(.WIDTH(WIDTH)) mul00420049(.x(x_49), .z(tmp00_49_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420050(.x(x_50), .z(tmp00_50_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420051(.x(x_51), .z(tmp00_51_42));
	booth_0014 #(.WIDTH(WIDTH)) mul00420052(.x(x_52), .z(tmp00_52_42));
	booth__010 #(.WIDTH(WIDTH)) mul00420053(.x(x_53), .z(tmp00_53_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420054(.x(x_54), .z(tmp00_54_42));
	booth_0014 #(.WIDTH(WIDTH)) mul00420055(.x(x_55), .z(tmp00_55_42));
	booth_0024 #(.WIDTH(WIDTH)) mul00420056(.x(x_56), .z(tmp00_56_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420057(.x(x_57), .z(tmp00_57_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420058(.x(x_58), .z(tmp00_58_42));
	booth__002 #(.WIDTH(WIDTH)) mul00420059(.x(x_59), .z(tmp00_59_42));
	booth_0010 #(.WIDTH(WIDTH)) mul00420060(.x(x_60), .z(tmp00_60_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420061(.x(x_61), .z(tmp00_61_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420062(.x(x_62), .z(tmp00_62_42));
	booth_0012 #(.WIDTH(WIDTH)) mul00420063(.x(x_63), .z(tmp00_63_42));
	booth_0002 #(.WIDTH(WIDTH)) mul00420064(.x(x_64), .z(tmp00_64_42));
	booth_0002 #(.WIDTH(WIDTH)) mul00420065(.x(x_65), .z(tmp00_65_42));
	booth_0016 #(.WIDTH(WIDTH)) mul00420066(.x(x_66), .z(tmp00_66_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420067(.x(x_67), .z(tmp00_67_42));
	booth_0020 #(.WIDTH(WIDTH)) mul00420068(.x(x_68), .z(tmp00_68_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420069(.x(x_69), .z(tmp00_69_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420070(.x(x_70), .z(tmp00_70_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420071(.x(x_71), .z(tmp00_71_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420072(.x(x_72), .z(tmp00_72_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420073(.x(x_73), .z(tmp00_73_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420074(.x(x_74), .z(tmp00_74_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420075(.x(x_75), .z(tmp00_75_42));
	booth__012 #(.WIDTH(WIDTH)) mul00420076(.x(x_76), .z(tmp00_76_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420077(.x(x_77), .z(tmp00_77_42));
	booth__006 #(.WIDTH(WIDTH)) mul00420078(.x(x_78), .z(tmp00_78_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420079(.x(x_79), .z(tmp00_79_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420080(.x(x_80), .z(tmp00_80_42));
	booth_0020 #(.WIDTH(WIDTH)) mul00420081(.x(x_81), .z(tmp00_81_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420082(.x(x_82), .z(tmp00_82_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420083(.x(x_83), .z(tmp00_83_42));
	booth__006 #(.WIDTH(WIDTH)) mul00420084(.x(x_84), .z(tmp00_84_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420085(.x(x_85), .z(tmp00_85_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420086(.x(x_86), .z(tmp00_86_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420087(.x(x_87), .z(tmp00_87_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420088(.x(x_88), .z(tmp00_88_42));
	booth_0016 #(.WIDTH(WIDTH)) mul00420089(.x(x_89), .z(tmp00_89_42));
	booth_0004 #(.WIDTH(WIDTH)) mul00420090(.x(x_90), .z(tmp00_90_42));
	booth_0016 #(.WIDTH(WIDTH)) mul00420091(.x(x_91), .z(tmp00_91_42));
	booth__012 #(.WIDTH(WIDTH)) mul00420092(.x(x_92), .z(tmp00_92_42));
	booth__010 #(.WIDTH(WIDTH)) mul00420093(.x(x_93), .z(tmp00_93_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420094(.x(x_94), .z(tmp00_94_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420095(.x(x_95), .z(tmp00_95_42));
	booth__002 #(.WIDTH(WIDTH)) mul00420096(.x(x_96), .z(tmp00_96_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420097(.x(x_97), .z(tmp00_97_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420098(.x(x_98), .z(tmp00_98_42));
	booth__012 #(.WIDTH(WIDTH)) mul00420099(.x(x_99), .z(tmp00_99_42));
	booth__016 #(.WIDTH(WIDTH)) mul00420100(.x(x_100), .z(tmp00_100_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420101(.x(x_101), .z(tmp00_101_42));
	booth__012 #(.WIDTH(WIDTH)) mul00420102(.x(x_102), .z(tmp00_102_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420103(.x(x_103), .z(tmp00_103_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420104(.x(x_104), .z(tmp00_104_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420105(.x(x_105), .z(tmp00_105_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420106(.x(x_106), .z(tmp00_106_42));
	booth__008 #(.WIDTH(WIDTH)) mul00420107(.x(x_107), .z(tmp00_107_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420108(.x(x_108), .z(tmp00_108_42));
	booth__016 #(.WIDTH(WIDTH)) mul00420109(.x(x_109), .z(tmp00_109_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420110(.x(x_110), .z(tmp00_110_42));
	booth_0008 #(.WIDTH(WIDTH)) mul00420111(.x(x_111), .z(tmp00_111_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420112(.x(x_112), .z(tmp00_112_42));
	booth_0016 #(.WIDTH(WIDTH)) mul00420113(.x(x_113), .z(tmp00_113_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420114(.x(x_114), .z(tmp00_114_42));
	booth_0010 #(.WIDTH(WIDTH)) mul00420115(.x(x_115), .z(tmp00_115_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420116(.x(x_116), .z(tmp00_116_42));
	booth__006 #(.WIDTH(WIDTH)) mul00420117(.x(x_117), .z(tmp00_117_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420118(.x(x_118), .z(tmp00_118_42));
	booth_0012 #(.WIDTH(WIDTH)) mul00420119(.x(x_119), .z(tmp00_119_42));
	booth_0012 #(.WIDTH(WIDTH)) mul00420120(.x(x_120), .z(tmp00_120_42));
	booth__006 #(.WIDTH(WIDTH)) mul00420121(.x(x_121), .z(tmp00_121_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420122(.x(x_122), .z(tmp00_122_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420123(.x(x_123), .z(tmp00_123_42));
	booth__004 #(.WIDTH(WIDTH)) mul00420124(.x(x_124), .z(tmp00_124_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420125(.x(x_125), .z(tmp00_125_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420126(.x(x_126), .z(tmp00_126_42));
	booth_0000 #(.WIDTH(WIDTH)) mul00420127(.x(x_127), .z(tmp00_127_42));
	booth__008 #(.WIDTH(WIDTH)) mul00430000(.x(x_0), .z(tmp00_0_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430001(.x(x_1), .z(tmp00_1_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430002(.x(x_2), .z(tmp00_2_43));
	booth_0010 #(.WIDTH(WIDTH)) mul00430003(.x(x_3), .z(tmp00_3_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430004(.x(x_4), .z(tmp00_4_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430005(.x(x_5), .z(tmp00_5_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430006(.x(x_6), .z(tmp00_6_43));
	booth__012 #(.WIDTH(WIDTH)) mul00430007(.x(x_7), .z(tmp00_7_43));
	booth_0014 #(.WIDTH(WIDTH)) mul00430008(.x(x_8), .z(tmp00_8_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430009(.x(x_9), .z(tmp00_9_43));
	booth__006 #(.WIDTH(WIDTH)) mul00430010(.x(x_10), .z(tmp00_10_43));
	booth_0010 #(.WIDTH(WIDTH)) mul00430011(.x(x_11), .z(tmp00_11_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430012(.x(x_12), .z(tmp00_12_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430013(.x(x_13), .z(tmp00_13_43));
	booth_0004 #(.WIDTH(WIDTH)) mul00430014(.x(x_14), .z(tmp00_14_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430015(.x(x_15), .z(tmp00_15_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430016(.x(x_16), .z(tmp00_16_43));
	booth__010 #(.WIDTH(WIDTH)) mul00430017(.x(x_17), .z(tmp00_17_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430018(.x(x_18), .z(tmp00_18_43));
	booth_0012 #(.WIDTH(WIDTH)) mul00430019(.x(x_19), .z(tmp00_19_43));
	booth_0010 #(.WIDTH(WIDTH)) mul00430020(.x(x_20), .z(tmp00_20_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430021(.x(x_21), .z(tmp00_21_43));
	booth_0004 #(.WIDTH(WIDTH)) mul00430022(.x(x_22), .z(tmp00_22_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430023(.x(x_23), .z(tmp00_23_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430024(.x(x_24), .z(tmp00_24_43));
	booth__012 #(.WIDTH(WIDTH)) mul00430025(.x(x_25), .z(tmp00_25_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430026(.x(x_26), .z(tmp00_26_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430027(.x(x_27), .z(tmp00_27_43));
	booth_0004 #(.WIDTH(WIDTH)) mul00430028(.x(x_28), .z(tmp00_28_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430029(.x(x_29), .z(tmp00_29_43));
	booth_0002 #(.WIDTH(WIDTH)) mul00430030(.x(x_30), .z(tmp00_30_43));
	booth__004 #(.WIDTH(WIDTH)) mul00430031(.x(x_31), .z(tmp00_31_43));
	booth_0002 #(.WIDTH(WIDTH)) mul00430032(.x(x_32), .z(tmp00_32_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430033(.x(x_33), .z(tmp00_33_43));
	booth__010 #(.WIDTH(WIDTH)) mul00430034(.x(x_34), .z(tmp00_34_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430035(.x(x_35), .z(tmp00_35_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430036(.x(x_36), .z(tmp00_36_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430037(.x(x_37), .z(tmp00_37_43));
	booth_0020 #(.WIDTH(WIDTH)) mul00430038(.x(x_38), .z(tmp00_38_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430039(.x(x_39), .z(tmp00_39_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430040(.x(x_40), .z(tmp00_40_43));
	booth_0016 #(.WIDTH(WIDTH)) mul00430041(.x(x_41), .z(tmp00_41_43));
	booth__004 #(.WIDTH(WIDTH)) mul00430042(.x(x_42), .z(tmp00_42_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430043(.x(x_43), .z(tmp00_43_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430044(.x(x_44), .z(tmp00_44_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430045(.x(x_45), .z(tmp00_45_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430046(.x(x_46), .z(tmp00_46_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430047(.x(x_47), .z(tmp00_47_43));
	booth__010 #(.WIDTH(WIDTH)) mul00430048(.x(x_48), .z(tmp00_48_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430049(.x(x_49), .z(tmp00_49_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430050(.x(x_50), .z(tmp00_50_43));
	booth_0006 #(.WIDTH(WIDTH)) mul00430051(.x(x_51), .z(tmp00_51_43));
	booth_0012 #(.WIDTH(WIDTH)) mul00430052(.x(x_52), .z(tmp00_52_43));
	booth_0010 #(.WIDTH(WIDTH)) mul00430053(.x(x_53), .z(tmp00_53_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430054(.x(x_54), .z(tmp00_54_43));
	booth_0006 #(.WIDTH(WIDTH)) mul00430055(.x(x_55), .z(tmp00_55_43));
	booth__010 #(.WIDTH(WIDTH)) mul00430056(.x(x_56), .z(tmp00_56_43));
	booth_0004 #(.WIDTH(WIDTH)) mul00430057(.x(x_57), .z(tmp00_57_43));
	booth_0016 #(.WIDTH(WIDTH)) mul00430058(.x(x_58), .z(tmp00_58_43));
	booth_0004 #(.WIDTH(WIDTH)) mul00430059(.x(x_59), .z(tmp00_59_43));
	booth_0006 #(.WIDTH(WIDTH)) mul00430060(.x(x_60), .z(tmp00_60_43));
	booth__004 #(.WIDTH(WIDTH)) mul00430061(.x(x_61), .z(tmp00_61_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430062(.x(x_62), .z(tmp00_62_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430063(.x(x_63), .z(tmp00_63_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430064(.x(x_64), .z(tmp00_64_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430065(.x(x_65), .z(tmp00_65_43));
	booth_0016 #(.WIDTH(WIDTH)) mul00430066(.x(x_66), .z(tmp00_66_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430067(.x(x_67), .z(tmp00_67_43));
	booth__012 #(.WIDTH(WIDTH)) mul00430068(.x(x_68), .z(tmp00_68_43));
	booth__004 #(.WIDTH(WIDTH)) mul00430069(.x(x_69), .z(tmp00_69_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430070(.x(x_70), .z(tmp00_70_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430071(.x(x_71), .z(tmp00_71_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430072(.x(x_72), .z(tmp00_72_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430073(.x(x_73), .z(tmp00_73_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430074(.x(x_74), .z(tmp00_74_43));
	booth_0016 #(.WIDTH(WIDTH)) mul00430075(.x(x_75), .z(tmp00_75_43));
	booth__004 #(.WIDTH(WIDTH)) mul00430076(.x(x_76), .z(tmp00_76_43));
	booth__002 #(.WIDTH(WIDTH)) mul00430077(.x(x_77), .z(tmp00_77_43));
	booth_0004 #(.WIDTH(WIDTH)) mul00430078(.x(x_78), .z(tmp00_78_43));
	booth__002 #(.WIDTH(WIDTH)) mul00430079(.x(x_79), .z(tmp00_79_43));
	booth__004 #(.WIDTH(WIDTH)) mul00430080(.x(x_80), .z(tmp00_80_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430081(.x(x_81), .z(tmp00_81_43));
	booth__004 #(.WIDTH(WIDTH)) mul00430082(.x(x_82), .z(tmp00_82_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430083(.x(x_83), .z(tmp00_83_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430084(.x(x_84), .z(tmp00_84_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430085(.x(x_85), .z(tmp00_85_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430086(.x(x_86), .z(tmp00_86_43));
	booth_0004 #(.WIDTH(WIDTH)) mul00430087(.x(x_87), .z(tmp00_87_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430088(.x(x_88), .z(tmp00_88_43));
	booth__012 #(.WIDTH(WIDTH)) mul00430089(.x(x_89), .z(tmp00_89_43));
	booth__016 #(.WIDTH(WIDTH)) mul00430090(.x(x_90), .z(tmp00_90_43));
	booth__016 #(.WIDTH(WIDTH)) mul00430091(.x(x_91), .z(tmp00_91_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430092(.x(x_92), .z(tmp00_92_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430093(.x(x_93), .z(tmp00_93_43));
	booth_0010 #(.WIDTH(WIDTH)) mul00430094(.x(x_94), .z(tmp00_94_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430095(.x(x_95), .z(tmp00_95_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430096(.x(x_96), .z(tmp00_96_43));
	booth_0002 #(.WIDTH(WIDTH)) mul00430097(.x(x_97), .z(tmp00_97_43));
	booth__012 #(.WIDTH(WIDTH)) mul00430098(.x(x_98), .z(tmp00_98_43));
	booth_0012 #(.WIDTH(WIDTH)) mul00430099(.x(x_99), .z(tmp00_99_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430100(.x(x_100), .z(tmp00_100_43));
	booth__012 #(.WIDTH(WIDTH)) mul00430101(.x(x_101), .z(tmp00_101_43));
	booth_0012 #(.WIDTH(WIDTH)) mul00430102(.x(x_102), .z(tmp00_102_43));
	booth__004 #(.WIDTH(WIDTH)) mul00430103(.x(x_103), .z(tmp00_103_43));
	booth_0006 #(.WIDTH(WIDTH)) mul00430104(.x(x_104), .z(tmp00_104_43));
	booth_0004 #(.WIDTH(WIDTH)) mul00430105(.x(x_105), .z(tmp00_105_43));
	booth__008 #(.WIDTH(WIDTH)) mul00430106(.x(x_106), .z(tmp00_106_43));
	booth__006 #(.WIDTH(WIDTH)) mul00430107(.x(x_107), .z(tmp00_107_43));
	booth_0010 #(.WIDTH(WIDTH)) mul00430108(.x(x_108), .z(tmp00_108_43));
	booth_0016 #(.WIDTH(WIDTH)) mul00430109(.x(x_109), .z(tmp00_109_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430110(.x(x_110), .z(tmp00_110_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430111(.x(x_111), .z(tmp00_111_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430112(.x(x_112), .z(tmp00_112_43));
	booth__016 #(.WIDTH(WIDTH)) mul00430113(.x(x_113), .z(tmp00_113_43));
	booth__010 #(.WIDTH(WIDTH)) mul00430114(.x(x_114), .z(tmp00_114_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430115(.x(x_115), .z(tmp00_115_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430116(.x(x_116), .z(tmp00_116_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430117(.x(x_117), .z(tmp00_117_43));
	booth_0012 #(.WIDTH(WIDTH)) mul00430118(.x(x_118), .z(tmp00_118_43));
	booth_0008 #(.WIDTH(WIDTH)) mul00430119(.x(x_119), .z(tmp00_119_43));
	booth__016 #(.WIDTH(WIDTH)) mul00430120(.x(x_120), .z(tmp00_120_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430121(.x(x_121), .z(tmp00_121_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430122(.x(x_122), .z(tmp00_122_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430123(.x(x_123), .z(tmp00_123_43));
	booth_0000 #(.WIDTH(WIDTH)) mul00430124(.x(x_124), .z(tmp00_124_43));
	booth__010 #(.WIDTH(WIDTH)) mul00430125(.x(x_125), .z(tmp00_125_43));
	booth_0014 #(.WIDTH(WIDTH)) mul00430126(.x(x_126), .z(tmp00_126_43));
	booth_0016 #(.WIDTH(WIDTH)) mul00430127(.x(x_127), .z(tmp00_127_43));
	booth__008 #(.WIDTH(WIDTH)) mul00440000(.x(x_0), .z(tmp00_0_44));
	booth_0010 #(.WIDTH(WIDTH)) mul00440001(.x(x_1), .z(tmp00_1_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440002(.x(x_2), .z(tmp00_2_44));
	booth_0012 #(.WIDTH(WIDTH)) mul00440003(.x(x_3), .z(tmp00_3_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440004(.x(x_4), .z(tmp00_4_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440005(.x(x_5), .z(tmp00_5_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440006(.x(x_6), .z(tmp00_6_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440007(.x(x_7), .z(tmp00_7_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440008(.x(x_8), .z(tmp00_8_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440009(.x(x_9), .z(tmp00_9_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440010(.x(x_10), .z(tmp00_10_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440011(.x(x_11), .z(tmp00_11_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440012(.x(x_12), .z(tmp00_12_44));
	booth__010 #(.WIDTH(WIDTH)) mul00440013(.x(x_13), .z(tmp00_13_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440014(.x(x_14), .z(tmp00_14_44));
	booth__012 #(.WIDTH(WIDTH)) mul00440015(.x(x_15), .z(tmp00_15_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440016(.x(x_16), .z(tmp00_16_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440017(.x(x_17), .z(tmp00_17_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440018(.x(x_18), .z(tmp00_18_44));
	booth__012 #(.WIDTH(WIDTH)) mul00440019(.x(x_19), .z(tmp00_19_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440020(.x(x_20), .z(tmp00_20_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440021(.x(x_21), .z(tmp00_21_44));
	booth__006 #(.WIDTH(WIDTH)) mul00440022(.x(x_22), .z(tmp00_22_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440023(.x(x_23), .z(tmp00_23_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440024(.x(x_24), .z(tmp00_24_44));
	booth__010 #(.WIDTH(WIDTH)) mul00440025(.x(x_25), .z(tmp00_25_44));
	booth_0010 #(.WIDTH(WIDTH)) mul00440026(.x(x_26), .z(tmp00_26_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440027(.x(x_27), .z(tmp00_27_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440028(.x(x_28), .z(tmp00_28_44));
	booth__010 #(.WIDTH(WIDTH)) mul00440029(.x(x_29), .z(tmp00_29_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440030(.x(x_30), .z(tmp00_30_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440031(.x(x_31), .z(tmp00_31_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440032(.x(x_32), .z(tmp00_32_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440033(.x(x_33), .z(tmp00_33_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440034(.x(x_34), .z(tmp00_34_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440035(.x(x_35), .z(tmp00_35_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440036(.x(x_36), .z(tmp00_36_44));
	booth__002 #(.WIDTH(WIDTH)) mul00440037(.x(x_37), .z(tmp00_37_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440038(.x(x_38), .z(tmp00_38_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440039(.x(x_39), .z(tmp00_39_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440040(.x(x_40), .z(tmp00_40_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440041(.x(x_41), .z(tmp00_41_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440042(.x(x_42), .z(tmp00_42_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440043(.x(x_43), .z(tmp00_43_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440044(.x(x_44), .z(tmp00_44_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440045(.x(x_45), .z(tmp00_45_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440046(.x(x_46), .z(tmp00_46_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440047(.x(x_47), .z(tmp00_47_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440048(.x(x_48), .z(tmp00_48_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440049(.x(x_49), .z(tmp00_49_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440050(.x(x_50), .z(tmp00_50_44));
	booth__006 #(.WIDTH(WIDTH)) mul00440051(.x(x_51), .z(tmp00_51_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440052(.x(x_52), .z(tmp00_52_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440053(.x(x_53), .z(tmp00_53_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440054(.x(x_54), .z(tmp00_54_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440055(.x(x_55), .z(tmp00_55_44));
	booth_0002 #(.WIDTH(WIDTH)) mul00440056(.x(x_56), .z(tmp00_56_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440057(.x(x_57), .z(tmp00_57_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440058(.x(x_58), .z(tmp00_58_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440059(.x(x_59), .z(tmp00_59_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440060(.x(x_60), .z(tmp00_60_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440061(.x(x_61), .z(tmp00_61_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440062(.x(x_62), .z(tmp00_62_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440063(.x(x_63), .z(tmp00_63_44));
	booth__002 #(.WIDTH(WIDTH)) mul00440064(.x(x_64), .z(tmp00_64_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440065(.x(x_65), .z(tmp00_65_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440066(.x(x_66), .z(tmp00_66_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440067(.x(x_67), .z(tmp00_67_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440068(.x(x_68), .z(tmp00_68_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440069(.x(x_69), .z(tmp00_69_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440070(.x(x_70), .z(tmp00_70_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440071(.x(x_71), .z(tmp00_71_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440072(.x(x_72), .z(tmp00_72_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440073(.x(x_73), .z(tmp00_73_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440074(.x(x_74), .z(tmp00_74_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440075(.x(x_75), .z(tmp00_75_44));
	booth__010 #(.WIDTH(WIDTH)) mul00440076(.x(x_76), .z(tmp00_76_44));
	booth__010 #(.WIDTH(WIDTH)) mul00440077(.x(x_77), .z(tmp00_77_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440078(.x(x_78), .z(tmp00_78_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440079(.x(x_79), .z(tmp00_79_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440080(.x(x_80), .z(tmp00_80_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440081(.x(x_81), .z(tmp00_81_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440082(.x(x_82), .z(tmp00_82_44));
	booth__002 #(.WIDTH(WIDTH)) mul00440083(.x(x_83), .z(tmp00_83_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440084(.x(x_84), .z(tmp00_84_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440085(.x(x_85), .z(tmp00_85_44));
	booth_0002 #(.WIDTH(WIDTH)) mul00440086(.x(x_86), .z(tmp00_86_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440087(.x(x_87), .z(tmp00_87_44));
	booth__006 #(.WIDTH(WIDTH)) mul00440088(.x(x_88), .z(tmp00_88_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440089(.x(x_89), .z(tmp00_89_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440090(.x(x_90), .z(tmp00_90_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440091(.x(x_91), .z(tmp00_91_44));
	booth_0010 #(.WIDTH(WIDTH)) mul00440092(.x(x_92), .z(tmp00_92_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440093(.x(x_93), .z(tmp00_93_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440094(.x(x_94), .z(tmp00_94_44));
	booth__010 #(.WIDTH(WIDTH)) mul00440095(.x(x_95), .z(tmp00_95_44));
	booth__002 #(.WIDTH(WIDTH)) mul00440096(.x(x_96), .z(tmp00_96_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440097(.x(x_97), .z(tmp00_97_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440098(.x(x_98), .z(tmp00_98_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440099(.x(x_99), .z(tmp00_99_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440100(.x(x_100), .z(tmp00_100_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440101(.x(x_101), .z(tmp00_101_44));
	booth_0010 #(.WIDTH(WIDTH)) mul00440102(.x(x_102), .z(tmp00_102_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440103(.x(x_103), .z(tmp00_103_44));
	booth_0010 #(.WIDTH(WIDTH)) mul00440104(.x(x_104), .z(tmp00_104_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440105(.x(x_105), .z(tmp00_105_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440106(.x(x_106), .z(tmp00_106_44));
	booth_0010 #(.WIDTH(WIDTH)) mul00440107(.x(x_107), .z(tmp00_107_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440108(.x(x_108), .z(tmp00_108_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440109(.x(x_109), .z(tmp00_109_44));
	booth__006 #(.WIDTH(WIDTH)) mul00440110(.x(x_110), .z(tmp00_110_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440111(.x(x_111), .z(tmp00_111_44));
	booth_0002 #(.WIDTH(WIDTH)) mul00440112(.x(x_112), .z(tmp00_112_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440113(.x(x_113), .z(tmp00_113_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440114(.x(x_114), .z(tmp00_114_44));
	booth__008 #(.WIDTH(WIDTH)) mul00440115(.x(x_115), .z(tmp00_115_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440116(.x(x_116), .z(tmp00_116_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440117(.x(x_117), .z(tmp00_117_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440118(.x(x_118), .z(tmp00_118_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440119(.x(x_119), .z(tmp00_119_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440120(.x(x_120), .z(tmp00_120_44));
	booth_0004 #(.WIDTH(WIDTH)) mul00440121(.x(x_121), .z(tmp00_121_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440122(.x(x_122), .z(tmp00_122_44));
	booth_0000 #(.WIDTH(WIDTH)) mul00440123(.x(x_123), .z(tmp00_123_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440124(.x(x_124), .z(tmp00_124_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440125(.x(x_125), .z(tmp00_125_44));
	booth_0008 #(.WIDTH(WIDTH)) mul00440126(.x(x_126), .z(tmp00_126_44));
	booth__004 #(.WIDTH(WIDTH)) mul00440127(.x(x_127), .z(tmp00_127_44));
	booth_0006 #(.WIDTH(WIDTH)) mul00450000(.x(x_0), .z(tmp00_0_45));
	booth_0012 #(.WIDTH(WIDTH)) mul00450001(.x(x_1), .z(tmp00_1_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450002(.x(x_2), .z(tmp00_2_45));
	booth_0002 #(.WIDTH(WIDTH)) mul00450003(.x(x_3), .z(tmp00_3_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450004(.x(x_4), .z(tmp00_4_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450005(.x(x_5), .z(tmp00_5_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450006(.x(x_6), .z(tmp00_6_45));
	booth_0002 #(.WIDTH(WIDTH)) mul00450007(.x(x_7), .z(tmp00_7_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450008(.x(x_8), .z(tmp00_8_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450009(.x(x_9), .z(tmp00_9_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450010(.x(x_10), .z(tmp00_10_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450011(.x(x_11), .z(tmp00_11_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450012(.x(x_12), .z(tmp00_12_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450013(.x(x_13), .z(tmp00_13_45));
	booth__006 #(.WIDTH(WIDTH)) mul00450014(.x(x_14), .z(tmp00_14_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450015(.x(x_15), .z(tmp00_15_45));
	booth_0010 #(.WIDTH(WIDTH)) mul00450016(.x(x_16), .z(tmp00_16_45));
	booth_0010 #(.WIDTH(WIDTH)) mul00450017(.x(x_17), .z(tmp00_17_45));
	booth__002 #(.WIDTH(WIDTH)) mul00450018(.x(x_18), .z(tmp00_18_45));
	booth_0014 #(.WIDTH(WIDTH)) mul00450019(.x(x_19), .z(tmp00_19_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450020(.x(x_20), .z(tmp00_20_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450021(.x(x_21), .z(tmp00_21_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450022(.x(x_22), .z(tmp00_22_45));
	booth_0006 #(.WIDTH(WIDTH)) mul00450023(.x(x_23), .z(tmp00_23_45));
	booth__002 #(.WIDTH(WIDTH)) mul00450024(.x(x_24), .z(tmp00_24_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450025(.x(x_25), .z(tmp00_25_45));
	booth__002 #(.WIDTH(WIDTH)) mul00450026(.x(x_26), .z(tmp00_26_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450027(.x(x_27), .z(tmp00_27_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450028(.x(x_28), .z(tmp00_28_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450029(.x(x_29), .z(tmp00_29_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450030(.x(x_30), .z(tmp00_30_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450031(.x(x_31), .z(tmp00_31_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450032(.x(x_32), .z(tmp00_32_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450033(.x(x_33), .z(tmp00_33_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450034(.x(x_34), .z(tmp00_34_45));
	booth_0006 #(.WIDTH(WIDTH)) mul00450035(.x(x_35), .z(tmp00_35_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450036(.x(x_36), .z(tmp00_36_45));
	booth_0006 #(.WIDTH(WIDTH)) mul00450037(.x(x_37), .z(tmp00_37_45));
	booth_0006 #(.WIDTH(WIDTH)) mul00450038(.x(x_38), .z(tmp00_38_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450039(.x(x_39), .z(tmp00_39_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450040(.x(x_40), .z(tmp00_40_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450041(.x(x_41), .z(tmp00_41_45));
	booth_0006 #(.WIDTH(WIDTH)) mul00450042(.x(x_42), .z(tmp00_42_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450043(.x(x_43), .z(tmp00_43_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450044(.x(x_44), .z(tmp00_44_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450045(.x(x_45), .z(tmp00_45_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450046(.x(x_46), .z(tmp00_46_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450047(.x(x_47), .z(tmp00_47_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450048(.x(x_48), .z(tmp00_48_45));
	booth_0016 #(.WIDTH(WIDTH)) mul00450049(.x(x_49), .z(tmp00_49_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450050(.x(x_50), .z(tmp00_50_45));
	booth_0006 #(.WIDTH(WIDTH)) mul00450051(.x(x_51), .z(tmp00_51_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450052(.x(x_52), .z(tmp00_52_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450053(.x(x_53), .z(tmp00_53_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450054(.x(x_54), .z(tmp00_54_45));
	booth_0006 #(.WIDTH(WIDTH)) mul00450055(.x(x_55), .z(tmp00_55_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450056(.x(x_56), .z(tmp00_56_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450057(.x(x_57), .z(tmp00_57_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450058(.x(x_58), .z(tmp00_58_45));
	booth_0018 #(.WIDTH(WIDTH)) mul00450059(.x(x_59), .z(tmp00_59_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450060(.x(x_60), .z(tmp00_60_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450061(.x(x_61), .z(tmp00_61_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450062(.x(x_62), .z(tmp00_62_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450063(.x(x_63), .z(tmp00_63_45));
	booth__006 #(.WIDTH(WIDTH)) mul00450064(.x(x_64), .z(tmp00_64_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450065(.x(x_65), .z(tmp00_65_45));
	booth_0014 #(.WIDTH(WIDTH)) mul00450066(.x(x_66), .z(tmp00_66_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450067(.x(x_67), .z(tmp00_67_45));
	booth__012 #(.WIDTH(WIDTH)) mul00450068(.x(x_68), .z(tmp00_68_45));
	booth_0006 #(.WIDTH(WIDTH)) mul00450069(.x(x_69), .z(tmp00_69_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450070(.x(x_70), .z(tmp00_70_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450071(.x(x_71), .z(tmp00_71_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450072(.x(x_72), .z(tmp00_72_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450073(.x(x_73), .z(tmp00_73_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450074(.x(x_74), .z(tmp00_74_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450075(.x(x_75), .z(tmp00_75_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450076(.x(x_76), .z(tmp00_76_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450077(.x(x_77), .z(tmp00_77_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450078(.x(x_78), .z(tmp00_78_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450079(.x(x_79), .z(tmp00_79_45));
	booth_0014 #(.WIDTH(WIDTH)) mul00450080(.x(x_80), .z(tmp00_80_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450081(.x(x_81), .z(tmp00_81_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450082(.x(x_82), .z(tmp00_82_45));
	booth__010 #(.WIDTH(WIDTH)) mul00450083(.x(x_83), .z(tmp00_83_45));
	booth_0010 #(.WIDTH(WIDTH)) mul00450084(.x(x_84), .z(tmp00_84_45));
	booth__010 #(.WIDTH(WIDTH)) mul00450085(.x(x_85), .z(tmp00_85_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450086(.x(x_86), .z(tmp00_86_45));
	booth__012 #(.WIDTH(WIDTH)) mul00450087(.x(x_87), .z(tmp00_87_45));
	booth__010 #(.WIDTH(WIDTH)) mul00450088(.x(x_88), .z(tmp00_88_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450089(.x(x_89), .z(tmp00_89_45));
	booth__016 #(.WIDTH(WIDTH)) mul00450090(.x(x_90), .z(tmp00_90_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450091(.x(x_91), .z(tmp00_91_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450092(.x(x_92), .z(tmp00_92_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450093(.x(x_93), .z(tmp00_93_45));
	booth_0002 #(.WIDTH(WIDTH)) mul00450094(.x(x_94), .z(tmp00_94_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450095(.x(x_95), .z(tmp00_95_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450096(.x(x_96), .z(tmp00_96_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450097(.x(x_97), .z(tmp00_97_45));
	booth_0012 #(.WIDTH(WIDTH)) mul00450098(.x(x_98), .z(tmp00_98_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450099(.x(x_99), .z(tmp00_99_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450100(.x(x_100), .z(tmp00_100_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450101(.x(x_101), .z(tmp00_101_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450102(.x(x_102), .z(tmp00_102_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450103(.x(x_103), .z(tmp00_103_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450104(.x(x_104), .z(tmp00_104_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450105(.x(x_105), .z(tmp00_105_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450106(.x(x_106), .z(tmp00_106_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450107(.x(x_107), .z(tmp00_107_45));
	booth__012 #(.WIDTH(WIDTH)) mul00450108(.x(x_108), .z(tmp00_108_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450109(.x(x_109), .z(tmp00_109_45));
	booth__010 #(.WIDTH(WIDTH)) mul00450110(.x(x_110), .z(tmp00_110_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450111(.x(x_111), .z(tmp00_111_45));
	booth__012 #(.WIDTH(WIDTH)) mul00450112(.x(x_112), .z(tmp00_112_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450113(.x(x_113), .z(tmp00_113_45));
	booth_0002 #(.WIDTH(WIDTH)) mul00450114(.x(x_114), .z(tmp00_114_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450115(.x(x_115), .z(tmp00_115_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450116(.x(x_116), .z(tmp00_116_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450117(.x(x_117), .z(tmp00_117_45));
	booth__004 #(.WIDTH(WIDTH)) mul00450118(.x(x_118), .z(tmp00_118_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450119(.x(x_119), .z(tmp00_119_45));
	booth__008 #(.WIDTH(WIDTH)) mul00450120(.x(x_120), .z(tmp00_120_45));
	booth_0020 #(.WIDTH(WIDTH)) mul00450121(.x(x_121), .z(tmp00_121_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450122(.x(x_122), .z(tmp00_122_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450123(.x(x_123), .z(tmp00_123_45));
	booth_0010 #(.WIDTH(WIDTH)) mul00450124(.x(x_124), .z(tmp00_124_45));
	booth_0000 #(.WIDTH(WIDTH)) mul00450125(.x(x_125), .z(tmp00_125_45));
	booth_0004 #(.WIDTH(WIDTH)) mul00450126(.x(x_126), .z(tmp00_126_45));
	booth_0008 #(.WIDTH(WIDTH)) mul00450127(.x(x_127), .z(tmp00_127_45));
	booth__008 #(.WIDTH(WIDTH)) mul00460000(.x(x_0), .z(tmp00_0_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460001(.x(x_1), .z(tmp00_1_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460002(.x(x_2), .z(tmp00_2_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460003(.x(x_3), .z(tmp00_3_46));
	booth_0010 #(.WIDTH(WIDTH)) mul00460004(.x(x_4), .z(tmp00_4_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460005(.x(x_5), .z(tmp00_5_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460006(.x(x_6), .z(tmp00_6_46));
	booth__002 #(.WIDTH(WIDTH)) mul00460007(.x(x_7), .z(tmp00_7_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460008(.x(x_8), .z(tmp00_8_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460009(.x(x_9), .z(tmp00_9_46));
	booth_0010 #(.WIDTH(WIDTH)) mul00460010(.x(x_10), .z(tmp00_10_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460011(.x(x_11), .z(tmp00_11_46));
	booth_0002 #(.WIDTH(WIDTH)) mul00460012(.x(x_12), .z(tmp00_12_46));
	booth__010 #(.WIDTH(WIDTH)) mul00460013(.x(x_13), .z(tmp00_13_46));
	booth__002 #(.WIDTH(WIDTH)) mul00460014(.x(x_14), .z(tmp00_14_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460015(.x(x_15), .z(tmp00_15_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460016(.x(x_16), .z(tmp00_16_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460017(.x(x_17), .z(tmp00_17_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460018(.x(x_18), .z(tmp00_18_46));
	booth_0002 #(.WIDTH(WIDTH)) mul00460019(.x(x_19), .z(tmp00_19_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460020(.x(x_20), .z(tmp00_20_46));
	booth__006 #(.WIDTH(WIDTH)) mul00460021(.x(x_21), .z(tmp00_21_46));
	booth_0010 #(.WIDTH(WIDTH)) mul00460022(.x(x_22), .z(tmp00_22_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460023(.x(x_23), .z(tmp00_23_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460024(.x(x_24), .z(tmp00_24_46));
	booth__006 #(.WIDTH(WIDTH)) mul00460025(.x(x_25), .z(tmp00_25_46));
	booth_0010 #(.WIDTH(WIDTH)) mul00460026(.x(x_26), .z(tmp00_26_46));
	booth_0002 #(.WIDTH(WIDTH)) mul00460027(.x(x_27), .z(tmp00_27_46));
	booth_0006 #(.WIDTH(WIDTH)) mul00460028(.x(x_28), .z(tmp00_28_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460029(.x(x_29), .z(tmp00_29_46));
	booth_0006 #(.WIDTH(WIDTH)) mul00460030(.x(x_30), .z(tmp00_30_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460031(.x(x_31), .z(tmp00_31_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460032(.x(x_32), .z(tmp00_32_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460033(.x(x_33), .z(tmp00_33_46));
	booth_0002 #(.WIDTH(WIDTH)) mul00460034(.x(x_34), .z(tmp00_34_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460035(.x(x_35), .z(tmp00_35_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460036(.x(x_36), .z(tmp00_36_46));
	booth_0002 #(.WIDTH(WIDTH)) mul00460037(.x(x_37), .z(tmp00_37_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460038(.x(x_38), .z(tmp00_38_46));
	booth__002 #(.WIDTH(WIDTH)) mul00460039(.x(x_39), .z(tmp00_39_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460040(.x(x_40), .z(tmp00_40_46));
	booth__012 #(.WIDTH(WIDTH)) mul00460041(.x(x_41), .z(tmp00_41_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460042(.x(x_42), .z(tmp00_42_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460043(.x(x_43), .z(tmp00_43_46));
	booth__006 #(.WIDTH(WIDTH)) mul00460044(.x(x_44), .z(tmp00_44_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460045(.x(x_45), .z(tmp00_45_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460046(.x(x_46), .z(tmp00_46_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460047(.x(x_47), .z(tmp00_47_46));
	booth_0010 #(.WIDTH(WIDTH)) mul00460048(.x(x_48), .z(tmp00_48_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460049(.x(x_49), .z(tmp00_49_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460050(.x(x_50), .z(tmp00_50_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460051(.x(x_51), .z(tmp00_51_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460052(.x(x_52), .z(tmp00_52_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460053(.x(x_53), .z(tmp00_53_46));
	booth__010 #(.WIDTH(WIDTH)) mul00460054(.x(x_54), .z(tmp00_54_46));
	booth_0006 #(.WIDTH(WIDTH)) mul00460055(.x(x_55), .z(tmp00_55_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460056(.x(x_56), .z(tmp00_56_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460057(.x(x_57), .z(tmp00_57_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460058(.x(x_58), .z(tmp00_58_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460059(.x(x_59), .z(tmp00_59_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460060(.x(x_60), .z(tmp00_60_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460061(.x(x_61), .z(tmp00_61_46));
	booth__006 #(.WIDTH(WIDTH)) mul00460062(.x(x_62), .z(tmp00_62_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460063(.x(x_63), .z(tmp00_63_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460064(.x(x_64), .z(tmp00_64_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460065(.x(x_65), .z(tmp00_65_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460066(.x(x_66), .z(tmp00_66_46));
	booth__012 #(.WIDTH(WIDTH)) mul00460067(.x(x_67), .z(tmp00_67_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460068(.x(x_68), .z(tmp00_68_46));
	booth__006 #(.WIDTH(WIDTH)) mul00460069(.x(x_69), .z(tmp00_69_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460070(.x(x_70), .z(tmp00_70_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460071(.x(x_71), .z(tmp00_71_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460072(.x(x_72), .z(tmp00_72_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460073(.x(x_73), .z(tmp00_73_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460074(.x(x_74), .z(tmp00_74_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460075(.x(x_75), .z(tmp00_75_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460076(.x(x_76), .z(tmp00_76_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460077(.x(x_77), .z(tmp00_77_46));
	booth__006 #(.WIDTH(WIDTH)) mul00460078(.x(x_78), .z(tmp00_78_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460079(.x(x_79), .z(tmp00_79_46));
	booth_0006 #(.WIDTH(WIDTH)) mul00460080(.x(x_80), .z(tmp00_80_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460081(.x(x_81), .z(tmp00_81_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460082(.x(x_82), .z(tmp00_82_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460083(.x(x_83), .z(tmp00_83_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460084(.x(x_84), .z(tmp00_84_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460085(.x(x_85), .z(tmp00_85_46));
	booth__012 #(.WIDTH(WIDTH)) mul00460086(.x(x_86), .z(tmp00_86_46));
	booth_0002 #(.WIDTH(WIDTH)) mul00460087(.x(x_87), .z(tmp00_87_46));
	booth_0002 #(.WIDTH(WIDTH)) mul00460088(.x(x_88), .z(tmp00_88_46));
	booth_0006 #(.WIDTH(WIDTH)) mul00460089(.x(x_89), .z(tmp00_89_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460090(.x(x_90), .z(tmp00_90_46));
	booth__006 #(.WIDTH(WIDTH)) mul00460091(.x(x_91), .z(tmp00_91_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460092(.x(x_92), .z(tmp00_92_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460093(.x(x_93), .z(tmp00_93_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460094(.x(x_94), .z(tmp00_94_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460095(.x(x_95), .z(tmp00_95_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460096(.x(x_96), .z(tmp00_96_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460097(.x(x_97), .z(tmp00_97_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460098(.x(x_98), .z(tmp00_98_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460099(.x(x_99), .z(tmp00_99_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460100(.x(x_100), .z(tmp00_100_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460101(.x(x_101), .z(tmp00_101_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460102(.x(x_102), .z(tmp00_102_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460103(.x(x_103), .z(tmp00_103_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460104(.x(x_104), .z(tmp00_104_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460105(.x(x_105), .z(tmp00_105_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460106(.x(x_106), .z(tmp00_106_46));
	booth__004 #(.WIDTH(WIDTH)) mul00460107(.x(x_107), .z(tmp00_107_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460108(.x(x_108), .z(tmp00_108_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460109(.x(x_109), .z(tmp00_109_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460110(.x(x_110), .z(tmp00_110_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460111(.x(x_111), .z(tmp00_111_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460112(.x(x_112), .z(tmp00_112_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460113(.x(x_113), .z(tmp00_113_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460114(.x(x_114), .z(tmp00_114_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460115(.x(x_115), .z(tmp00_115_46));
	booth__002 #(.WIDTH(WIDTH)) mul00460116(.x(x_116), .z(tmp00_116_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460117(.x(x_117), .z(tmp00_117_46));
	booth_0012 #(.WIDTH(WIDTH)) mul00460118(.x(x_118), .z(tmp00_118_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460119(.x(x_119), .z(tmp00_119_46));
	booth__002 #(.WIDTH(WIDTH)) mul00460120(.x(x_120), .z(tmp00_120_46));
	booth_0004 #(.WIDTH(WIDTH)) mul00460121(.x(x_121), .z(tmp00_121_46));
	booth__010 #(.WIDTH(WIDTH)) mul00460122(.x(x_122), .z(tmp00_122_46));
	booth__008 #(.WIDTH(WIDTH)) mul00460123(.x(x_123), .z(tmp00_123_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460124(.x(x_124), .z(tmp00_124_46));
	booth_0008 #(.WIDTH(WIDTH)) mul00460125(.x(x_125), .z(tmp00_125_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00460126(.x(x_126), .z(tmp00_126_46));
	booth__002 #(.WIDTH(WIDTH)) mul00460127(.x(x_127), .z(tmp00_127_46));
	booth_0000 #(.WIDTH(WIDTH)) mul00470000(.x(x_0), .z(tmp00_0_47));
	booth__002 #(.WIDTH(WIDTH)) mul00470001(.x(x_1), .z(tmp00_1_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470002(.x(x_2), .z(tmp00_2_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470003(.x(x_3), .z(tmp00_3_47));
	booth__002 #(.WIDTH(WIDTH)) mul00470004(.x(x_4), .z(tmp00_4_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470005(.x(x_5), .z(tmp00_5_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470006(.x(x_6), .z(tmp00_6_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470007(.x(x_7), .z(tmp00_7_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470008(.x(x_8), .z(tmp00_8_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470009(.x(x_9), .z(tmp00_9_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470010(.x(x_10), .z(tmp00_10_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470011(.x(x_11), .z(tmp00_11_47));
	booth__012 #(.WIDTH(WIDTH)) mul00470012(.x(x_12), .z(tmp00_12_47));
	booth__006 #(.WIDTH(WIDTH)) mul00470013(.x(x_13), .z(tmp00_13_47));
	booth__006 #(.WIDTH(WIDTH)) mul00470014(.x(x_14), .z(tmp00_14_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470015(.x(x_15), .z(tmp00_15_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470016(.x(x_16), .z(tmp00_16_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470017(.x(x_17), .z(tmp00_17_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470018(.x(x_18), .z(tmp00_18_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470019(.x(x_19), .z(tmp00_19_47));
	booth_0002 #(.WIDTH(WIDTH)) mul00470020(.x(x_20), .z(tmp00_20_47));
	booth_0002 #(.WIDTH(WIDTH)) mul00470021(.x(x_21), .z(tmp00_21_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470022(.x(x_22), .z(tmp00_22_47));
	booth_0002 #(.WIDTH(WIDTH)) mul00470023(.x(x_23), .z(tmp00_23_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470024(.x(x_24), .z(tmp00_24_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470025(.x(x_25), .z(tmp00_25_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470026(.x(x_26), .z(tmp00_26_47));
	booth_0002 #(.WIDTH(WIDTH)) mul00470027(.x(x_27), .z(tmp00_27_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470028(.x(x_28), .z(tmp00_28_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470029(.x(x_29), .z(tmp00_29_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470030(.x(x_30), .z(tmp00_30_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470031(.x(x_31), .z(tmp00_31_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470032(.x(x_32), .z(tmp00_32_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470033(.x(x_33), .z(tmp00_33_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470034(.x(x_34), .z(tmp00_34_47));
	booth_0006 #(.WIDTH(WIDTH)) mul00470035(.x(x_35), .z(tmp00_35_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470036(.x(x_36), .z(tmp00_36_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470037(.x(x_37), .z(tmp00_37_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470038(.x(x_38), .z(tmp00_38_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470039(.x(x_39), .z(tmp00_39_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470040(.x(x_40), .z(tmp00_40_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470041(.x(x_41), .z(tmp00_41_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470042(.x(x_42), .z(tmp00_42_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470043(.x(x_43), .z(tmp00_43_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470044(.x(x_44), .z(tmp00_44_47));
	booth_0006 #(.WIDTH(WIDTH)) mul00470045(.x(x_45), .z(tmp00_45_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470046(.x(x_46), .z(tmp00_46_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470047(.x(x_47), .z(tmp00_47_47));
	booth_0010 #(.WIDTH(WIDTH)) mul00470048(.x(x_48), .z(tmp00_48_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470049(.x(x_49), .z(tmp00_49_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470050(.x(x_50), .z(tmp00_50_47));
	booth__006 #(.WIDTH(WIDTH)) mul00470051(.x(x_51), .z(tmp00_51_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470052(.x(x_52), .z(tmp00_52_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470053(.x(x_53), .z(tmp00_53_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470054(.x(x_54), .z(tmp00_54_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470055(.x(x_55), .z(tmp00_55_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470056(.x(x_56), .z(tmp00_56_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470057(.x(x_57), .z(tmp00_57_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470058(.x(x_58), .z(tmp00_58_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470059(.x(x_59), .z(tmp00_59_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470060(.x(x_60), .z(tmp00_60_47));
	booth_0012 #(.WIDTH(WIDTH)) mul00470061(.x(x_61), .z(tmp00_61_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470062(.x(x_62), .z(tmp00_62_47));
	booth__006 #(.WIDTH(WIDTH)) mul00470063(.x(x_63), .z(tmp00_63_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470064(.x(x_64), .z(tmp00_64_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470065(.x(x_65), .z(tmp00_65_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470066(.x(x_66), .z(tmp00_66_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470067(.x(x_67), .z(tmp00_67_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470068(.x(x_68), .z(tmp00_68_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470069(.x(x_69), .z(tmp00_69_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470070(.x(x_70), .z(tmp00_70_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470071(.x(x_71), .z(tmp00_71_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470072(.x(x_72), .z(tmp00_72_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470073(.x(x_73), .z(tmp00_73_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470074(.x(x_74), .z(tmp00_74_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470075(.x(x_75), .z(tmp00_75_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470076(.x(x_76), .z(tmp00_76_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470077(.x(x_77), .z(tmp00_77_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470078(.x(x_78), .z(tmp00_78_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470079(.x(x_79), .z(tmp00_79_47));
	booth_0002 #(.WIDTH(WIDTH)) mul00470080(.x(x_80), .z(tmp00_80_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470081(.x(x_81), .z(tmp00_81_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470082(.x(x_82), .z(tmp00_82_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470083(.x(x_83), .z(tmp00_83_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470084(.x(x_84), .z(tmp00_84_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470085(.x(x_85), .z(tmp00_85_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470086(.x(x_86), .z(tmp00_86_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470087(.x(x_87), .z(tmp00_87_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470088(.x(x_88), .z(tmp00_88_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470089(.x(x_89), .z(tmp00_89_47));
	booth_0002 #(.WIDTH(WIDTH)) mul00470090(.x(x_90), .z(tmp00_90_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470091(.x(x_91), .z(tmp00_91_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470092(.x(x_92), .z(tmp00_92_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470093(.x(x_93), .z(tmp00_93_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470094(.x(x_94), .z(tmp00_94_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470095(.x(x_95), .z(tmp00_95_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470096(.x(x_96), .z(tmp00_96_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470097(.x(x_97), .z(tmp00_97_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470098(.x(x_98), .z(tmp00_98_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470099(.x(x_99), .z(tmp00_99_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470100(.x(x_100), .z(tmp00_100_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470101(.x(x_101), .z(tmp00_101_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470102(.x(x_102), .z(tmp00_102_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470103(.x(x_103), .z(tmp00_103_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470104(.x(x_104), .z(tmp00_104_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470105(.x(x_105), .z(tmp00_105_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470106(.x(x_106), .z(tmp00_106_47));
	booth_0008 #(.WIDTH(WIDTH)) mul00470107(.x(x_107), .z(tmp00_107_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470108(.x(x_108), .z(tmp00_108_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470109(.x(x_109), .z(tmp00_109_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470110(.x(x_110), .z(tmp00_110_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470111(.x(x_111), .z(tmp00_111_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470112(.x(x_112), .z(tmp00_112_47));
	booth__010 #(.WIDTH(WIDTH)) mul00470113(.x(x_113), .z(tmp00_113_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470114(.x(x_114), .z(tmp00_114_47));
	booth_0004 #(.WIDTH(WIDTH)) mul00470115(.x(x_115), .z(tmp00_115_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470116(.x(x_116), .z(tmp00_116_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470117(.x(x_117), .z(tmp00_117_47));
	booth__002 #(.WIDTH(WIDTH)) mul00470118(.x(x_118), .z(tmp00_118_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470119(.x(x_119), .z(tmp00_119_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470120(.x(x_120), .z(tmp00_120_47));
	booth__008 #(.WIDTH(WIDTH)) mul00470121(.x(x_121), .z(tmp00_121_47));
	booth__002 #(.WIDTH(WIDTH)) mul00470122(.x(x_122), .z(tmp00_122_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470123(.x(x_123), .z(tmp00_123_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00470124(.x(x_124), .z(tmp00_124_47));
	booth__004 #(.WIDTH(WIDTH)) mul00470125(.x(x_125), .z(tmp00_125_47));
	booth_0006 #(.WIDTH(WIDTH)) mul00470126(.x(x_126), .z(tmp00_126_47));
	booth_0006 #(.WIDTH(WIDTH)) mul00470127(.x(x_127), .z(tmp00_127_47));
	booth_0000 #(.WIDTH(WIDTH)) mul00480000(.x(x_0), .z(tmp00_0_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480001(.x(x_1), .z(tmp00_1_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480002(.x(x_2), .z(tmp00_2_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480003(.x(x_3), .z(tmp00_3_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480004(.x(x_4), .z(tmp00_4_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480005(.x(x_5), .z(tmp00_5_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480006(.x(x_6), .z(tmp00_6_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480007(.x(x_7), .z(tmp00_7_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480008(.x(x_8), .z(tmp00_8_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480009(.x(x_9), .z(tmp00_9_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480010(.x(x_10), .z(tmp00_10_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480011(.x(x_11), .z(tmp00_11_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480012(.x(x_12), .z(tmp00_12_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480013(.x(x_13), .z(tmp00_13_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480014(.x(x_14), .z(tmp00_14_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480015(.x(x_15), .z(tmp00_15_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480016(.x(x_16), .z(tmp00_16_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480017(.x(x_17), .z(tmp00_17_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480018(.x(x_18), .z(tmp00_18_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480019(.x(x_19), .z(tmp00_19_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480020(.x(x_20), .z(tmp00_20_48));
	booth_0010 #(.WIDTH(WIDTH)) mul00480021(.x(x_21), .z(tmp00_21_48));
	booth_0010 #(.WIDTH(WIDTH)) mul00480022(.x(x_22), .z(tmp00_22_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480023(.x(x_23), .z(tmp00_23_48));
	booth__006 #(.WIDTH(WIDTH)) mul00480024(.x(x_24), .z(tmp00_24_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480025(.x(x_25), .z(tmp00_25_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480026(.x(x_26), .z(tmp00_26_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480027(.x(x_27), .z(tmp00_27_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480028(.x(x_28), .z(tmp00_28_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480029(.x(x_29), .z(tmp00_29_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480030(.x(x_30), .z(tmp00_30_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480031(.x(x_31), .z(tmp00_31_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480032(.x(x_32), .z(tmp00_32_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480033(.x(x_33), .z(tmp00_33_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480034(.x(x_34), .z(tmp00_34_48));
	booth_0006 #(.WIDTH(WIDTH)) mul00480035(.x(x_35), .z(tmp00_35_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480036(.x(x_36), .z(tmp00_36_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480037(.x(x_37), .z(tmp00_37_48));
	booth_0010 #(.WIDTH(WIDTH)) mul00480038(.x(x_38), .z(tmp00_38_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480039(.x(x_39), .z(tmp00_39_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480040(.x(x_40), .z(tmp00_40_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480041(.x(x_41), .z(tmp00_41_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480042(.x(x_42), .z(tmp00_42_48));
	booth__002 #(.WIDTH(WIDTH)) mul00480043(.x(x_43), .z(tmp00_43_48));
	booth__012 #(.WIDTH(WIDTH)) mul00480044(.x(x_44), .z(tmp00_44_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480045(.x(x_45), .z(tmp00_45_48));
	booth__006 #(.WIDTH(WIDTH)) mul00480046(.x(x_46), .z(tmp00_46_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480047(.x(x_47), .z(tmp00_47_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480048(.x(x_48), .z(tmp00_48_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480049(.x(x_49), .z(tmp00_49_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480050(.x(x_50), .z(tmp00_50_48));
	booth_0002 #(.WIDTH(WIDTH)) mul00480051(.x(x_51), .z(tmp00_51_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480052(.x(x_52), .z(tmp00_52_48));
	booth__002 #(.WIDTH(WIDTH)) mul00480053(.x(x_53), .z(tmp00_53_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480054(.x(x_54), .z(tmp00_54_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480055(.x(x_55), .z(tmp00_55_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480056(.x(x_56), .z(tmp00_56_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480057(.x(x_57), .z(tmp00_57_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480058(.x(x_58), .z(tmp00_58_48));
	booth_0002 #(.WIDTH(WIDTH)) mul00480059(.x(x_59), .z(tmp00_59_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480060(.x(x_60), .z(tmp00_60_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480061(.x(x_61), .z(tmp00_61_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480062(.x(x_62), .z(tmp00_62_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480063(.x(x_63), .z(tmp00_63_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480064(.x(x_64), .z(tmp00_64_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480065(.x(x_65), .z(tmp00_65_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480066(.x(x_66), .z(tmp00_66_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480067(.x(x_67), .z(tmp00_67_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480068(.x(x_68), .z(tmp00_68_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480069(.x(x_69), .z(tmp00_69_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480070(.x(x_70), .z(tmp00_70_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480071(.x(x_71), .z(tmp00_71_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480072(.x(x_72), .z(tmp00_72_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480073(.x(x_73), .z(tmp00_73_48));
	booth_0006 #(.WIDTH(WIDTH)) mul00480074(.x(x_74), .z(tmp00_74_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480075(.x(x_75), .z(tmp00_75_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480076(.x(x_76), .z(tmp00_76_48));
	booth_0002 #(.WIDTH(WIDTH)) mul00480077(.x(x_77), .z(tmp00_77_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480078(.x(x_78), .z(tmp00_78_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480079(.x(x_79), .z(tmp00_79_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480080(.x(x_80), .z(tmp00_80_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480081(.x(x_81), .z(tmp00_81_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480082(.x(x_82), .z(tmp00_82_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480083(.x(x_83), .z(tmp00_83_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480084(.x(x_84), .z(tmp00_84_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480085(.x(x_85), .z(tmp00_85_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480086(.x(x_86), .z(tmp00_86_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480087(.x(x_87), .z(tmp00_87_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480088(.x(x_88), .z(tmp00_88_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480089(.x(x_89), .z(tmp00_89_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480090(.x(x_90), .z(tmp00_90_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480091(.x(x_91), .z(tmp00_91_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480092(.x(x_92), .z(tmp00_92_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480093(.x(x_93), .z(tmp00_93_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480094(.x(x_94), .z(tmp00_94_48));
	booth_0010 #(.WIDTH(WIDTH)) mul00480095(.x(x_95), .z(tmp00_95_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480096(.x(x_96), .z(tmp00_96_48));
	booth_0012 #(.WIDTH(WIDTH)) mul00480097(.x(x_97), .z(tmp00_97_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480098(.x(x_98), .z(tmp00_98_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480099(.x(x_99), .z(tmp00_99_48));
	booth_0010 #(.WIDTH(WIDTH)) mul00480100(.x(x_100), .z(tmp00_100_48));
	booth__006 #(.WIDTH(WIDTH)) mul00480101(.x(x_101), .z(tmp00_101_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480102(.x(x_102), .z(tmp00_102_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480103(.x(x_103), .z(tmp00_103_48));
	booth__006 #(.WIDTH(WIDTH)) mul00480104(.x(x_104), .z(tmp00_104_48));
	booth__012 #(.WIDTH(WIDTH)) mul00480105(.x(x_105), .z(tmp00_105_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480106(.x(x_106), .z(tmp00_106_48));
	booth_0012 #(.WIDTH(WIDTH)) mul00480107(.x(x_107), .z(tmp00_107_48));
	booth__002 #(.WIDTH(WIDTH)) mul00480108(.x(x_108), .z(tmp00_108_48));
	booth__002 #(.WIDTH(WIDTH)) mul00480109(.x(x_109), .z(tmp00_109_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480110(.x(x_110), .z(tmp00_110_48));
	booth_0006 #(.WIDTH(WIDTH)) mul00480111(.x(x_111), .z(tmp00_111_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480112(.x(x_112), .z(tmp00_112_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480113(.x(x_113), .z(tmp00_113_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480114(.x(x_114), .z(tmp00_114_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480115(.x(x_115), .z(tmp00_115_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480116(.x(x_116), .z(tmp00_116_48));
	booth__002 #(.WIDTH(WIDTH)) mul00480117(.x(x_117), .z(tmp00_117_48));
	booth__004 #(.WIDTH(WIDTH)) mul00480118(.x(x_118), .z(tmp00_118_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480119(.x(x_119), .z(tmp00_119_48));
	booth_0010 #(.WIDTH(WIDTH)) mul00480120(.x(x_120), .z(tmp00_120_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480121(.x(x_121), .z(tmp00_121_48));
	booth_0008 #(.WIDTH(WIDTH)) mul00480122(.x(x_122), .z(tmp00_122_48));
	booth__008 #(.WIDTH(WIDTH)) mul00480123(.x(x_123), .z(tmp00_123_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480124(.x(x_124), .z(tmp00_124_48));
	booth_0000 #(.WIDTH(WIDTH)) mul00480125(.x(x_125), .z(tmp00_125_48));
	booth_0004 #(.WIDTH(WIDTH)) mul00480126(.x(x_126), .z(tmp00_126_48));
	booth__010 #(.WIDTH(WIDTH)) mul00480127(.x(x_127), .z(tmp00_127_48));
	booth__006 #(.WIDTH(WIDTH)) mul00490000(.x(x_0), .z(tmp00_0_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490001(.x(x_1), .z(tmp00_1_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490002(.x(x_2), .z(tmp00_2_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490003(.x(x_3), .z(tmp00_3_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490004(.x(x_4), .z(tmp00_4_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490005(.x(x_5), .z(tmp00_5_49));
	booth__002 #(.WIDTH(WIDTH)) mul00490006(.x(x_6), .z(tmp00_6_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490007(.x(x_7), .z(tmp00_7_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490008(.x(x_8), .z(tmp00_8_49));
	booth_0006 #(.WIDTH(WIDTH)) mul00490009(.x(x_9), .z(tmp00_9_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490010(.x(x_10), .z(tmp00_10_49));
	booth_0006 #(.WIDTH(WIDTH)) mul00490011(.x(x_11), .z(tmp00_11_49));
	booth__006 #(.WIDTH(WIDTH)) mul00490012(.x(x_12), .z(tmp00_12_49));
	booth__010 #(.WIDTH(WIDTH)) mul00490013(.x(x_13), .z(tmp00_13_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490014(.x(x_14), .z(tmp00_14_49));
	booth__002 #(.WIDTH(WIDTH)) mul00490015(.x(x_15), .z(tmp00_15_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490016(.x(x_16), .z(tmp00_16_49));
	booth_0006 #(.WIDTH(WIDTH)) mul00490017(.x(x_17), .z(tmp00_17_49));
	booth__010 #(.WIDTH(WIDTH)) mul00490018(.x(x_18), .z(tmp00_18_49));
	booth__006 #(.WIDTH(WIDTH)) mul00490019(.x(x_19), .z(tmp00_19_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490020(.x(x_20), .z(tmp00_20_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490021(.x(x_21), .z(tmp00_21_49));
	booth_0010 #(.WIDTH(WIDTH)) mul00490022(.x(x_22), .z(tmp00_22_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490023(.x(x_23), .z(tmp00_23_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490024(.x(x_24), .z(tmp00_24_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490025(.x(x_25), .z(tmp00_25_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490026(.x(x_26), .z(tmp00_26_49));
	booth_0010 #(.WIDTH(WIDTH)) mul00490027(.x(x_27), .z(tmp00_27_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490028(.x(x_28), .z(tmp00_28_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490029(.x(x_29), .z(tmp00_29_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490030(.x(x_30), .z(tmp00_30_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490031(.x(x_31), .z(tmp00_31_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490032(.x(x_32), .z(tmp00_32_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490033(.x(x_33), .z(tmp00_33_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490034(.x(x_34), .z(tmp00_34_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490035(.x(x_35), .z(tmp00_35_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490036(.x(x_36), .z(tmp00_36_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490037(.x(x_37), .z(tmp00_37_49));
	booth__006 #(.WIDTH(WIDTH)) mul00490038(.x(x_38), .z(tmp00_38_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490039(.x(x_39), .z(tmp00_39_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490040(.x(x_40), .z(tmp00_40_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490041(.x(x_41), .z(tmp00_41_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490042(.x(x_42), .z(tmp00_42_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490043(.x(x_43), .z(tmp00_43_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490044(.x(x_44), .z(tmp00_44_49));
	booth_0002 #(.WIDTH(WIDTH)) mul00490045(.x(x_45), .z(tmp00_45_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490046(.x(x_46), .z(tmp00_46_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490047(.x(x_47), .z(tmp00_47_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490048(.x(x_48), .z(tmp00_48_49));
	booth__010 #(.WIDTH(WIDTH)) mul00490049(.x(x_49), .z(tmp00_49_49));
	booth_0006 #(.WIDTH(WIDTH)) mul00490050(.x(x_50), .z(tmp00_50_49));
	booth__006 #(.WIDTH(WIDTH)) mul00490051(.x(x_51), .z(tmp00_51_49));
	booth_0002 #(.WIDTH(WIDTH)) mul00490052(.x(x_52), .z(tmp00_52_49));
	booth_0010 #(.WIDTH(WIDTH)) mul00490053(.x(x_53), .z(tmp00_53_49));
	booth__010 #(.WIDTH(WIDTH)) mul00490054(.x(x_54), .z(tmp00_54_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490055(.x(x_55), .z(tmp00_55_49));
	booth_0012 #(.WIDTH(WIDTH)) mul00490056(.x(x_56), .z(tmp00_56_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490057(.x(x_57), .z(tmp00_57_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490058(.x(x_58), .z(tmp00_58_49));
	booth__006 #(.WIDTH(WIDTH)) mul00490059(.x(x_59), .z(tmp00_59_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490060(.x(x_60), .z(tmp00_60_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490061(.x(x_61), .z(tmp00_61_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490062(.x(x_62), .z(tmp00_62_49));
	booth__010 #(.WIDTH(WIDTH)) mul00490063(.x(x_63), .z(tmp00_63_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490064(.x(x_64), .z(tmp00_64_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490065(.x(x_65), .z(tmp00_65_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490066(.x(x_66), .z(tmp00_66_49));
	booth__012 #(.WIDTH(WIDTH)) mul00490067(.x(x_67), .z(tmp00_67_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490068(.x(x_68), .z(tmp00_68_49));
	booth_0010 #(.WIDTH(WIDTH)) mul00490069(.x(x_69), .z(tmp00_69_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490070(.x(x_70), .z(tmp00_70_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490071(.x(x_71), .z(tmp00_71_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490072(.x(x_72), .z(tmp00_72_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490073(.x(x_73), .z(tmp00_73_49));
	booth__010 #(.WIDTH(WIDTH)) mul00490074(.x(x_74), .z(tmp00_74_49));
	booth_0006 #(.WIDTH(WIDTH)) mul00490075(.x(x_75), .z(tmp00_75_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490076(.x(x_76), .z(tmp00_76_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490077(.x(x_77), .z(tmp00_77_49));
	booth_0012 #(.WIDTH(WIDTH)) mul00490078(.x(x_78), .z(tmp00_78_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490079(.x(x_79), .z(tmp00_79_49));
	booth_0010 #(.WIDTH(WIDTH)) mul00490080(.x(x_80), .z(tmp00_80_49));
	booth_0010 #(.WIDTH(WIDTH)) mul00490081(.x(x_81), .z(tmp00_81_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490082(.x(x_82), .z(tmp00_82_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490083(.x(x_83), .z(tmp00_83_49));
	booth_0010 #(.WIDTH(WIDTH)) mul00490084(.x(x_84), .z(tmp00_84_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490085(.x(x_85), .z(tmp00_85_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490086(.x(x_86), .z(tmp00_86_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490087(.x(x_87), .z(tmp00_87_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490088(.x(x_88), .z(tmp00_88_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490089(.x(x_89), .z(tmp00_89_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490090(.x(x_90), .z(tmp00_90_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490091(.x(x_91), .z(tmp00_91_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490092(.x(x_92), .z(tmp00_92_49));
	booth_0012 #(.WIDTH(WIDTH)) mul00490093(.x(x_93), .z(tmp00_93_49));
	booth__002 #(.WIDTH(WIDTH)) mul00490094(.x(x_94), .z(tmp00_94_49));
	booth__002 #(.WIDTH(WIDTH)) mul00490095(.x(x_95), .z(tmp00_95_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490096(.x(x_96), .z(tmp00_96_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490097(.x(x_97), .z(tmp00_97_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490098(.x(x_98), .z(tmp00_98_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490099(.x(x_99), .z(tmp00_99_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490100(.x(x_100), .z(tmp00_100_49));
	booth__008 #(.WIDTH(WIDTH)) mul00490101(.x(x_101), .z(tmp00_101_49));
	booth_0006 #(.WIDTH(WIDTH)) mul00490102(.x(x_102), .z(tmp00_102_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490103(.x(x_103), .z(tmp00_103_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490104(.x(x_104), .z(tmp00_104_49));
	booth__012 #(.WIDTH(WIDTH)) mul00490105(.x(x_105), .z(tmp00_105_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490106(.x(x_106), .z(tmp00_106_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490107(.x(x_107), .z(tmp00_107_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490108(.x(x_108), .z(tmp00_108_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490109(.x(x_109), .z(tmp00_109_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490110(.x(x_110), .z(tmp00_110_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490111(.x(x_111), .z(tmp00_111_49));
	booth__010 #(.WIDTH(WIDTH)) mul00490112(.x(x_112), .z(tmp00_112_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490113(.x(x_113), .z(tmp00_113_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490114(.x(x_114), .z(tmp00_114_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490115(.x(x_115), .z(tmp00_115_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490116(.x(x_116), .z(tmp00_116_49));
	booth__004 #(.WIDTH(WIDTH)) mul00490117(.x(x_117), .z(tmp00_117_49));
	booth__002 #(.WIDTH(WIDTH)) mul00490118(.x(x_118), .z(tmp00_118_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490119(.x(x_119), .z(tmp00_119_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490120(.x(x_120), .z(tmp00_120_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490121(.x(x_121), .z(tmp00_121_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490122(.x(x_122), .z(tmp00_122_49));
	booth__010 #(.WIDTH(WIDTH)) mul00490123(.x(x_123), .z(tmp00_123_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490124(.x(x_124), .z(tmp00_124_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00490125(.x(x_125), .z(tmp00_125_49));
	booth_0008 #(.WIDTH(WIDTH)) mul00490126(.x(x_126), .z(tmp00_126_49));
	booth_0004 #(.WIDTH(WIDTH)) mul00490127(.x(x_127), .z(tmp00_127_49));
	booth_0000 #(.WIDTH(WIDTH)) mul00500000(.x(x_0), .z(tmp00_0_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500001(.x(x_1), .z(tmp00_1_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500002(.x(x_2), .z(tmp00_2_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500003(.x(x_3), .z(tmp00_3_50));
	booth_0012 #(.WIDTH(WIDTH)) mul00500004(.x(x_4), .z(tmp00_4_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500005(.x(x_5), .z(tmp00_5_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500006(.x(x_6), .z(tmp00_6_50));
	booth_0006 #(.WIDTH(WIDTH)) mul00500007(.x(x_7), .z(tmp00_7_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500008(.x(x_8), .z(tmp00_8_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500009(.x(x_9), .z(tmp00_9_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500010(.x(x_10), .z(tmp00_10_50));
	booth_0010 #(.WIDTH(WIDTH)) mul00500011(.x(x_11), .z(tmp00_11_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500012(.x(x_12), .z(tmp00_12_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500013(.x(x_13), .z(tmp00_13_50));
	booth__012 #(.WIDTH(WIDTH)) mul00500014(.x(x_14), .z(tmp00_14_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500015(.x(x_15), .z(tmp00_15_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500016(.x(x_16), .z(tmp00_16_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500017(.x(x_17), .z(tmp00_17_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500018(.x(x_18), .z(tmp00_18_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500019(.x(x_19), .z(tmp00_19_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500020(.x(x_20), .z(tmp00_20_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500021(.x(x_21), .z(tmp00_21_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500022(.x(x_22), .z(tmp00_22_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500023(.x(x_23), .z(tmp00_23_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500024(.x(x_24), .z(tmp00_24_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500025(.x(x_25), .z(tmp00_25_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500026(.x(x_26), .z(tmp00_26_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500027(.x(x_27), .z(tmp00_27_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500028(.x(x_28), .z(tmp00_28_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500029(.x(x_29), .z(tmp00_29_50));
	booth_0012 #(.WIDTH(WIDTH)) mul00500030(.x(x_30), .z(tmp00_30_50));
	booth__002 #(.WIDTH(WIDTH)) mul00500031(.x(x_31), .z(tmp00_31_50));
	booth__002 #(.WIDTH(WIDTH)) mul00500032(.x(x_32), .z(tmp00_32_50));
	booth_0002 #(.WIDTH(WIDTH)) mul00500033(.x(x_33), .z(tmp00_33_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500034(.x(x_34), .z(tmp00_34_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500035(.x(x_35), .z(tmp00_35_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500036(.x(x_36), .z(tmp00_36_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500037(.x(x_37), .z(tmp00_37_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500038(.x(x_38), .z(tmp00_38_50));
	booth__002 #(.WIDTH(WIDTH)) mul00500039(.x(x_39), .z(tmp00_39_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500040(.x(x_40), .z(tmp00_40_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500041(.x(x_41), .z(tmp00_41_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500042(.x(x_42), .z(tmp00_42_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500043(.x(x_43), .z(tmp00_43_50));
	booth_0010 #(.WIDTH(WIDTH)) mul00500044(.x(x_44), .z(tmp00_44_50));
	booth_0010 #(.WIDTH(WIDTH)) mul00500045(.x(x_45), .z(tmp00_45_50));
	booth__012 #(.WIDTH(WIDTH)) mul00500046(.x(x_46), .z(tmp00_46_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500047(.x(x_47), .z(tmp00_47_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500048(.x(x_48), .z(tmp00_48_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500049(.x(x_49), .z(tmp00_49_50));
	booth__010 #(.WIDTH(WIDTH)) mul00500050(.x(x_50), .z(tmp00_50_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500051(.x(x_51), .z(tmp00_51_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500052(.x(x_52), .z(tmp00_52_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500053(.x(x_53), .z(tmp00_53_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500054(.x(x_54), .z(tmp00_54_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500055(.x(x_55), .z(tmp00_55_50));
	booth__002 #(.WIDTH(WIDTH)) mul00500056(.x(x_56), .z(tmp00_56_50));
	booth_0012 #(.WIDTH(WIDTH)) mul00500057(.x(x_57), .z(tmp00_57_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500058(.x(x_58), .z(tmp00_58_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500059(.x(x_59), .z(tmp00_59_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500060(.x(x_60), .z(tmp00_60_50));
	booth_0006 #(.WIDTH(WIDTH)) mul00500061(.x(x_61), .z(tmp00_61_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500062(.x(x_62), .z(tmp00_62_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500063(.x(x_63), .z(tmp00_63_50));
	booth_0002 #(.WIDTH(WIDTH)) mul00500064(.x(x_64), .z(tmp00_64_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500065(.x(x_65), .z(tmp00_65_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500066(.x(x_66), .z(tmp00_66_50));
	booth_0006 #(.WIDTH(WIDTH)) mul00500067(.x(x_67), .z(tmp00_67_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500068(.x(x_68), .z(tmp00_68_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500069(.x(x_69), .z(tmp00_69_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500070(.x(x_70), .z(tmp00_70_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500071(.x(x_71), .z(tmp00_71_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500072(.x(x_72), .z(tmp00_72_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500073(.x(x_73), .z(tmp00_73_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500074(.x(x_74), .z(tmp00_74_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500075(.x(x_75), .z(tmp00_75_50));
	booth_0012 #(.WIDTH(WIDTH)) mul00500076(.x(x_76), .z(tmp00_76_50));
	booth_0010 #(.WIDTH(WIDTH)) mul00500077(.x(x_77), .z(tmp00_77_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500078(.x(x_78), .z(tmp00_78_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500079(.x(x_79), .z(tmp00_79_50));
	booth__002 #(.WIDTH(WIDTH)) mul00500080(.x(x_80), .z(tmp00_80_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500081(.x(x_81), .z(tmp00_81_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500082(.x(x_82), .z(tmp00_82_50));
	booth_0002 #(.WIDTH(WIDTH)) mul00500083(.x(x_83), .z(tmp00_83_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500084(.x(x_84), .z(tmp00_84_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500085(.x(x_85), .z(tmp00_85_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500086(.x(x_86), .z(tmp00_86_50));
	booth_0002 #(.WIDTH(WIDTH)) mul00500087(.x(x_87), .z(tmp00_87_50));
	booth_0002 #(.WIDTH(WIDTH)) mul00500088(.x(x_88), .z(tmp00_88_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500089(.x(x_89), .z(tmp00_89_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500090(.x(x_90), .z(tmp00_90_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500091(.x(x_91), .z(tmp00_91_50));
	booth_0002 #(.WIDTH(WIDTH)) mul00500092(.x(x_92), .z(tmp00_92_50));
	booth__002 #(.WIDTH(WIDTH)) mul00500093(.x(x_93), .z(tmp00_93_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500094(.x(x_94), .z(tmp00_94_50));
	booth_0006 #(.WIDTH(WIDTH)) mul00500095(.x(x_95), .z(tmp00_95_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500096(.x(x_96), .z(tmp00_96_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500097(.x(x_97), .z(tmp00_97_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500098(.x(x_98), .z(tmp00_98_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500099(.x(x_99), .z(tmp00_99_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500100(.x(x_100), .z(tmp00_100_50));
	booth_0006 #(.WIDTH(WIDTH)) mul00500101(.x(x_101), .z(tmp00_101_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500102(.x(x_102), .z(tmp00_102_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500103(.x(x_103), .z(tmp00_103_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500104(.x(x_104), .z(tmp00_104_50));
	booth_0010 #(.WIDTH(WIDTH)) mul00500105(.x(x_105), .z(tmp00_105_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500106(.x(x_106), .z(tmp00_106_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500107(.x(x_107), .z(tmp00_107_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500108(.x(x_108), .z(tmp00_108_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500109(.x(x_109), .z(tmp00_109_50));
	booth__006 #(.WIDTH(WIDTH)) mul00500110(.x(x_110), .z(tmp00_110_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500111(.x(x_111), .z(tmp00_111_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500112(.x(x_112), .z(tmp00_112_50));
	booth__004 #(.WIDTH(WIDTH)) mul00500113(.x(x_113), .z(tmp00_113_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500114(.x(x_114), .z(tmp00_114_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500115(.x(x_115), .z(tmp00_115_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500116(.x(x_116), .z(tmp00_116_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500117(.x(x_117), .z(tmp00_117_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500118(.x(x_118), .z(tmp00_118_50));
	booth_0006 #(.WIDTH(WIDTH)) mul00500119(.x(x_119), .z(tmp00_119_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500120(.x(x_120), .z(tmp00_120_50));
	booth_0008 #(.WIDTH(WIDTH)) mul00500121(.x(x_121), .z(tmp00_121_50));
	booth_0002 #(.WIDTH(WIDTH)) mul00500122(.x(x_122), .z(tmp00_122_50));
	booth_0010 #(.WIDTH(WIDTH)) mul00500123(.x(x_123), .z(tmp00_123_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500124(.x(x_124), .z(tmp00_124_50));
	booth_0000 #(.WIDTH(WIDTH)) mul00500125(.x(x_125), .z(tmp00_125_50));
	booth__008 #(.WIDTH(WIDTH)) mul00500126(.x(x_126), .z(tmp00_126_50));
	booth_0004 #(.WIDTH(WIDTH)) mul00500127(.x(x_127), .z(tmp00_127_50));
	booth_0010 #(.WIDTH(WIDTH)) mul00510000(.x(x_0), .z(tmp00_0_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510001(.x(x_1), .z(tmp00_1_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510002(.x(x_2), .z(tmp00_2_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510003(.x(x_3), .z(tmp00_3_51));
	booth__012 #(.WIDTH(WIDTH)) mul00510004(.x(x_4), .z(tmp00_4_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510005(.x(x_5), .z(tmp00_5_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510006(.x(x_6), .z(tmp00_6_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510007(.x(x_7), .z(tmp00_7_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510008(.x(x_8), .z(tmp00_8_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510009(.x(x_9), .z(tmp00_9_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510010(.x(x_10), .z(tmp00_10_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510011(.x(x_11), .z(tmp00_11_51));
	booth__006 #(.WIDTH(WIDTH)) mul00510012(.x(x_12), .z(tmp00_12_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510013(.x(x_13), .z(tmp00_13_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510014(.x(x_14), .z(tmp00_14_51));
	booth__002 #(.WIDTH(WIDTH)) mul00510015(.x(x_15), .z(tmp00_15_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510016(.x(x_16), .z(tmp00_16_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510017(.x(x_17), .z(tmp00_17_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510018(.x(x_18), .z(tmp00_18_51));
	booth_0012 #(.WIDTH(WIDTH)) mul00510019(.x(x_19), .z(tmp00_19_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510020(.x(x_20), .z(tmp00_20_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510021(.x(x_21), .z(tmp00_21_51));
	booth_0006 #(.WIDTH(WIDTH)) mul00510022(.x(x_22), .z(tmp00_22_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510023(.x(x_23), .z(tmp00_23_51));
	booth_0002 #(.WIDTH(WIDTH)) mul00510024(.x(x_24), .z(tmp00_24_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510025(.x(x_25), .z(tmp00_25_51));
	booth_0010 #(.WIDTH(WIDTH)) mul00510026(.x(x_26), .z(tmp00_26_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510027(.x(x_27), .z(tmp00_27_51));
	booth_0016 #(.WIDTH(WIDTH)) mul00510028(.x(x_28), .z(tmp00_28_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510029(.x(x_29), .z(tmp00_29_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510030(.x(x_30), .z(tmp00_30_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510031(.x(x_31), .z(tmp00_31_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510032(.x(x_32), .z(tmp00_32_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510033(.x(x_33), .z(tmp00_33_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510034(.x(x_34), .z(tmp00_34_51));
	booth_0012 #(.WIDTH(WIDTH)) mul00510035(.x(x_35), .z(tmp00_35_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510036(.x(x_36), .z(tmp00_36_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510037(.x(x_37), .z(tmp00_37_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510038(.x(x_38), .z(tmp00_38_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510039(.x(x_39), .z(tmp00_39_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510040(.x(x_40), .z(tmp00_40_51));
	booth__010 #(.WIDTH(WIDTH)) mul00510041(.x(x_41), .z(tmp00_41_51));
	booth_0014 #(.WIDTH(WIDTH)) mul00510042(.x(x_42), .z(tmp00_42_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510043(.x(x_43), .z(tmp00_43_51));
	booth_0010 #(.WIDTH(WIDTH)) mul00510044(.x(x_44), .z(tmp00_44_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510045(.x(x_45), .z(tmp00_45_51));
	booth_0016 #(.WIDTH(WIDTH)) mul00510046(.x(x_46), .z(tmp00_46_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510047(.x(x_47), .z(tmp00_47_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510048(.x(x_48), .z(tmp00_48_51));
	booth_0016 #(.WIDTH(WIDTH)) mul00510049(.x(x_49), .z(tmp00_49_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510050(.x(x_50), .z(tmp00_50_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510051(.x(x_51), .z(tmp00_51_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510052(.x(x_52), .z(tmp00_52_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510053(.x(x_53), .z(tmp00_53_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510054(.x(x_54), .z(tmp00_54_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510055(.x(x_55), .z(tmp00_55_51));
	booth_0012 #(.WIDTH(WIDTH)) mul00510056(.x(x_56), .z(tmp00_56_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510057(.x(x_57), .z(tmp00_57_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510058(.x(x_58), .z(tmp00_58_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510059(.x(x_59), .z(tmp00_59_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510060(.x(x_60), .z(tmp00_60_51));
	booth_0012 #(.WIDTH(WIDTH)) mul00510061(.x(x_61), .z(tmp00_61_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510062(.x(x_62), .z(tmp00_62_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510063(.x(x_63), .z(tmp00_63_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510064(.x(x_64), .z(tmp00_64_51));
	booth__006 #(.WIDTH(WIDTH)) mul00510065(.x(x_65), .z(tmp00_65_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510066(.x(x_66), .z(tmp00_66_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510067(.x(x_67), .z(tmp00_67_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510068(.x(x_68), .z(tmp00_68_51));
	booth__012 #(.WIDTH(WIDTH)) mul00510069(.x(x_69), .z(tmp00_69_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510070(.x(x_70), .z(tmp00_70_51));
	booth_0012 #(.WIDTH(WIDTH)) mul00510071(.x(x_71), .z(tmp00_71_51));
	booth__012 #(.WIDTH(WIDTH)) mul00510072(.x(x_72), .z(tmp00_72_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510073(.x(x_73), .z(tmp00_73_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510074(.x(x_74), .z(tmp00_74_51));
	booth_0014 #(.WIDTH(WIDTH)) mul00510075(.x(x_75), .z(tmp00_75_51));
	booth__002 #(.WIDTH(WIDTH)) mul00510076(.x(x_76), .z(tmp00_76_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510077(.x(x_77), .z(tmp00_77_51));
	booth_0002 #(.WIDTH(WIDTH)) mul00510078(.x(x_78), .z(tmp00_78_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510079(.x(x_79), .z(tmp00_79_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510080(.x(x_80), .z(tmp00_80_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510081(.x(x_81), .z(tmp00_81_51));
	booth__016 #(.WIDTH(WIDTH)) mul00510082(.x(x_82), .z(tmp00_82_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510083(.x(x_83), .z(tmp00_83_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510084(.x(x_84), .z(tmp00_84_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510085(.x(x_85), .z(tmp00_85_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510086(.x(x_86), .z(tmp00_86_51));
	booth_0012 #(.WIDTH(WIDTH)) mul00510087(.x(x_87), .z(tmp00_87_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510088(.x(x_88), .z(tmp00_88_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510089(.x(x_89), .z(tmp00_89_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510090(.x(x_90), .z(tmp00_90_51));
	booth_0002 #(.WIDTH(WIDTH)) mul00510091(.x(x_91), .z(tmp00_91_51));
	booth_0006 #(.WIDTH(WIDTH)) mul00510092(.x(x_92), .z(tmp00_92_51));
	booth_0012 #(.WIDTH(WIDTH)) mul00510093(.x(x_93), .z(tmp00_93_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510094(.x(x_94), .z(tmp00_94_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510095(.x(x_95), .z(tmp00_95_51));
	booth_0006 #(.WIDTH(WIDTH)) mul00510096(.x(x_96), .z(tmp00_96_51));
	booth__006 #(.WIDTH(WIDTH)) mul00510097(.x(x_97), .z(tmp00_97_51));
	booth__014 #(.WIDTH(WIDTH)) mul00510098(.x(x_98), .z(tmp00_98_51));
	booth_0006 #(.WIDTH(WIDTH)) mul00510099(.x(x_99), .z(tmp00_99_51));
	booth_0016 #(.WIDTH(WIDTH)) mul00510100(.x(x_100), .z(tmp00_100_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510101(.x(x_101), .z(tmp00_101_51));
	booth_0012 #(.WIDTH(WIDTH)) mul00510102(.x(x_102), .z(tmp00_102_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510103(.x(x_103), .z(tmp00_103_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510104(.x(x_104), .z(tmp00_104_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510105(.x(x_105), .z(tmp00_105_51));
	booth_0010 #(.WIDTH(WIDTH)) mul00510106(.x(x_106), .z(tmp00_106_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510107(.x(x_107), .z(tmp00_107_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510108(.x(x_108), .z(tmp00_108_51));
	booth_0008 #(.WIDTH(WIDTH)) mul00510109(.x(x_109), .z(tmp00_109_51));
	booth__002 #(.WIDTH(WIDTH)) mul00510110(.x(x_110), .z(tmp00_110_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510111(.x(x_111), .z(tmp00_111_51));
	booth_0006 #(.WIDTH(WIDTH)) mul00510112(.x(x_112), .z(tmp00_112_51));
	booth__012 #(.WIDTH(WIDTH)) mul00510113(.x(x_113), .z(tmp00_113_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510114(.x(x_114), .z(tmp00_114_51));
	booth__016 #(.WIDTH(WIDTH)) mul00510115(.x(x_115), .z(tmp00_115_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510116(.x(x_116), .z(tmp00_116_51));
	booth_0006 #(.WIDTH(WIDTH)) mul00510117(.x(x_117), .z(tmp00_117_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510118(.x(x_118), .z(tmp00_118_51));
	booth__004 #(.WIDTH(WIDTH)) mul00510119(.x(x_119), .z(tmp00_119_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510120(.x(x_120), .z(tmp00_120_51));
	booth__002 #(.WIDTH(WIDTH)) mul00510121(.x(x_121), .z(tmp00_121_51));
	booth__008 #(.WIDTH(WIDTH)) mul00510122(.x(x_122), .z(tmp00_122_51));
	booth_0000 #(.WIDTH(WIDTH)) mul00510123(.x(x_123), .z(tmp00_123_51));
	booth_0016 #(.WIDTH(WIDTH)) mul00510124(.x(x_124), .z(tmp00_124_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510125(.x(x_125), .z(tmp00_125_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00510126(.x(x_126), .z(tmp00_126_51));
	booth_0014 #(.WIDTH(WIDTH)) mul00510127(.x(x_127), .z(tmp00_127_51));
	booth_0004 #(.WIDTH(WIDTH)) mul00520000(.x(x_0), .z(tmp00_0_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520001(.x(x_1), .z(tmp00_1_52));
	booth_0006 #(.WIDTH(WIDTH)) mul00520002(.x(x_2), .z(tmp00_2_52));
	booth_0006 #(.WIDTH(WIDTH)) mul00520003(.x(x_3), .z(tmp00_3_52));
	booth__004 #(.WIDTH(WIDTH)) mul00520004(.x(x_4), .z(tmp00_4_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520005(.x(x_5), .z(tmp00_5_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520006(.x(x_6), .z(tmp00_6_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520007(.x(x_7), .z(tmp00_7_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520008(.x(x_8), .z(tmp00_8_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520009(.x(x_9), .z(tmp00_9_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520010(.x(x_10), .z(tmp00_10_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520011(.x(x_11), .z(tmp00_11_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520012(.x(x_12), .z(tmp00_12_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520013(.x(x_13), .z(tmp00_13_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520014(.x(x_14), .z(tmp00_14_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520015(.x(x_15), .z(tmp00_15_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520016(.x(x_16), .z(tmp00_16_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520017(.x(x_17), .z(tmp00_17_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520018(.x(x_18), .z(tmp00_18_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520019(.x(x_19), .z(tmp00_19_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520020(.x(x_20), .z(tmp00_20_52));
	booth_0010 #(.WIDTH(WIDTH)) mul00520021(.x(x_21), .z(tmp00_21_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520022(.x(x_22), .z(tmp00_22_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520023(.x(x_23), .z(tmp00_23_52));
	booth_0006 #(.WIDTH(WIDTH)) mul00520024(.x(x_24), .z(tmp00_24_52));
	booth__004 #(.WIDTH(WIDTH)) mul00520025(.x(x_25), .z(tmp00_25_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520026(.x(x_26), .z(tmp00_26_52));
	booth__010 #(.WIDTH(WIDTH)) mul00520027(.x(x_27), .z(tmp00_27_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520028(.x(x_28), .z(tmp00_28_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520029(.x(x_29), .z(tmp00_29_52));
	booth_0012 #(.WIDTH(WIDTH)) mul00520030(.x(x_30), .z(tmp00_30_52));
	booth_0002 #(.WIDTH(WIDTH)) mul00520031(.x(x_31), .z(tmp00_31_52));
	booth__004 #(.WIDTH(WIDTH)) mul00520032(.x(x_32), .z(tmp00_32_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520033(.x(x_33), .z(tmp00_33_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520034(.x(x_34), .z(tmp00_34_52));
	booth_0012 #(.WIDTH(WIDTH)) mul00520035(.x(x_35), .z(tmp00_35_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520036(.x(x_36), .z(tmp00_36_52));
	booth__004 #(.WIDTH(WIDTH)) mul00520037(.x(x_37), .z(tmp00_37_52));
	booth__002 #(.WIDTH(WIDTH)) mul00520038(.x(x_38), .z(tmp00_38_52));
	booth_0012 #(.WIDTH(WIDTH)) mul00520039(.x(x_39), .z(tmp00_39_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520040(.x(x_40), .z(tmp00_40_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520041(.x(x_41), .z(tmp00_41_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520042(.x(x_42), .z(tmp00_42_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520043(.x(x_43), .z(tmp00_43_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520044(.x(x_44), .z(tmp00_44_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520045(.x(x_45), .z(tmp00_45_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520046(.x(x_46), .z(tmp00_46_52));
	booth_0010 #(.WIDTH(WIDTH)) mul00520047(.x(x_47), .z(tmp00_47_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520048(.x(x_48), .z(tmp00_48_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520049(.x(x_49), .z(tmp00_49_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520050(.x(x_50), .z(tmp00_50_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520051(.x(x_51), .z(tmp00_51_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520052(.x(x_52), .z(tmp00_52_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520053(.x(x_53), .z(tmp00_53_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520054(.x(x_54), .z(tmp00_54_52));
	booth__010 #(.WIDTH(WIDTH)) mul00520055(.x(x_55), .z(tmp00_55_52));
	booth__006 #(.WIDTH(WIDTH)) mul00520056(.x(x_56), .z(tmp00_56_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520057(.x(x_57), .z(tmp00_57_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520058(.x(x_58), .z(tmp00_58_52));
	booth__010 #(.WIDTH(WIDTH)) mul00520059(.x(x_59), .z(tmp00_59_52));
	booth__006 #(.WIDTH(WIDTH)) mul00520060(.x(x_60), .z(tmp00_60_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520061(.x(x_61), .z(tmp00_61_52));
	booth_0002 #(.WIDTH(WIDTH)) mul00520062(.x(x_62), .z(tmp00_62_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520063(.x(x_63), .z(tmp00_63_52));
	booth__010 #(.WIDTH(WIDTH)) mul00520064(.x(x_64), .z(tmp00_64_52));
	booth__002 #(.WIDTH(WIDTH)) mul00520065(.x(x_65), .z(tmp00_65_52));
	booth_0012 #(.WIDTH(WIDTH)) mul00520066(.x(x_66), .z(tmp00_66_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520067(.x(x_67), .z(tmp00_67_52));
	booth__006 #(.WIDTH(WIDTH)) mul00520068(.x(x_68), .z(tmp00_68_52));
	booth__004 #(.WIDTH(WIDTH)) mul00520069(.x(x_69), .z(tmp00_69_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520070(.x(x_70), .z(tmp00_70_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520071(.x(x_71), .z(tmp00_71_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520072(.x(x_72), .z(tmp00_72_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520073(.x(x_73), .z(tmp00_73_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520074(.x(x_74), .z(tmp00_74_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520075(.x(x_75), .z(tmp00_75_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520076(.x(x_76), .z(tmp00_76_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520077(.x(x_77), .z(tmp00_77_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520078(.x(x_78), .z(tmp00_78_52));
	booth__004 #(.WIDTH(WIDTH)) mul00520079(.x(x_79), .z(tmp00_79_52));
	booth_0002 #(.WIDTH(WIDTH)) mul00520080(.x(x_80), .z(tmp00_80_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520081(.x(x_81), .z(tmp00_81_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520082(.x(x_82), .z(tmp00_82_52));
	booth__012 #(.WIDTH(WIDTH)) mul00520083(.x(x_83), .z(tmp00_83_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520084(.x(x_84), .z(tmp00_84_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520085(.x(x_85), .z(tmp00_85_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520086(.x(x_86), .z(tmp00_86_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520087(.x(x_87), .z(tmp00_87_52));
	booth__004 #(.WIDTH(WIDTH)) mul00520088(.x(x_88), .z(tmp00_88_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520089(.x(x_89), .z(tmp00_89_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520090(.x(x_90), .z(tmp00_90_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520091(.x(x_91), .z(tmp00_91_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520092(.x(x_92), .z(tmp00_92_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520093(.x(x_93), .z(tmp00_93_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520094(.x(x_94), .z(tmp00_94_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520095(.x(x_95), .z(tmp00_95_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520096(.x(x_96), .z(tmp00_96_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520097(.x(x_97), .z(tmp00_97_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520098(.x(x_98), .z(tmp00_98_52));
	booth__006 #(.WIDTH(WIDTH)) mul00520099(.x(x_99), .z(tmp00_99_52));
	booth_0012 #(.WIDTH(WIDTH)) mul00520100(.x(x_100), .z(tmp00_100_52));
	booth_0010 #(.WIDTH(WIDTH)) mul00520101(.x(x_101), .z(tmp00_101_52));
	booth_0006 #(.WIDTH(WIDTH)) mul00520102(.x(x_102), .z(tmp00_102_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520103(.x(x_103), .z(tmp00_103_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520104(.x(x_104), .z(tmp00_104_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520105(.x(x_105), .z(tmp00_105_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520106(.x(x_106), .z(tmp00_106_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520107(.x(x_107), .z(tmp00_107_52));
	booth__002 #(.WIDTH(WIDTH)) mul00520108(.x(x_108), .z(tmp00_108_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520109(.x(x_109), .z(tmp00_109_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520110(.x(x_110), .z(tmp00_110_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520111(.x(x_111), .z(tmp00_111_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520112(.x(x_112), .z(tmp00_112_52));
	booth__010 #(.WIDTH(WIDTH)) mul00520113(.x(x_113), .z(tmp00_113_52));
	booth__002 #(.WIDTH(WIDTH)) mul00520114(.x(x_114), .z(tmp00_114_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520115(.x(x_115), .z(tmp00_115_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520116(.x(x_116), .z(tmp00_116_52));
	booth__010 #(.WIDTH(WIDTH)) mul00520117(.x(x_117), .z(tmp00_117_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520118(.x(x_118), .z(tmp00_118_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520119(.x(x_119), .z(tmp00_119_52));
	booth__004 #(.WIDTH(WIDTH)) mul00520120(.x(x_120), .z(tmp00_120_52));
	booth__012 #(.WIDTH(WIDTH)) mul00520121(.x(x_121), .z(tmp00_121_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520122(.x(x_122), .z(tmp00_122_52));
	booth_0004 #(.WIDTH(WIDTH)) mul00520123(.x(x_123), .z(tmp00_123_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00520124(.x(x_124), .z(tmp00_124_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520125(.x(x_125), .z(tmp00_125_52));
	booth__008 #(.WIDTH(WIDTH)) mul00520126(.x(x_126), .z(tmp00_126_52));
	booth_0008 #(.WIDTH(WIDTH)) mul00520127(.x(x_127), .z(tmp00_127_52));
	booth_0000 #(.WIDTH(WIDTH)) mul00530000(.x(x_0), .z(tmp00_0_53));
	booth_0006 #(.WIDTH(WIDTH)) mul00530001(.x(x_1), .z(tmp00_1_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530002(.x(x_2), .z(tmp00_2_53));
	booth_0002 #(.WIDTH(WIDTH)) mul00530003(.x(x_3), .z(tmp00_3_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530004(.x(x_4), .z(tmp00_4_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530005(.x(x_5), .z(tmp00_5_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530006(.x(x_6), .z(tmp00_6_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530007(.x(x_7), .z(tmp00_7_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530008(.x(x_8), .z(tmp00_8_53));
	booth__006 #(.WIDTH(WIDTH)) mul00530009(.x(x_9), .z(tmp00_9_53));
	booth__006 #(.WIDTH(WIDTH)) mul00530010(.x(x_10), .z(tmp00_10_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530011(.x(x_11), .z(tmp00_11_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530012(.x(x_12), .z(tmp00_12_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530013(.x(x_13), .z(tmp00_13_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530014(.x(x_14), .z(tmp00_14_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530015(.x(x_15), .z(tmp00_15_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530016(.x(x_16), .z(tmp00_16_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530017(.x(x_17), .z(tmp00_17_53));
	booth__006 #(.WIDTH(WIDTH)) mul00530018(.x(x_18), .z(tmp00_18_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530019(.x(x_19), .z(tmp00_19_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530020(.x(x_20), .z(tmp00_20_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530021(.x(x_21), .z(tmp00_21_53));
	booth_0010 #(.WIDTH(WIDTH)) mul00530022(.x(x_22), .z(tmp00_22_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530023(.x(x_23), .z(tmp00_23_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530024(.x(x_24), .z(tmp00_24_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530025(.x(x_25), .z(tmp00_25_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530026(.x(x_26), .z(tmp00_26_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530027(.x(x_27), .z(tmp00_27_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530028(.x(x_28), .z(tmp00_28_53));
	booth_0010 #(.WIDTH(WIDTH)) mul00530029(.x(x_29), .z(tmp00_29_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530030(.x(x_30), .z(tmp00_30_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530031(.x(x_31), .z(tmp00_31_53));
	booth_0006 #(.WIDTH(WIDTH)) mul00530032(.x(x_32), .z(tmp00_32_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530033(.x(x_33), .z(tmp00_33_53));
	booth__012 #(.WIDTH(WIDTH)) mul00530034(.x(x_34), .z(tmp00_34_53));
	booth_0010 #(.WIDTH(WIDTH)) mul00530035(.x(x_35), .z(tmp00_35_53));
	booth_0012 #(.WIDTH(WIDTH)) mul00530036(.x(x_36), .z(tmp00_36_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530037(.x(x_37), .z(tmp00_37_53));
	booth__002 #(.WIDTH(WIDTH)) mul00530038(.x(x_38), .z(tmp00_38_53));
	booth__006 #(.WIDTH(WIDTH)) mul00530039(.x(x_39), .z(tmp00_39_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530040(.x(x_40), .z(tmp00_40_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530041(.x(x_41), .z(tmp00_41_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530042(.x(x_42), .z(tmp00_42_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530043(.x(x_43), .z(tmp00_43_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530044(.x(x_44), .z(tmp00_44_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530045(.x(x_45), .z(tmp00_45_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530046(.x(x_46), .z(tmp00_46_53));
	booth__002 #(.WIDTH(WIDTH)) mul00530047(.x(x_47), .z(tmp00_47_53));
	booth_0006 #(.WIDTH(WIDTH)) mul00530048(.x(x_48), .z(tmp00_48_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530049(.x(x_49), .z(tmp00_49_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530050(.x(x_50), .z(tmp00_50_53));
	booth__010 #(.WIDTH(WIDTH)) mul00530051(.x(x_51), .z(tmp00_51_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530052(.x(x_52), .z(tmp00_52_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530053(.x(x_53), .z(tmp00_53_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530054(.x(x_54), .z(tmp00_54_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530055(.x(x_55), .z(tmp00_55_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530056(.x(x_56), .z(tmp00_56_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530057(.x(x_57), .z(tmp00_57_53));
	booth__012 #(.WIDTH(WIDTH)) mul00530058(.x(x_58), .z(tmp00_58_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530059(.x(x_59), .z(tmp00_59_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530060(.x(x_60), .z(tmp00_60_53));
	booth_0006 #(.WIDTH(WIDTH)) mul00530061(.x(x_61), .z(tmp00_61_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530062(.x(x_62), .z(tmp00_62_53));
	booth__002 #(.WIDTH(WIDTH)) mul00530063(.x(x_63), .z(tmp00_63_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530064(.x(x_64), .z(tmp00_64_53));
	booth__002 #(.WIDTH(WIDTH)) mul00530065(.x(x_65), .z(tmp00_65_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530066(.x(x_66), .z(tmp00_66_53));
	booth__006 #(.WIDTH(WIDTH)) mul00530067(.x(x_67), .z(tmp00_67_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530068(.x(x_68), .z(tmp00_68_53));
	booth__006 #(.WIDTH(WIDTH)) mul00530069(.x(x_69), .z(tmp00_69_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530070(.x(x_70), .z(tmp00_70_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530071(.x(x_71), .z(tmp00_71_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530072(.x(x_72), .z(tmp00_72_53));
	booth__006 #(.WIDTH(WIDTH)) mul00530073(.x(x_73), .z(tmp00_73_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530074(.x(x_74), .z(tmp00_74_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530075(.x(x_75), .z(tmp00_75_53));
	booth_0002 #(.WIDTH(WIDTH)) mul00530076(.x(x_76), .z(tmp00_76_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530077(.x(x_77), .z(tmp00_77_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530078(.x(x_78), .z(tmp00_78_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530079(.x(x_79), .z(tmp00_79_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530080(.x(x_80), .z(tmp00_80_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530081(.x(x_81), .z(tmp00_81_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530082(.x(x_82), .z(tmp00_82_53));
	booth_0002 #(.WIDTH(WIDTH)) mul00530083(.x(x_83), .z(tmp00_83_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530084(.x(x_84), .z(tmp00_84_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530085(.x(x_85), .z(tmp00_85_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530086(.x(x_86), .z(tmp00_86_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530087(.x(x_87), .z(tmp00_87_53));
	booth__010 #(.WIDTH(WIDTH)) mul00530088(.x(x_88), .z(tmp00_88_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530089(.x(x_89), .z(tmp00_89_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530090(.x(x_90), .z(tmp00_90_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530091(.x(x_91), .z(tmp00_91_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530092(.x(x_92), .z(tmp00_92_53));
	booth_0006 #(.WIDTH(WIDTH)) mul00530093(.x(x_93), .z(tmp00_93_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530094(.x(x_94), .z(tmp00_94_53));
	booth_0010 #(.WIDTH(WIDTH)) mul00530095(.x(x_95), .z(tmp00_95_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530096(.x(x_96), .z(tmp00_96_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530097(.x(x_97), .z(tmp00_97_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530098(.x(x_98), .z(tmp00_98_53));
	booth__010 #(.WIDTH(WIDTH)) mul00530099(.x(x_99), .z(tmp00_99_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530100(.x(x_100), .z(tmp00_100_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530101(.x(x_101), .z(tmp00_101_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530102(.x(x_102), .z(tmp00_102_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530103(.x(x_103), .z(tmp00_103_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530104(.x(x_104), .z(tmp00_104_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530105(.x(x_105), .z(tmp00_105_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530106(.x(x_106), .z(tmp00_106_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530107(.x(x_107), .z(tmp00_107_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530108(.x(x_108), .z(tmp00_108_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530109(.x(x_109), .z(tmp00_109_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530110(.x(x_110), .z(tmp00_110_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530111(.x(x_111), .z(tmp00_111_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530112(.x(x_112), .z(tmp00_112_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530113(.x(x_113), .z(tmp00_113_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530114(.x(x_114), .z(tmp00_114_53));
	booth_0006 #(.WIDTH(WIDTH)) mul00530115(.x(x_115), .z(tmp00_115_53));
	booth__012 #(.WIDTH(WIDTH)) mul00530116(.x(x_116), .z(tmp00_116_53));
	booth_0008 #(.WIDTH(WIDTH)) mul00530117(.x(x_117), .z(tmp00_117_53));
	booth_0002 #(.WIDTH(WIDTH)) mul00530118(.x(x_118), .z(tmp00_118_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530119(.x(x_119), .z(tmp00_119_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530120(.x(x_120), .z(tmp00_120_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530121(.x(x_121), .z(tmp00_121_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530122(.x(x_122), .z(tmp00_122_53));
	booth__004 #(.WIDTH(WIDTH)) mul00530123(.x(x_123), .z(tmp00_123_53));
	booth_0004 #(.WIDTH(WIDTH)) mul00530124(.x(x_124), .z(tmp00_124_53));
	booth__008 #(.WIDTH(WIDTH)) mul00530125(.x(x_125), .z(tmp00_125_53));
	booth_0010 #(.WIDTH(WIDTH)) mul00530126(.x(x_126), .z(tmp00_126_53));
	booth_0000 #(.WIDTH(WIDTH)) mul00530127(.x(x_127), .z(tmp00_127_53));
	booth__008 #(.WIDTH(WIDTH)) mul00540000(.x(x_0), .z(tmp00_0_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540001(.x(x_1), .z(tmp00_1_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540002(.x(x_2), .z(tmp00_2_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540003(.x(x_3), .z(tmp00_3_54));
	booth_0016 #(.WIDTH(WIDTH)) mul00540004(.x(x_4), .z(tmp00_4_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540005(.x(x_5), .z(tmp00_5_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540006(.x(x_6), .z(tmp00_6_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540007(.x(x_7), .z(tmp00_7_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540008(.x(x_8), .z(tmp00_8_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540009(.x(x_9), .z(tmp00_9_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540010(.x(x_10), .z(tmp00_10_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540011(.x(x_11), .z(tmp00_11_54));
	booth_0010 #(.WIDTH(WIDTH)) mul00540012(.x(x_12), .z(tmp00_12_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540013(.x(x_13), .z(tmp00_13_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540014(.x(x_14), .z(tmp00_14_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540015(.x(x_15), .z(tmp00_15_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540016(.x(x_16), .z(tmp00_16_54));
	booth_0012 #(.WIDTH(WIDTH)) mul00540017(.x(x_17), .z(tmp00_17_54));
	booth_0014 #(.WIDTH(WIDTH)) mul00540018(.x(x_18), .z(tmp00_18_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540019(.x(x_19), .z(tmp00_19_54));
	booth_0010 #(.WIDTH(WIDTH)) mul00540020(.x(x_20), .z(tmp00_20_54));
	booth_0006 #(.WIDTH(WIDTH)) mul00540021(.x(x_21), .z(tmp00_21_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540022(.x(x_22), .z(tmp00_22_54));
	booth_0016 #(.WIDTH(WIDTH)) mul00540023(.x(x_23), .z(tmp00_23_54));
	booth_0012 #(.WIDTH(WIDTH)) mul00540024(.x(x_24), .z(tmp00_24_54));
	booth__010 #(.WIDTH(WIDTH)) mul00540025(.x(x_25), .z(tmp00_25_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540026(.x(x_26), .z(tmp00_26_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540027(.x(x_27), .z(tmp00_27_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540028(.x(x_28), .z(tmp00_28_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540029(.x(x_29), .z(tmp00_29_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540030(.x(x_30), .z(tmp00_30_54));
	booth_0002 #(.WIDTH(WIDTH)) mul00540031(.x(x_31), .z(tmp00_31_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540032(.x(x_32), .z(tmp00_32_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540033(.x(x_33), .z(tmp00_33_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540034(.x(x_34), .z(tmp00_34_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540035(.x(x_35), .z(tmp00_35_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540036(.x(x_36), .z(tmp00_36_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540037(.x(x_37), .z(tmp00_37_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540038(.x(x_38), .z(tmp00_38_54));
	booth__002 #(.WIDTH(WIDTH)) mul00540039(.x(x_39), .z(tmp00_39_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540040(.x(x_40), .z(tmp00_40_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540041(.x(x_41), .z(tmp00_41_54));
	booth__016 #(.WIDTH(WIDTH)) mul00540042(.x(x_42), .z(tmp00_42_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540043(.x(x_43), .z(tmp00_43_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540044(.x(x_44), .z(tmp00_44_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540045(.x(x_45), .z(tmp00_45_54));
	booth_0010 #(.WIDTH(WIDTH)) mul00540046(.x(x_46), .z(tmp00_46_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540047(.x(x_47), .z(tmp00_47_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540048(.x(x_48), .z(tmp00_48_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540049(.x(x_49), .z(tmp00_49_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540050(.x(x_50), .z(tmp00_50_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540051(.x(x_51), .z(tmp00_51_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540052(.x(x_52), .z(tmp00_52_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540053(.x(x_53), .z(tmp00_53_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540054(.x(x_54), .z(tmp00_54_54));
	booth_0010 #(.WIDTH(WIDTH)) mul00540055(.x(x_55), .z(tmp00_55_54));
	booth__012 #(.WIDTH(WIDTH)) mul00540056(.x(x_56), .z(tmp00_56_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540057(.x(x_57), .z(tmp00_57_54));
	booth_0010 #(.WIDTH(WIDTH)) mul00540058(.x(x_58), .z(tmp00_58_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540059(.x(x_59), .z(tmp00_59_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540060(.x(x_60), .z(tmp00_60_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540061(.x(x_61), .z(tmp00_61_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540062(.x(x_62), .z(tmp00_62_54));
	booth_0006 #(.WIDTH(WIDTH)) mul00540063(.x(x_63), .z(tmp00_63_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540064(.x(x_64), .z(tmp00_64_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540065(.x(x_65), .z(tmp00_65_54));
	booth_0012 #(.WIDTH(WIDTH)) mul00540066(.x(x_66), .z(tmp00_66_54));
	booth_0002 #(.WIDTH(WIDTH)) mul00540067(.x(x_67), .z(tmp00_67_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540068(.x(x_68), .z(tmp00_68_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540069(.x(x_69), .z(tmp00_69_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540070(.x(x_70), .z(tmp00_70_54));
	booth__002 #(.WIDTH(WIDTH)) mul00540071(.x(x_71), .z(tmp00_71_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540072(.x(x_72), .z(tmp00_72_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540073(.x(x_73), .z(tmp00_73_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540074(.x(x_74), .z(tmp00_74_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540075(.x(x_75), .z(tmp00_75_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540076(.x(x_76), .z(tmp00_76_54));
	booth_0010 #(.WIDTH(WIDTH)) mul00540077(.x(x_77), .z(tmp00_77_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540078(.x(x_78), .z(tmp00_78_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540079(.x(x_79), .z(tmp00_79_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540080(.x(x_80), .z(tmp00_80_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540081(.x(x_81), .z(tmp00_81_54));
	booth_0012 #(.WIDTH(WIDTH)) mul00540082(.x(x_82), .z(tmp00_82_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540083(.x(x_83), .z(tmp00_83_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540084(.x(x_84), .z(tmp00_84_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540085(.x(x_85), .z(tmp00_85_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540086(.x(x_86), .z(tmp00_86_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540087(.x(x_87), .z(tmp00_87_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540088(.x(x_88), .z(tmp00_88_54));
	booth_0002 #(.WIDTH(WIDTH)) mul00540089(.x(x_89), .z(tmp00_89_54));
	booth__018 #(.WIDTH(WIDTH)) mul00540090(.x(x_90), .z(tmp00_90_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540091(.x(x_91), .z(tmp00_91_54));
	booth__010 #(.WIDTH(WIDTH)) mul00540092(.x(x_92), .z(tmp00_92_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540093(.x(x_93), .z(tmp00_93_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540094(.x(x_94), .z(tmp00_94_54));
	booth_0002 #(.WIDTH(WIDTH)) mul00540095(.x(x_95), .z(tmp00_95_54));
	booth_0020 #(.WIDTH(WIDTH)) mul00540096(.x(x_96), .z(tmp00_96_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540097(.x(x_97), .z(tmp00_97_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540098(.x(x_98), .z(tmp00_98_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540099(.x(x_99), .z(tmp00_99_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540100(.x(x_100), .z(tmp00_100_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540101(.x(x_101), .z(tmp00_101_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540102(.x(x_102), .z(tmp00_102_54));
	booth_0002 #(.WIDTH(WIDTH)) mul00540103(.x(x_103), .z(tmp00_103_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540104(.x(x_104), .z(tmp00_104_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540105(.x(x_105), .z(tmp00_105_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540106(.x(x_106), .z(tmp00_106_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540107(.x(x_107), .z(tmp00_107_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540108(.x(x_108), .z(tmp00_108_54));
	booth_0016 #(.WIDTH(WIDTH)) mul00540109(.x(x_109), .z(tmp00_109_54));
	booth_0016 #(.WIDTH(WIDTH)) mul00540110(.x(x_110), .z(tmp00_110_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540111(.x(x_111), .z(tmp00_111_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540112(.x(x_112), .z(tmp00_112_54));
	booth__016 #(.WIDTH(WIDTH)) mul00540113(.x(x_113), .z(tmp00_113_54));
	booth__008 #(.WIDTH(WIDTH)) mul00540114(.x(x_114), .z(tmp00_114_54));
	booth__004 #(.WIDTH(WIDTH)) mul00540115(.x(x_115), .z(tmp00_115_54));
	booth__006 #(.WIDTH(WIDTH)) mul00540116(.x(x_116), .z(tmp00_116_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540117(.x(x_117), .z(tmp00_117_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540118(.x(x_118), .z(tmp00_118_54));
	booth_0004 #(.WIDTH(WIDTH)) mul00540119(.x(x_119), .z(tmp00_119_54));
	booth_0000 #(.WIDTH(WIDTH)) mul00540120(.x(x_120), .z(tmp00_120_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540121(.x(x_121), .z(tmp00_121_54));
	booth_0010 #(.WIDTH(WIDTH)) mul00540122(.x(x_122), .z(tmp00_122_54));
	booth__010 #(.WIDTH(WIDTH)) mul00540123(.x(x_123), .z(tmp00_123_54));
	booth_0016 #(.WIDTH(WIDTH)) mul00540124(.x(x_124), .z(tmp00_124_54));
	booth_0008 #(.WIDTH(WIDTH)) mul00540125(.x(x_125), .z(tmp00_125_54));
	booth__006 #(.WIDTH(WIDTH)) mul00540126(.x(x_126), .z(tmp00_126_54));
	booth_0012 #(.WIDTH(WIDTH)) mul00540127(.x(x_127), .z(tmp00_127_54));
	booth__008 #(.WIDTH(WIDTH)) mul00550000(.x(x_0), .z(tmp00_0_55));
	booth_0010 #(.WIDTH(WIDTH)) mul00550001(.x(x_1), .z(tmp00_1_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550002(.x(x_2), .z(tmp00_2_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550003(.x(x_3), .z(tmp00_3_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550004(.x(x_4), .z(tmp00_4_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550005(.x(x_5), .z(tmp00_5_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550006(.x(x_6), .z(tmp00_6_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550007(.x(x_7), .z(tmp00_7_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550008(.x(x_8), .z(tmp00_8_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550009(.x(x_9), .z(tmp00_9_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550010(.x(x_10), .z(tmp00_10_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550011(.x(x_11), .z(tmp00_11_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550012(.x(x_12), .z(tmp00_12_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550013(.x(x_13), .z(tmp00_13_55));
	booth_0010 #(.WIDTH(WIDTH)) mul00550014(.x(x_14), .z(tmp00_14_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550015(.x(x_15), .z(tmp00_15_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550016(.x(x_16), .z(tmp00_16_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550017(.x(x_17), .z(tmp00_17_55));
	booth_0010 #(.WIDTH(WIDTH)) mul00550018(.x(x_18), .z(tmp00_18_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550019(.x(x_19), .z(tmp00_19_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550020(.x(x_20), .z(tmp00_20_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550021(.x(x_21), .z(tmp00_21_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550022(.x(x_22), .z(tmp00_22_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550023(.x(x_23), .z(tmp00_23_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550024(.x(x_24), .z(tmp00_24_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550025(.x(x_25), .z(tmp00_25_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550026(.x(x_26), .z(tmp00_26_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550027(.x(x_27), .z(tmp00_27_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550028(.x(x_28), .z(tmp00_28_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550029(.x(x_29), .z(tmp00_29_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550030(.x(x_30), .z(tmp00_30_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550031(.x(x_31), .z(tmp00_31_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550032(.x(x_32), .z(tmp00_32_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550033(.x(x_33), .z(tmp00_33_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550034(.x(x_34), .z(tmp00_34_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550035(.x(x_35), .z(tmp00_35_55));
	booth__010 #(.WIDTH(WIDTH)) mul00550036(.x(x_36), .z(tmp00_36_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550037(.x(x_37), .z(tmp00_37_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550038(.x(x_38), .z(tmp00_38_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550039(.x(x_39), .z(tmp00_39_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550040(.x(x_40), .z(tmp00_40_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550041(.x(x_41), .z(tmp00_41_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550042(.x(x_42), .z(tmp00_42_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550043(.x(x_43), .z(tmp00_43_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550044(.x(x_44), .z(tmp00_44_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550045(.x(x_45), .z(tmp00_45_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550046(.x(x_46), .z(tmp00_46_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550047(.x(x_47), .z(tmp00_47_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550048(.x(x_48), .z(tmp00_48_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550049(.x(x_49), .z(tmp00_49_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550050(.x(x_50), .z(tmp00_50_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550051(.x(x_51), .z(tmp00_51_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550052(.x(x_52), .z(tmp00_52_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550053(.x(x_53), .z(tmp00_53_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550054(.x(x_54), .z(tmp00_54_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550055(.x(x_55), .z(tmp00_55_55));
	booth__002 #(.WIDTH(WIDTH)) mul00550056(.x(x_56), .z(tmp00_56_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550057(.x(x_57), .z(tmp00_57_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550058(.x(x_58), .z(tmp00_58_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550059(.x(x_59), .z(tmp00_59_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550060(.x(x_60), .z(tmp00_60_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550061(.x(x_61), .z(tmp00_61_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550062(.x(x_62), .z(tmp00_62_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550063(.x(x_63), .z(tmp00_63_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550064(.x(x_64), .z(tmp00_64_55));
	booth__010 #(.WIDTH(WIDTH)) mul00550065(.x(x_65), .z(tmp00_65_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550066(.x(x_66), .z(tmp00_66_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550067(.x(x_67), .z(tmp00_67_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550068(.x(x_68), .z(tmp00_68_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550069(.x(x_69), .z(tmp00_69_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550070(.x(x_70), .z(tmp00_70_55));
	booth_0002 #(.WIDTH(WIDTH)) mul00550071(.x(x_71), .z(tmp00_71_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550072(.x(x_72), .z(tmp00_72_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550073(.x(x_73), .z(tmp00_73_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550074(.x(x_74), .z(tmp00_74_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550075(.x(x_75), .z(tmp00_75_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550076(.x(x_76), .z(tmp00_76_55));
	booth__012 #(.WIDTH(WIDTH)) mul00550077(.x(x_77), .z(tmp00_77_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550078(.x(x_78), .z(tmp00_78_55));
	booth_0012 #(.WIDTH(WIDTH)) mul00550079(.x(x_79), .z(tmp00_79_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550080(.x(x_80), .z(tmp00_80_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550081(.x(x_81), .z(tmp00_81_55));
	booth__012 #(.WIDTH(WIDTH)) mul00550082(.x(x_82), .z(tmp00_82_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550083(.x(x_83), .z(tmp00_83_55));
	booth_0010 #(.WIDTH(WIDTH)) mul00550084(.x(x_84), .z(tmp00_84_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550085(.x(x_85), .z(tmp00_85_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550086(.x(x_86), .z(tmp00_86_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550087(.x(x_87), .z(tmp00_87_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550088(.x(x_88), .z(tmp00_88_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550089(.x(x_89), .z(tmp00_89_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550090(.x(x_90), .z(tmp00_90_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550091(.x(x_91), .z(tmp00_91_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550092(.x(x_92), .z(tmp00_92_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550093(.x(x_93), .z(tmp00_93_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550094(.x(x_94), .z(tmp00_94_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550095(.x(x_95), .z(tmp00_95_55));
	booth_0006 #(.WIDTH(WIDTH)) mul00550096(.x(x_96), .z(tmp00_96_55));
	booth__002 #(.WIDTH(WIDTH)) mul00550097(.x(x_97), .z(tmp00_97_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550098(.x(x_98), .z(tmp00_98_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550099(.x(x_99), .z(tmp00_99_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550100(.x(x_100), .z(tmp00_100_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550101(.x(x_101), .z(tmp00_101_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550102(.x(x_102), .z(tmp00_102_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550103(.x(x_103), .z(tmp00_103_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550104(.x(x_104), .z(tmp00_104_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550105(.x(x_105), .z(tmp00_105_55));
	booth__008 #(.WIDTH(WIDTH)) mul00550106(.x(x_106), .z(tmp00_106_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550107(.x(x_107), .z(tmp00_107_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550108(.x(x_108), .z(tmp00_108_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550109(.x(x_109), .z(tmp00_109_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550110(.x(x_110), .z(tmp00_110_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550111(.x(x_111), .z(tmp00_111_55));
	booth_0006 #(.WIDTH(WIDTH)) mul00550112(.x(x_112), .z(tmp00_112_55));
	booth_0012 #(.WIDTH(WIDTH)) mul00550113(.x(x_113), .z(tmp00_113_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550114(.x(x_114), .z(tmp00_114_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550115(.x(x_115), .z(tmp00_115_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550116(.x(x_116), .z(tmp00_116_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550117(.x(x_117), .z(tmp00_117_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550118(.x(x_118), .z(tmp00_118_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550119(.x(x_119), .z(tmp00_119_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550120(.x(x_120), .z(tmp00_120_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550121(.x(x_121), .z(tmp00_121_55));
	booth__006 #(.WIDTH(WIDTH)) mul00550122(.x(x_122), .z(tmp00_122_55));
	booth_0008 #(.WIDTH(WIDTH)) mul00550123(.x(x_123), .z(tmp00_123_55));
	booth_0004 #(.WIDTH(WIDTH)) mul00550124(.x(x_124), .z(tmp00_124_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550125(.x(x_125), .z(tmp00_125_55));
	booth__004 #(.WIDTH(WIDTH)) mul00550126(.x(x_126), .z(tmp00_126_55));
	booth_0000 #(.WIDTH(WIDTH)) mul00550127(.x(x_127), .z(tmp00_127_55));
	booth__008 #(.WIDTH(WIDTH)) mul00560000(.x(x_0), .z(tmp00_0_56));
	booth_0002 #(.WIDTH(WIDTH)) mul00560001(.x(x_1), .z(tmp00_1_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560002(.x(x_2), .z(tmp00_2_56));
	booth__002 #(.WIDTH(WIDTH)) mul00560003(.x(x_3), .z(tmp00_3_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560004(.x(x_4), .z(tmp00_4_56));
	booth__010 #(.WIDTH(WIDTH)) mul00560005(.x(x_5), .z(tmp00_5_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560006(.x(x_6), .z(tmp00_6_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560007(.x(x_7), .z(tmp00_7_56));
	booth_0010 #(.WIDTH(WIDTH)) mul00560008(.x(x_8), .z(tmp00_8_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560009(.x(x_9), .z(tmp00_9_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560010(.x(x_10), .z(tmp00_10_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560011(.x(x_11), .z(tmp00_11_56));
	booth_0002 #(.WIDTH(WIDTH)) mul00560012(.x(x_12), .z(tmp00_12_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560013(.x(x_13), .z(tmp00_13_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560014(.x(x_14), .z(tmp00_14_56));
	booth__010 #(.WIDTH(WIDTH)) mul00560015(.x(x_15), .z(tmp00_15_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560016(.x(x_16), .z(tmp00_16_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560017(.x(x_17), .z(tmp00_17_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560018(.x(x_18), .z(tmp00_18_56));
	booth_0010 #(.WIDTH(WIDTH)) mul00560019(.x(x_19), .z(tmp00_19_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560020(.x(x_20), .z(tmp00_20_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560021(.x(x_21), .z(tmp00_21_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560022(.x(x_22), .z(tmp00_22_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560023(.x(x_23), .z(tmp00_23_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560024(.x(x_24), .z(tmp00_24_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560025(.x(x_25), .z(tmp00_25_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560026(.x(x_26), .z(tmp00_26_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560027(.x(x_27), .z(tmp00_27_56));
	booth_0010 #(.WIDTH(WIDTH)) mul00560028(.x(x_28), .z(tmp00_28_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560029(.x(x_29), .z(tmp00_29_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560030(.x(x_30), .z(tmp00_30_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560031(.x(x_31), .z(tmp00_31_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560032(.x(x_32), .z(tmp00_32_56));
	booth__010 #(.WIDTH(WIDTH)) mul00560033(.x(x_33), .z(tmp00_33_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560034(.x(x_34), .z(tmp00_34_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560035(.x(x_35), .z(tmp00_35_56));
	booth_0006 #(.WIDTH(WIDTH)) mul00560036(.x(x_36), .z(tmp00_36_56));
	booth_0010 #(.WIDTH(WIDTH)) mul00560037(.x(x_37), .z(tmp00_37_56));
	booth_0006 #(.WIDTH(WIDTH)) mul00560038(.x(x_38), .z(tmp00_38_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560039(.x(x_39), .z(tmp00_39_56));
	booth__002 #(.WIDTH(WIDTH)) mul00560040(.x(x_40), .z(tmp00_40_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560041(.x(x_41), .z(tmp00_41_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560042(.x(x_42), .z(tmp00_42_56));
	booth__010 #(.WIDTH(WIDTH)) mul00560043(.x(x_43), .z(tmp00_43_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560044(.x(x_44), .z(tmp00_44_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560045(.x(x_45), .z(tmp00_45_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560046(.x(x_46), .z(tmp00_46_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560047(.x(x_47), .z(tmp00_47_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560048(.x(x_48), .z(tmp00_48_56));
	booth__002 #(.WIDTH(WIDTH)) mul00560049(.x(x_49), .z(tmp00_49_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560050(.x(x_50), .z(tmp00_50_56));
	booth_0002 #(.WIDTH(WIDTH)) mul00560051(.x(x_51), .z(tmp00_51_56));
	booth_0010 #(.WIDTH(WIDTH)) mul00560052(.x(x_52), .z(tmp00_52_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560053(.x(x_53), .z(tmp00_53_56));
	booth__002 #(.WIDTH(WIDTH)) mul00560054(.x(x_54), .z(tmp00_54_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560055(.x(x_55), .z(tmp00_55_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560056(.x(x_56), .z(tmp00_56_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560057(.x(x_57), .z(tmp00_57_56));
	booth__002 #(.WIDTH(WIDTH)) mul00560058(.x(x_58), .z(tmp00_58_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560059(.x(x_59), .z(tmp00_59_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560060(.x(x_60), .z(tmp00_60_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560061(.x(x_61), .z(tmp00_61_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560062(.x(x_62), .z(tmp00_62_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560063(.x(x_63), .z(tmp00_63_56));
	booth__006 #(.WIDTH(WIDTH)) mul00560064(.x(x_64), .z(tmp00_64_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560065(.x(x_65), .z(tmp00_65_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560066(.x(x_66), .z(tmp00_66_56));
	booth__010 #(.WIDTH(WIDTH)) mul00560067(.x(x_67), .z(tmp00_67_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560068(.x(x_68), .z(tmp00_68_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560069(.x(x_69), .z(tmp00_69_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560070(.x(x_70), .z(tmp00_70_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560071(.x(x_71), .z(tmp00_71_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560072(.x(x_72), .z(tmp00_72_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560073(.x(x_73), .z(tmp00_73_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560074(.x(x_74), .z(tmp00_74_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560075(.x(x_75), .z(tmp00_75_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560076(.x(x_76), .z(tmp00_76_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560077(.x(x_77), .z(tmp00_77_56));
	booth__002 #(.WIDTH(WIDTH)) mul00560078(.x(x_78), .z(tmp00_78_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560079(.x(x_79), .z(tmp00_79_56));
	booth__002 #(.WIDTH(WIDTH)) mul00560080(.x(x_80), .z(tmp00_80_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560081(.x(x_81), .z(tmp00_81_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560082(.x(x_82), .z(tmp00_82_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560083(.x(x_83), .z(tmp00_83_56));
	booth__006 #(.WIDTH(WIDTH)) mul00560084(.x(x_84), .z(tmp00_84_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560085(.x(x_85), .z(tmp00_85_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560086(.x(x_86), .z(tmp00_86_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560087(.x(x_87), .z(tmp00_87_56));
	booth__010 #(.WIDTH(WIDTH)) mul00560088(.x(x_88), .z(tmp00_88_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560089(.x(x_89), .z(tmp00_89_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560090(.x(x_90), .z(tmp00_90_56));
	booth__006 #(.WIDTH(WIDTH)) mul00560091(.x(x_91), .z(tmp00_91_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560092(.x(x_92), .z(tmp00_92_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560093(.x(x_93), .z(tmp00_93_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560094(.x(x_94), .z(tmp00_94_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560095(.x(x_95), .z(tmp00_95_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560096(.x(x_96), .z(tmp00_96_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560097(.x(x_97), .z(tmp00_97_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560098(.x(x_98), .z(tmp00_98_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560099(.x(x_99), .z(tmp00_99_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560100(.x(x_100), .z(tmp00_100_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560101(.x(x_101), .z(tmp00_101_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560102(.x(x_102), .z(tmp00_102_56));
	booth__006 #(.WIDTH(WIDTH)) mul00560103(.x(x_103), .z(tmp00_103_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560104(.x(x_104), .z(tmp00_104_56));
	booth__002 #(.WIDTH(WIDTH)) mul00560105(.x(x_105), .z(tmp00_105_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560106(.x(x_106), .z(tmp00_106_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560107(.x(x_107), .z(tmp00_107_56));
	booth_0002 #(.WIDTH(WIDTH)) mul00560108(.x(x_108), .z(tmp00_108_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560109(.x(x_109), .z(tmp00_109_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560110(.x(x_110), .z(tmp00_110_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560111(.x(x_111), .z(tmp00_111_56));
	booth_0008 #(.WIDTH(WIDTH)) mul00560112(.x(x_112), .z(tmp00_112_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560113(.x(x_113), .z(tmp00_113_56));
	booth_0006 #(.WIDTH(WIDTH)) mul00560114(.x(x_114), .z(tmp00_114_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560115(.x(x_115), .z(tmp00_115_56));
	booth__004 #(.WIDTH(WIDTH)) mul00560116(.x(x_116), .z(tmp00_116_56));
	booth_0004 #(.WIDTH(WIDTH)) mul00560117(.x(x_117), .z(tmp00_117_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560118(.x(x_118), .z(tmp00_118_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560119(.x(x_119), .z(tmp00_119_56));
	booth__010 #(.WIDTH(WIDTH)) mul00560120(.x(x_120), .z(tmp00_120_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560121(.x(x_121), .z(tmp00_121_56));
	booth_0002 #(.WIDTH(WIDTH)) mul00560122(.x(x_122), .z(tmp00_122_56));
	booth__008 #(.WIDTH(WIDTH)) mul00560123(.x(x_123), .z(tmp00_123_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560124(.x(x_124), .z(tmp00_124_56));
	booth_0010 #(.WIDTH(WIDTH)) mul00560125(.x(x_125), .z(tmp00_125_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00560126(.x(x_126), .z(tmp00_126_56));
	booth__010 #(.WIDTH(WIDTH)) mul00560127(.x(x_127), .z(tmp00_127_56));
	booth_0000 #(.WIDTH(WIDTH)) mul00570000(.x(x_0), .z(tmp00_0_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570001(.x(x_1), .z(tmp00_1_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570002(.x(x_2), .z(tmp00_2_57));
	booth__006 #(.WIDTH(WIDTH)) mul00570003(.x(x_3), .z(tmp00_3_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570004(.x(x_4), .z(tmp00_4_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570005(.x(x_5), .z(tmp00_5_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570006(.x(x_6), .z(tmp00_6_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570007(.x(x_7), .z(tmp00_7_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570008(.x(x_8), .z(tmp00_8_57));
	booth_0010 #(.WIDTH(WIDTH)) mul00570009(.x(x_9), .z(tmp00_9_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570010(.x(x_10), .z(tmp00_10_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570011(.x(x_11), .z(tmp00_11_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570012(.x(x_12), .z(tmp00_12_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570013(.x(x_13), .z(tmp00_13_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570014(.x(x_14), .z(tmp00_14_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570015(.x(x_15), .z(tmp00_15_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570016(.x(x_16), .z(tmp00_16_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570017(.x(x_17), .z(tmp00_17_57));
	booth__006 #(.WIDTH(WIDTH)) mul00570018(.x(x_18), .z(tmp00_18_57));
	booth__010 #(.WIDTH(WIDTH)) mul00570019(.x(x_19), .z(tmp00_19_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570020(.x(x_20), .z(tmp00_20_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570021(.x(x_21), .z(tmp00_21_57));
	booth_0002 #(.WIDTH(WIDTH)) mul00570022(.x(x_22), .z(tmp00_22_57));
	booth__012 #(.WIDTH(WIDTH)) mul00570023(.x(x_23), .z(tmp00_23_57));
	booth_0002 #(.WIDTH(WIDTH)) mul00570024(.x(x_24), .z(tmp00_24_57));
	booth_0012 #(.WIDTH(WIDTH)) mul00570025(.x(x_25), .z(tmp00_25_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570026(.x(x_26), .z(tmp00_26_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570027(.x(x_27), .z(tmp00_27_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570028(.x(x_28), .z(tmp00_28_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570029(.x(x_29), .z(tmp00_29_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570030(.x(x_30), .z(tmp00_30_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570031(.x(x_31), .z(tmp00_31_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570032(.x(x_32), .z(tmp00_32_57));
	booth__002 #(.WIDTH(WIDTH)) mul00570033(.x(x_33), .z(tmp00_33_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570034(.x(x_34), .z(tmp00_34_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570035(.x(x_35), .z(tmp00_35_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570036(.x(x_36), .z(tmp00_36_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570037(.x(x_37), .z(tmp00_37_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570038(.x(x_38), .z(tmp00_38_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570039(.x(x_39), .z(tmp00_39_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570040(.x(x_40), .z(tmp00_40_57));
	booth_0006 #(.WIDTH(WIDTH)) mul00570041(.x(x_41), .z(tmp00_41_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570042(.x(x_42), .z(tmp00_42_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570043(.x(x_43), .z(tmp00_43_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570044(.x(x_44), .z(tmp00_44_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570045(.x(x_45), .z(tmp00_45_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570046(.x(x_46), .z(tmp00_46_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570047(.x(x_47), .z(tmp00_47_57));
	booth_0002 #(.WIDTH(WIDTH)) mul00570048(.x(x_48), .z(tmp00_48_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570049(.x(x_49), .z(tmp00_49_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570050(.x(x_50), .z(tmp00_50_57));
	booth__010 #(.WIDTH(WIDTH)) mul00570051(.x(x_51), .z(tmp00_51_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570052(.x(x_52), .z(tmp00_52_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570053(.x(x_53), .z(tmp00_53_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570054(.x(x_54), .z(tmp00_54_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570055(.x(x_55), .z(tmp00_55_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570056(.x(x_56), .z(tmp00_56_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570057(.x(x_57), .z(tmp00_57_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570058(.x(x_58), .z(tmp00_58_57));
	booth_0012 #(.WIDTH(WIDTH)) mul00570059(.x(x_59), .z(tmp00_59_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570060(.x(x_60), .z(tmp00_60_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570061(.x(x_61), .z(tmp00_61_57));
	booth_0006 #(.WIDTH(WIDTH)) mul00570062(.x(x_62), .z(tmp00_62_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570063(.x(x_63), .z(tmp00_63_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570064(.x(x_64), .z(tmp00_64_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570065(.x(x_65), .z(tmp00_65_57));
	booth__002 #(.WIDTH(WIDTH)) mul00570066(.x(x_66), .z(tmp00_66_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570067(.x(x_67), .z(tmp00_67_57));
	booth_0012 #(.WIDTH(WIDTH)) mul00570068(.x(x_68), .z(tmp00_68_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570069(.x(x_69), .z(tmp00_69_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570070(.x(x_70), .z(tmp00_70_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570071(.x(x_71), .z(tmp00_71_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570072(.x(x_72), .z(tmp00_72_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570073(.x(x_73), .z(tmp00_73_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570074(.x(x_74), .z(tmp00_74_57));
	booth_0012 #(.WIDTH(WIDTH)) mul00570075(.x(x_75), .z(tmp00_75_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570076(.x(x_76), .z(tmp00_76_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570077(.x(x_77), .z(tmp00_77_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570078(.x(x_78), .z(tmp00_78_57));
	booth__010 #(.WIDTH(WIDTH)) mul00570079(.x(x_79), .z(tmp00_79_57));
	booth_0006 #(.WIDTH(WIDTH)) mul00570080(.x(x_80), .z(tmp00_80_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570081(.x(x_81), .z(tmp00_81_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570082(.x(x_82), .z(tmp00_82_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570083(.x(x_83), .z(tmp00_83_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570084(.x(x_84), .z(tmp00_84_57));
	booth_0012 #(.WIDTH(WIDTH)) mul00570085(.x(x_85), .z(tmp00_85_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570086(.x(x_86), .z(tmp00_86_57));
	booth_0012 #(.WIDTH(WIDTH)) mul00570087(.x(x_87), .z(tmp00_87_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570088(.x(x_88), .z(tmp00_88_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570089(.x(x_89), .z(tmp00_89_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570090(.x(x_90), .z(tmp00_90_57));
	booth__010 #(.WIDTH(WIDTH)) mul00570091(.x(x_91), .z(tmp00_91_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570092(.x(x_92), .z(tmp00_92_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570093(.x(x_93), .z(tmp00_93_57));
	booth__006 #(.WIDTH(WIDTH)) mul00570094(.x(x_94), .z(tmp00_94_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570095(.x(x_95), .z(tmp00_95_57));
	booth__004 #(.WIDTH(WIDTH)) mul00570096(.x(x_96), .z(tmp00_96_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570097(.x(x_97), .z(tmp00_97_57));
	booth__002 #(.WIDTH(WIDTH)) mul00570098(.x(x_98), .z(tmp00_98_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570099(.x(x_99), .z(tmp00_99_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570100(.x(x_100), .z(tmp00_100_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570101(.x(x_101), .z(tmp00_101_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570102(.x(x_102), .z(tmp00_102_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570103(.x(x_103), .z(tmp00_103_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570104(.x(x_104), .z(tmp00_104_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570105(.x(x_105), .z(tmp00_105_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570106(.x(x_106), .z(tmp00_106_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570107(.x(x_107), .z(tmp00_107_57));
	booth_0012 #(.WIDTH(WIDTH)) mul00570108(.x(x_108), .z(tmp00_108_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570109(.x(x_109), .z(tmp00_109_57));
	booth_0002 #(.WIDTH(WIDTH)) mul00570110(.x(x_110), .z(tmp00_110_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570111(.x(x_111), .z(tmp00_111_57));
	booth_0010 #(.WIDTH(WIDTH)) mul00570112(.x(x_112), .z(tmp00_112_57));
	booth_0008 #(.WIDTH(WIDTH)) mul00570113(.x(x_113), .z(tmp00_113_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570114(.x(x_114), .z(tmp00_114_57));
	booth__002 #(.WIDTH(WIDTH)) mul00570115(.x(x_115), .z(tmp00_115_57));
	booth__010 #(.WIDTH(WIDTH)) mul00570116(.x(x_116), .z(tmp00_116_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570117(.x(x_117), .z(tmp00_117_57));
	booth__002 #(.WIDTH(WIDTH)) mul00570118(.x(x_118), .z(tmp00_118_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570119(.x(x_119), .z(tmp00_119_57));
	booth_0012 #(.WIDTH(WIDTH)) mul00570120(.x(x_120), .z(tmp00_120_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570121(.x(x_121), .z(tmp00_121_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570122(.x(x_122), .z(tmp00_122_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570123(.x(x_123), .z(tmp00_123_57));
	booth__008 #(.WIDTH(WIDTH)) mul00570124(.x(x_124), .z(tmp00_124_57));
	booth_0004 #(.WIDTH(WIDTH)) mul00570125(.x(x_125), .z(tmp00_125_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570126(.x(x_126), .z(tmp00_126_57));
	booth_0000 #(.WIDTH(WIDTH)) mul00570127(.x(x_127), .z(tmp00_127_57));
	booth_0002 #(.WIDTH(WIDTH)) mul00580000(.x(x_0), .z(tmp00_0_58));
	booth_0010 #(.WIDTH(WIDTH)) mul00580001(.x(x_1), .z(tmp00_1_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580002(.x(x_2), .z(tmp00_2_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580003(.x(x_3), .z(tmp00_3_58));
	booth__004 #(.WIDTH(WIDTH)) mul00580004(.x(x_4), .z(tmp00_4_58));
	booth_0006 #(.WIDTH(WIDTH)) mul00580005(.x(x_5), .z(tmp00_5_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580006(.x(x_6), .z(tmp00_6_58));
	booth_0010 #(.WIDTH(WIDTH)) mul00580007(.x(x_7), .z(tmp00_7_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580008(.x(x_8), .z(tmp00_8_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580009(.x(x_9), .z(tmp00_9_58));
	booth_0012 #(.WIDTH(WIDTH)) mul00580010(.x(x_10), .z(tmp00_10_58));
	booth_0010 #(.WIDTH(WIDTH)) mul00580011(.x(x_11), .z(tmp00_11_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580012(.x(x_12), .z(tmp00_12_58));
	booth_0012 #(.WIDTH(WIDTH)) mul00580013(.x(x_13), .z(tmp00_13_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580014(.x(x_14), .z(tmp00_14_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580015(.x(x_15), .z(tmp00_15_58));
	booth_0012 #(.WIDTH(WIDTH)) mul00580016(.x(x_16), .z(tmp00_16_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580017(.x(x_17), .z(tmp00_17_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580018(.x(x_18), .z(tmp00_18_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580019(.x(x_19), .z(tmp00_19_58));
	booth__014 #(.WIDTH(WIDTH)) mul00580020(.x(x_20), .z(tmp00_20_58));
	booth__006 #(.WIDTH(WIDTH)) mul00580021(.x(x_21), .z(tmp00_21_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580022(.x(x_22), .z(tmp00_22_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580023(.x(x_23), .z(tmp00_23_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580024(.x(x_24), .z(tmp00_24_58));
	booth_0014 #(.WIDTH(WIDTH)) mul00580025(.x(x_25), .z(tmp00_25_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580026(.x(x_26), .z(tmp00_26_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580027(.x(x_27), .z(tmp00_27_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580028(.x(x_28), .z(tmp00_28_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580029(.x(x_29), .z(tmp00_29_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580030(.x(x_30), .z(tmp00_30_58));
	booth__004 #(.WIDTH(WIDTH)) mul00580031(.x(x_31), .z(tmp00_31_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580032(.x(x_32), .z(tmp00_32_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580033(.x(x_33), .z(tmp00_33_58));
	booth_0006 #(.WIDTH(WIDTH)) mul00580034(.x(x_34), .z(tmp00_34_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580035(.x(x_35), .z(tmp00_35_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580036(.x(x_36), .z(tmp00_36_58));
	booth_0002 #(.WIDTH(WIDTH)) mul00580037(.x(x_37), .z(tmp00_37_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580038(.x(x_38), .z(tmp00_38_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580039(.x(x_39), .z(tmp00_39_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580040(.x(x_40), .z(tmp00_40_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580041(.x(x_41), .z(tmp00_41_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580042(.x(x_42), .z(tmp00_42_58));
	booth_0010 #(.WIDTH(WIDTH)) mul00580043(.x(x_43), .z(tmp00_43_58));
	booth__004 #(.WIDTH(WIDTH)) mul00580044(.x(x_44), .z(tmp00_44_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580045(.x(x_45), .z(tmp00_45_58));
	booth__012 #(.WIDTH(WIDTH)) mul00580046(.x(x_46), .z(tmp00_46_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580047(.x(x_47), .z(tmp00_47_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580048(.x(x_48), .z(tmp00_48_58));
	booth_0012 #(.WIDTH(WIDTH)) mul00580049(.x(x_49), .z(tmp00_49_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580050(.x(x_50), .z(tmp00_50_58));
	booth__010 #(.WIDTH(WIDTH)) mul00580051(.x(x_51), .z(tmp00_51_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580052(.x(x_52), .z(tmp00_52_58));
	booth__004 #(.WIDTH(WIDTH)) mul00580053(.x(x_53), .z(tmp00_53_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580054(.x(x_54), .z(tmp00_54_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580055(.x(x_55), .z(tmp00_55_58));
	booth_0010 #(.WIDTH(WIDTH)) mul00580056(.x(x_56), .z(tmp00_56_58));
	booth_0010 #(.WIDTH(WIDTH)) mul00580057(.x(x_57), .z(tmp00_57_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580058(.x(x_58), .z(tmp00_58_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580059(.x(x_59), .z(tmp00_59_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580060(.x(x_60), .z(tmp00_60_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580061(.x(x_61), .z(tmp00_61_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580062(.x(x_62), .z(tmp00_62_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580063(.x(x_63), .z(tmp00_63_58));
	booth_0006 #(.WIDTH(WIDTH)) mul00580064(.x(x_64), .z(tmp00_64_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580065(.x(x_65), .z(tmp00_65_58));
	booth_0002 #(.WIDTH(WIDTH)) mul00580066(.x(x_66), .z(tmp00_66_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580067(.x(x_67), .z(tmp00_67_58));
	booth__004 #(.WIDTH(WIDTH)) mul00580068(.x(x_68), .z(tmp00_68_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580069(.x(x_69), .z(tmp00_69_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580070(.x(x_70), .z(tmp00_70_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580071(.x(x_71), .z(tmp00_71_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580072(.x(x_72), .z(tmp00_72_58));
	booth__004 #(.WIDTH(WIDTH)) mul00580073(.x(x_73), .z(tmp00_73_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580074(.x(x_74), .z(tmp00_74_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580075(.x(x_75), .z(tmp00_75_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580076(.x(x_76), .z(tmp00_76_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580077(.x(x_77), .z(tmp00_77_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580078(.x(x_78), .z(tmp00_78_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580079(.x(x_79), .z(tmp00_79_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580080(.x(x_80), .z(tmp00_80_58));
	booth__004 #(.WIDTH(WIDTH)) mul00580081(.x(x_81), .z(tmp00_81_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580082(.x(x_82), .z(tmp00_82_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580083(.x(x_83), .z(tmp00_83_58));
	booth__006 #(.WIDTH(WIDTH)) mul00580084(.x(x_84), .z(tmp00_84_58));
	booth__012 #(.WIDTH(WIDTH)) mul00580085(.x(x_85), .z(tmp00_85_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580086(.x(x_86), .z(tmp00_86_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580087(.x(x_87), .z(tmp00_87_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580088(.x(x_88), .z(tmp00_88_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580089(.x(x_89), .z(tmp00_89_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580090(.x(x_90), .z(tmp00_90_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580091(.x(x_91), .z(tmp00_91_58));
	booth_0002 #(.WIDTH(WIDTH)) mul00580092(.x(x_92), .z(tmp00_92_58));
	booth__006 #(.WIDTH(WIDTH)) mul00580093(.x(x_93), .z(tmp00_93_58));
	booth_0002 #(.WIDTH(WIDTH)) mul00580094(.x(x_94), .z(tmp00_94_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580095(.x(x_95), .z(tmp00_95_58));
	booth__010 #(.WIDTH(WIDTH)) mul00580096(.x(x_96), .z(tmp00_96_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580097(.x(x_97), .z(tmp00_97_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580098(.x(x_98), .z(tmp00_98_58));
	booth__002 #(.WIDTH(WIDTH)) mul00580099(.x(x_99), .z(tmp00_99_58));
	booth__010 #(.WIDTH(WIDTH)) mul00580100(.x(x_100), .z(tmp00_100_58));
	booth__002 #(.WIDTH(WIDTH)) mul00580101(.x(x_101), .z(tmp00_101_58));
	booth__012 #(.WIDTH(WIDTH)) mul00580102(.x(x_102), .z(tmp00_102_58));
	booth__004 #(.WIDTH(WIDTH)) mul00580103(.x(x_103), .z(tmp00_103_58));
	booth__010 #(.WIDTH(WIDTH)) mul00580104(.x(x_104), .z(tmp00_104_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580105(.x(x_105), .z(tmp00_105_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580106(.x(x_106), .z(tmp00_106_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580107(.x(x_107), .z(tmp00_107_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580108(.x(x_108), .z(tmp00_108_58));
	booth__016 #(.WIDTH(WIDTH)) mul00580109(.x(x_109), .z(tmp00_109_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580110(.x(x_110), .z(tmp00_110_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580111(.x(x_111), .z(tmp00_111_58));
	booth__008 #(.WIDTH(WIDTH)) mul00580112(.x(x_112), .z(tmp00_112_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580113(.x(x_113), .z(tmp00_113_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580114(.x(x_114), .z(tmp00_114_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580115(.x(x_115), .z(tmp00_115_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580116(.x(x_116), .z(tmp00_116_58));
	booth__002 #(.WIDTH(WIDTH)) mul00580117(.x(x_117), .z(tmp00_117_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580118(.x(x_118), .z(tmp00_118_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580119(.x(x_119), .z(tmp00_119_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580120(.x(x_120), .z(tmp00_120_58));
	booth__002 #(.WIDTH(WIDTH)) mul00580121(.x(x_121), .z(tmp00_121_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580122(.x(x_122), .z(tmp00_122_58));
	booth_0000 #(.WIDTH(WIDTH)) mul00580123(.x(x_123), .z(tmp00_123_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580124(.x(x_124), .z(tmp00_124_58));
	booth_0008 #(.WIDTH(WIDTH)) mul00580125(.x(x_125), .z(tmp00_125_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580126(.x(x_126), .z(tmp00_126_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00580127(.x(x_127), .z(tmp00_127_58));
	booth_0004 #(.WIDTH(WIDTH)) mul00590000(.x(x_0), .z(tmp00_0_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590001(.x(x_1), .z(tmp00_1_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590002(.x(x_2), .z(tmp00_2_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590003(.x(x_3), .z(tmp00_3_59));
	booth_0012 #(.WIDTH(WIDTH)) mul00590004(.x(x_4), .z(tmp00_4_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590005(.x(x_5), .z(tmp00_5_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590006(.x(x_6), .z(tmp00_6_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590007(.x(x_7), .z(tmp00_7_59));
	booth_0012 #(.WIDTH(WIDTH)) mul00590008(.x(x_8), .z(tmp00_8_59));
	booth_0002 #(.WIDTH(WIDTH)) mul00590009(.x(x_9), .z(tmp00_9_59));
	booth__006 #(.WIDTH(WIDTH)) mul00590010(.x(x_10), .z(tmp00_10_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590011(.x(x_11), .z(tmp00_11_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590012(.x(x_12), .z(tmp00_12_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590013(.x(x_13), .z(tmp00_13_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590014(.x(x_14), .z(tmp00_14_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590015(.x(x_15), .z(tmp00_15_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590016(.x(x_16), .z(tmp00_16_59));
	booth_0012 #(.WIDTH(WIDTH)) mul00590017(.x(x_17), .z(tmp00_17_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590018(.x(x_18), .z(tmp00_18_59));
	booth_0002 #(.WIDTH(WIDTH)) mul00590019(.x(x_19), .z(tmp00_19_59));
	booth_0014 #(.WIDTH(WIDTH)) mul00590020(.x(x_20), .z(tmp00_20_59));
	booth__002 #(.WIDTH(WIDTH)) mul00590021(.x(x_21), .z(tmp00_21_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590022(.x(x_22), .z(tmp00_22_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590023(.x(x_23), .z(tmp00_23_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590024(.x(x_24), .z(tmp00_24_59));
	booth__014 #(.WIDTH(WIDTH)) mul00590025(.x(x_25), .z(tmp00_25_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590026(.x(x_26), .z(tmp00_26_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590027(.x(x_27), .z(tmp00_27_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590028(.x(x_28), .z(tmp00_28_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590029(.x(x_29), .z(tmp00_29_59));
	booth__002 #(.WIDTH(WIDTH)) mul00590030(.x(x_30), .z(tmp00_30_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590031(.x(x_31), .z(tmp00_31_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590032(.x(x_32), .z(tmp00_32_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590033(.x(x_33), .z(tmp00_33_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590034(.x(x_34), .z(tmp00_34_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590035(.x(x_35), .z(tmp00_35_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590036(.x(x_36), .z(tmp00_36_59));
	booth__002 #(.WIDTH(WIDTH)) mul00590037(.x(x_37), .z(tmp00_37_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590038(.x(x_38), .z(tmp00_38_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590039(.x(x_39), .z(tmp00_39_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590040(.x(x_40), .z(tmp00_40_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590041(.x(x_41), .z(tmp00_41_59));
	booth__020 #(.WIDTH(WIDTH)) mul00590042(.x(x_42), .z(tmp00_42_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590043(.x(x_43), .z(tmp00_43_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590044(.x(x_44), .z(tmp00_44_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590045(.x(x_45), .z(tmp00_45_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590046(.x(x_46), .z(tmp00_46_59));
	booth__012 #(.WIDTH(WIDTH)) mul00590047(.x(x_47), .z(tmp00_47_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590048(.x(x_48), .z(tmp00_48_59));
	booth__002 #(.WIDTH(WIDTH)) mul00590049(.x(x_49), .z(tmp00_49_59));
	booth__010 #(.WIDTH(WIDTH)) mul00590050(.x(x_50), .z(tmp00_50_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590051(.x(x_51), .z(tmp00_51_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590052(.x(x_52), .z(tmp00_52_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590053(.x(x_53), .z(tmp00_53_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590054(.x(x_54), .z(tmp00_54_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590055(.x(x_55), .z(tmp00_55_59));
	booth__016 #(.WIDTH(WIDTH)) mul00590056(.x(x_56), .z(tmp00_56_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590057(.x(x_57), .z(tmp00_57_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590058(.x(x_58), .z(tmp00_58_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590059(.x(x_59), .z(tmp00_59_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590060(.x(x_60), .z(tmp00_60_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590061(.x(x_61), .z(tmp00_61_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590062(.x(x_62), .z(tmp00_62_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590063(.x(x_63), .z(tmp00_63_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590064(.x(x_64), .z(tmp00_64_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590065(.x(x_65), .z(tmp00_65_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590066(.x(x_66), .z(tmp00_66_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590067(.x(x_67), .z(tmp00_67_59));
	booth__014 #(.WIDTH(WIDTH)) mul00590068(.x(x_68), .z(tmp00_68_59));
	booth__002 #(.WIDTH(WIDTH)) mul00590069(.x(x_69), .z(tmp00_69_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590070(.x(x_70), .z(tmp00_70_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590071(.x(x_71), .z(tmp00_71_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590072(.x(x_72), .z(tmp00_72_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590073(.x(x_73), .z(tmp00_73_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590074(.x(x_74), .z(tmp00_74_59));
	booth_0024 #(.WIDTH(WIDTH)) mul00590075(.x(x_75), .z(tmp00_75_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590076(.x(x_76), .z(tmp00_76_59));
	booth_0002 #(.WIDTH(WIDTH)) mul00590077(.x(x_77), .z(tmp00_77_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590078(.x(x_78), .z(tmp00_78_59));
	booth__010 #(.WIDTH(WIDTH)) mul00590079(.x(x_79), .z(tmp00_79_59));
	booth__014 #(.WIDTH(WIDTH)) mul00590080(.x(x_80), .z(tmp00_80_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590081(.x(x_81), .z(tmp00_81_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590082(.x(x_82), .z(tmp00_82_59));
	booth_0010 #(.WIDTH(WIDTH)) mul00590083(.x(x_83), .z(tmp00_83_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590084(.x(x_84), .z(tmp00_84_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590085(.x(x_85), .z(tmp00_85_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590086(.x(x_86), .z(tmp00_86_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590087(.x(x_87), .z(tmp00_87_59));
	booth_0002 #(.WIDTH(WIDTH)) mul00590088(.x(x_88), .z(tmp00_88_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590089(.x(x_89), .z(tmp00_89_59));
	booth__020 #(.WIDTH(WIDTH)) mul00590090(.x(x_90), .z(tmp00_90_59));
	booth__002 #(.WIDTH(WIDTH)) mul00590091(.x(x_91), .z(tmp00_91_59));
	booth__006 #(.WIDTH(WIDTH)) mul00590092(.x(x_92), .z(tmp00_92_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590093(.x(x_93), .z(tmp00_93_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590094(.x(x_94), .z(tmp00_94_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590095(.x(x_95), .z(tmp00_95_59));
	booth_0020 #(.WIDTH(WIDTH)) mul00590096(.x(x_96), .z(tmp00_96_59));
	booth_0002 #(.WIDTH(WIDTH)) mul00590097(.x(x_97), .z(tmp00_97_59));
	booth_0010 #(.WIDTH(WIDTH)) mul00590098(.x(x_98), .z(tmp00_98_59));
	booth_0012 #(.WIDTH(WIDTH)) mul00590099(.x(x_99), .z(tmp00_99_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590100(.x(x_100), .z(tmp00_100_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590101(.x(x_101), .z(tmp00_101_59));
	booth_0002 #(.WIDTH(WIDTH)) mul00590102(.x(x_102), .z(tmp00_102_59));
	booth__012 #(.WIDTH(WIDTH)) mul00590103(.x(x_103), .z(tmp00_103_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590104(.x(x_104), .z(tmp00_104_59));
	booth_0006 #(.WIDTH(WIDTH)) mul00590105(.x(x_105), .z(tmp00_105_59));
	booth_0002 #(.WIDTH(WIDTH)) mul00590106(.x(x_106), .z(tmp00_106_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590107(.x(x_107), .z(tmp00_107_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590108(.x(x_108), .z(tmp00_108_59));
	booth_0020 #(.WIDTH(WIDTH)) mul00590109(.x(x_109), .z(tmp00_109_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590110(.x(x_110), .z(tmp00_110_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590111(.x(x_111), .z(tmp00_111_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590112(.x(x_112), .z(tmp00_112_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590113(.x(x_113), .z(tmp00_113_59));
	booth__012 #(.WIDTH(WIDTH)) mul00590114(.x(x_114), .z(tmp00_114_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590115(.x(x_115), .z(tmp00_115_59));
	booth__008 #(.WIDTH(WIDTH)) mul00590116(.x(x_116), .z(tmp00_116_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590117(.x(x_117), .z(tmp00_117_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590118(.x(x_118), .z(tmp00_118_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590119(.x(x_119), .z(tmp00_119_59));
	booth_0006 #(.WIDTH(WIDTH)) mul00590120(.x(x_120), .z(tmp00_120_59));
	booth_0008 #(.WIDTH(WIDTH)) mul00590121(.x(x_121), .z(tmp00_121_59));
	booth_0004 #(.WIDTH(WIDTH)) mul00590122(.x(x_122), .z(tmp00_122_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590123(.x(x_123), .z(tmp00_123_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590124(.x(x_124), .z(tmp00_124_59));
	booth_0000 #(.WIDTH(WIDTH)) mul00590125(.x(x_125), .z(tmp00_125_59));
	booth__004 #(.WIDTH(WIDTH)) mul00590126(.x(x_126), .z(tmp00_126_59));
	booth_0016 #(.WIDTH(WIDTH)) mul00590127(.x(x_127), .z(tmp00_127_59));
	booth_0002 #(.WIDTH(WIDTH)) mul00600000(.x(x_0), .z(tmp00_0_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600001(.x(x_1), .z(tmp00_1_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600002(.x(x_2), .z(tmp00_2_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600003(.x(x_3), .z(tmp00_3_60));
	booth__006 #(.WIDTH(WIDTH)) mul00600004(.x(x_4), .z(tmp00_4_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600005(.x(x_5), .z(tmp00_5_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600006(.x(x_6), .z(tmp00_6_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600007(.x(x_7), .z(tmp00_7_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600008(.x(x_8), .z(tmp00_8_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600009(.x(x_9), .z(tmp00_9_60));
	booth__010 #(.WIDTH(WIDTH)) mul00600010(.x(x_10), .z(tmp00_10_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600011(.x(x_11), .z(tmp00_11_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600012(.x(x_12), .z(tmp00_12_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600013(.x(x_13), .z(tmp00_13_60));
	booth__002 #(.WIDTH(WIDTH)) mul00600014(.x(x_14), .z(tmp00_14_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600015(.x(x_15), .z(tmp00_15_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600016(.x(x_16), .z(tmp00_16_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600017(.x(x_17), .z(tmp00_17_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600018(.x(x_18), .z(tmp00_18_60));
	booth_0006 #(.WIDTH(WIDTH)) mul00600019(.x(x_19), .z(tmp00_19_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600020(.x(x_20), .z(tmp00_20_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600021(.x(x_21), .z(tmp00_21_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600022(.x(x_22), .z(tmp00_22_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600023(.x(x_23), .z(tmp00_23_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600024(.x(x_24), .z(tmp00_24_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600025(.x(x_25), .z(tmp00_25_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600026(.x(x_26), .z(tmp00_26_60));
	booth__002 #(.WIDTH(WIDTH)) mul00600027(.x(x_27), .z(tmp00_27_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600028(.x(x_28), .z(tmp00_28_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600029(.x(x_29), .z(tmp00_29_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600030(.x(x_30), .z(tmp00_30_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600031(.x(x_31), .z(tmp00_31_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600032(.x(x_32), .z(tmp00_32_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600033(.x(x_33), .z(tmp00_33_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600034(.x(x_34), .z(tmp00_34_60));
	booth__006 #(.WIDTH(WIDTH)) mul00600035(.x(x_35), .z(tmp00_35_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600036(.x(x_36), .z(tmp00_36_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600037(.x(x_37), .z(tmp00_37_60));
	booth_0010 #(.WIDTH(WIDTH)) mul00600038(.x(x_38), .z(tmp00_38_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600039(.x(x_39), .z(tmp00_39_60));
	booth__006 #(.WIDTH(WIDTH)) mul00600040(.x(x_40), .z(tmp00_40_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600041(.x(x_41), .z(tmp00_41_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600042(.x(x_42), .z(tmp00_42_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600043(.x(x_43), .z(tmp00_43_60));
	booth_0006 #(.WIDTH(WIDTH)) mul00600044(.x(x_44), .z(tmp00_44_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600045(.x(x_45), .z(tmp00_45_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600046(.x(x_46), .z(tmp00_46_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600047(.x(x_47), .z(tmp00_47_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600048(.x(x_48), .z(tmp00_48_60));
	booth_0010 #(.WIDTH(WIDTH)) mul00600049(.x(x_49), .z(tmp00_49_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600050(.x(x_50), .z(tmp00_50_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600051(.x(x_51), .z(tmp00_51_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600052(.x(x_52), .z(tmp00_52_60));
	booth__010 #(.WIDTH(WIDTH)) mul00600053(.x(x_53), .z(tmp00_53_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600054(.x(x_54), .z(tmp00_54_60));
	booth__010 #(.WIDTH(WIDTH)) mul00600055(.x(x_55), .z(tmp00_55_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600056(.x(x_56), .z(tmp00_56_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600057(.x(x_57), .z(tmp00_57_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600058(.x(x_58), .z(tmp00_58_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600059(.x(x_59), .z(tmp00_59_60));
	booth_0002 #(.WIDTH(WIDTH)) mul00600060(.x(x_60), .z(tmp00_60_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600061(.x(x_61), .z(tmp00_61_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600062(.x(x_62), .z(tmp00_62_60));
	booth__002 #(.WIDTH(WIDTH)) mul00600063(.x(x_63), .z(tmp00_63_60));
	booth__006 #(.WIDTH(WIDTH)) mul00600064(.x(x_64), .z(tmp00_64_60));
	booth_0010 #(.WIDTH(WIDTH)) mul00600065(.x(x_65), .z(tmp00_65_60));
	booth__006 #(.WIDTH(WIDTH)) mul00600066(.x(x_66), .z(tmp00_66_60));
	booth__006 #(.WIDTH(WIDTH)) mul00600067(.x(x_67), .z(tmp00_67_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600068(.x(x_68), .z(tmp00_68_60));
	booth__010 #(.WIDTH(WIDTH)) mul00600069(.x(x_69), .z(tmp00_69_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600070(.x(x_70), .z(tmp00_70_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600071(.x(x_71), .z(tmp00_71_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600072(.x(x_72), .z(tmp00_72_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600073(.x(x_73), .z(tmp00_73_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600074(.x(x_74), .z(tmp00_74_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600075(.x(x_75), .z(tmp00_75_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600076(.x(x_76), .z(tmp00_76_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600077(.x(x_77), .z(tmp00_77_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600078(.x(x_78), .z(tmp00_78_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600079(.x(x_79), .z(tmp00_79_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600080(.x(x_80), .z(tmp00_80_60));
	booth_0010 #(.WIDTH(WIDTH)) mul00600081(.x(x_81), .z(tmp00_81_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600082(.x(x_82), .z(tmp00_82_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600083(.x(x_83), .z(tmp00_83_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600084(.x(x_84), .z(tmp00_84_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600085(.x(x_85), .z(tmp00_85_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600086(.x(x_86), .z(tmp00_86_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600087(.x(x_87), .z(tmp00_87_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600088(.x(x_88), .z(tmp00_88_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600089(.x(x_89), .z(tmp00_89_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600090(.x(x_90), .z(tmp00_90_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600091(.x(x_91), .z(tmp00_91_60));
	booth__002 #(.WIDTH(WIDTH)) mul00600092(.x(x_92), .z(tmp00_92_60));
	booth__006 #(.WIDTH(WIDTH)) mul00600093(.x(x_93), .z(tmp00_93_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600094(.x(x_94), .z(tmp00_94_60));
	booth_0010 #(.WIDTH(WIDTH)) mul00600095(.x(x_95), .z(tmp00_95_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600096(.x(x_96), .z(tmp00_96_60));
	booth__002 #(.WIDTH(WIDTH)) mul00600097(.x(x_97), .z(tmp00_97_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600098(.x(x_98), .z(tmp00_98_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600099(.x(x_99), .z(tmp00_99_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600100(.x(x_100), .z(tmp00_100_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600101(.x(x_101), .z(tmp00_101_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600102(.x(x_102), .z(tmp00_102_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600103(.x(x_103), .z(tmp00_103_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600104(.x(x_104), .z(tmp00_104_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600105(.x(x_105), .z(tmp00_105_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600106(.x(x_106), .z(tmp00_106_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600107(.x(x_107), .z(tmp00_107_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600108(.x(x_108), .z(tmp00_108_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600109(.x(x_109), .z(tmp00_109_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600110(.x(x_110), .z(tmp00_110_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600111(.x(x_111), .z(tmp00_111_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600112(.x(x_112), .z(tmp00_112_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600113(.x(x_113), .z(tmp00_113_60));
	booth_0008 #(.WIDTH(WIDTH)) mul00600114(.x(x_114), .z(tmp00_114_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600115(.x(x_115), .z(tmp00_115_60));
	booth__002 #(.WIDTH(WIDTH)) mul00600116(.x(x_116), .z(tmp00_116_60));
	booth_0006 #(.WIDTH(WIDTH)) mul00600117(.x(x_117), .z(tmp00_117_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600118(.x(x_118), .z(tmp00_118_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600119(.x(x_119), .z(tmp00_119_60));
	booth__008 #(.WIDTH(WIDTH)) mul00600120(.x(x_120), .z(tmp00_120_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600121(.x(x_121), .z(tmp00_121_60));
	booth_0004 #(.WIDTH(WIDTH)) mul00600122(.x(x_122), .z(tmp00_122_60));
	booth__004 #(.WIDTH(WIDTH)) mul00600123(.x(x_123), .z(tmp00_123_60));
	booth_0002 #(.WIDTH(WIDTH)) mul00600124(.x(x_124), .z(tmp00_124_60));
	booth__010 #(.WIDTH(WIDTH)) mul00600125(.x(x_125), .z(tmp00_125_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600126(.x(x_126), .z(tmp00_126_60));
	booth_0000 #(.WIDTH(WIDTH)) mul00600127(.x(x_127), .z(tmp00_127_60));
	booth__004 #(.WIDTH(WIDTH)) mul00610000(.x(x_0), .z(tmp00_0_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610001(.x(x_1), .z(tmp00_1_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610002(.x(x_2), .z(tmp00_2_61));
	booth__010 #(.WIDTH(WIDTH)) mul00610003(.x(x_3), .z(tmp00_3_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610004(.x(x_4), .z(tmp00_4_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610005(.x(x_5), .z(tmp00_5_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610006(.x(x_6), .z(tmp00_6_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610007(.x(x_7), .z(tmp00_7_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610008(.x(x_8), .z(tmp00_8_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610009(.x(x_9), .z(tmp00_9_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610010(.x(x_10), .z(tmp00_10_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610011(.x(x_11), .z(tmp00_11_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610012(.x(x_12), .z(tmp00_12_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610013(.x(x_13), .z(tmp00_13_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610014(.x(x_14), .z(tmp00_14_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610015(.x(x_15), .z(tmp00_15_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610016(.x(x_16), .z(tmp00_16_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610017(.x(x_17), .z(tmp00_17_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610018(.x(x_18), .z(tmp00_18_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610019(.x(x_19), .z(tmp00_19_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610020(.x(x_20), .z(tmp00_20_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610021(.x(x_21), .z(tmp00_21_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610022(.x(x_22), .z(tmp00_22_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610023(.x(x_23), .z(tmp00_23_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610024(.x(x_24), .z(tmp00_24_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610025(.x(x_25), .z(tmp00_25_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610026(.x(x_26), .z(tmp00_26_61));
	booth__002 #(.WIDTH(WIDTH)) mul00610027(.x(x_27), .z(tmp00_27_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610028(.x(x_28), .z(tmp00_28_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610029(.x(x_29), .z(tmp00_29_61));
	booth__010 #(.WIDTH(WIDTH)) mul00610030(.x(x_30), .z(tmp00_30_61));
	booth_0012 #(.WIDTH(WIDTH)) mul00610031(.x(x_31), .z(tmp00_31_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610032(.x(x_32), .z(tmp00_32_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610033(.x(x_33), .z(tmp00_33_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610034(.x(x_34), .z(tmp00_34_61));
	booth__006 #(.WIDTH(WIDTH)) mul00610035(.x(x_35), .z(tmp00_35_61));
	booth__012 #(.WIDTH(WIDTH)) mul00610036(.x(x_36), .z(tmp00_36_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610037(.x(x_37), .z(tmp00_37_61));
	booth__002 #(.WIDTH(WIDTH)) mul00610038(.x(x_38), .z(tmp00_38_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610039(.x(x_39), .z(tmp00_39_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610040(.x(x_40), .z(tmp00_40_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610041(.x(x_41), .z(tmp00_41_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610042(.x(x_42), .z(tmp00_42_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610043(.x(x_43), .z(tmp00_43_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610044(.x(x_44), .z(tmp00_44_61));
	booth_0012 #(.WIDTH(WIDTH)) mul00610045(.x(x_45), .z(tmp00_45_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610046(.x(x_46), .z(tmp00_46_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610047(.x(x_47), .z(tmp00_47_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610048(.x(x_48), .z(tmp00_48_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610049(.x(x_49), .z(tmp00_49_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610050(.x(x_50), .z(tmp00_50_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610051(.x(x_51), .z(tmp00_51_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610052(.x(x_52), .z(tmp00_52_61));
	booth_0006 #(.WIDTH(WIDTH)) mul00610053(.x(x_53), .z(tmp00_53_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610054(.x(x_54), .z(tmp00_54_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610055(.x(x_55), .z(tmp00_55_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610056(.x(x_56), .z(tmp00_56_61));
	booth__006 #(.WIDTH(WIDTH)) mul00610057(.x(x_57), .z(tmp00_57_61));
	booth__002 #(.WIDTH(WIDTH)) mul00610058(.x(x_58), .z(tmp00_58_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610059(.x(x_59), .z(tmp00_59_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610060(.x(x_60), .z(tmp00_60_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610061(.x(x_61), .z(tmp00_61_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610062(.x(x_62), .z(tmp00_62_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610063(.x(x_63), .z(tmp00_63_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610064(.x(x_64), .z(tmp00_64_61));
	booth__010 #(.WIDTH(WIDTH)) mul00610065(.x(x_65), .z(tmp00_65_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610066(.x(x_66), .z(tmp00_66_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610067(.x(x_67), .z(tmp00_67_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610068(.x(x_68), .z(tmp00_68_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610069(.x(x_69), .z(tmp00_69_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610070(.x(x_70), .z(tmp00_70_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610071(.x(x_71), .z(tmp00_71_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610072(.x(x_72), .z(tmp00_72_61));
	booth_0010 #(.WIDTH(WIDTH)) mul00610073(.x(x_73), .z(tmp00_73_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610074(.x(x_74), .z(tmp00_74_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610075(.x(x_75), .z(tmp00_75_61));
	booth_0010 #(.WIDTH(WIDTH)) mul00610076(.x(x_76), .z(tmp00_76_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610077(.x(x_77), .z(tmp00_77_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610078(.x(x_78), .z(tmp00_78_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610079(.x(x_79), .z(tmp00_79_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610080(.x(x_80), .z(tmp00_80_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610081(.x(x_81), .z(tmp00_81_61));
	booth_0006 #(.WIDTH(WIDTH)) mul00610082(.x(x_82), .z(tmp00_82_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610083(.x(x_83), .z(tmp00_83_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610084(.x(x_84), .z(tmp00_84_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610085(.x(x_85), .z(tmp00_85_61));
	booth_0006 #(.WIDTH(WIDTH)) mul00610086(.x(x_86), .z(tmp00_86_61));
	booth__002 #(.WIDTH(WIDTH)) mul00610087(.x(x_87), .z(tmp00_87_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610088(.x(x_88), .z(tmp00_88_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610089(.x(x_89), .z(tmp00_89_61));
	booth__012 #(.WIDTH(WIDTH)) mul00610090(.x(x_90), .z(tmp00_90_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610091(.x(x_91), .z(tmp00_91_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610092(.x(x_92), .z(tmp00_92_61));
	booth__010 #(.WIDTH(WIDTH)) mul00610093(.x(x_93), .z(tmp00_93_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610094(.x(x_94), .z(tmp00_94_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610095(.x(x_95), .z(tmp00_95_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610096(.x(x_96), .z(tmp00_96_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610097(.x(x_97), .z(tmp00_97_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610098(.x(x_98), .z(tmp00_98_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610099(.x(x_99), .z(tmp00_99_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610100(.x(x_100), .z(tmp00_100_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610101(.x(x_101), .z(tmp00_101_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610102(.x(x_102), .z(tmp00_102_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00610103(.x(x_103), .z(tmp00_103_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610104(.x(x_104), .z(tmp00_104_61));
	booth__006 #(.WIDTH(WIDTH)) mul00610105(.x(x_105), .z(tmp00_105_61));
	booth_0012 #(.WIDTH(WIDTH)) mul00610106(.x(x_106), .z(tmp00_106_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610107(.x(x_107), .z(tmp00_107_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610108(.x(x_108), .z(tmp00_108_61));
	booth_0012 #(.WIDTH(WIDTH)) mul00610109(.x(x_109), .z(tmp00_109_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610110(.x(x_110), .z(tmp00_110_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610111(.x(x_111), .z(tmp00_111_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610112(.x(x_112), .z(tmp00_112_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610113(.x(x_113), .z(tmp00_113_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610114(.x(x_114), .z(tmp00_114_61));
	booth__010 #(.WIDTH(WIDTH)) mul00610115(.x(x_115), .z(tmp00_115_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610116(.x(x_116), .z(tmp00_116_61));
	booth__008 #(.WIDTH(WIDTH)) mul00610117(.x(x_117), .z(tmp00_117_61));
	booth_0004 #(.WIDTH(WIDTH)) mul00610118(.x(x_118), .z(tmp00_118_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610119(.x(x_119), .z(tmp00_119_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610120(.x(x_120), .z(tmp00_120_61));
	booth__002 #(.WIDTH(WIDTH)) mul00610121(.x(x_121), .z(tmp00_121_61));
	booth__004 #(.WIDTH(WIDTH)) mul00610122(.x(x_122), .z(tmp00_122_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610123(.x(x_123), .z(tmp00_123_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610124(.x(x_124), .z(tmp00_124_61));
	booth_0008 #(.WIDTH(WIDTH)) mul00610125(.x(x_125), .z(tmp00_125_61));
	booth__006 #(.WIDTH(WIDTH)) mul00610126(.x(x_126), .z(tmp00_126_61));
	booth_0000 #(.WIDTH(WIDTH)) mul00610127(.x(x_127), .z(tmp00_127_61));
	booth_0002 #(.WIDTH(WIDTH)) mul00620000(.x(x_0), .z(tmp00_0_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620001(.x(x_1), .z(tmp00_1_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620002(.x(x_2), .z(tmp00_2_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620003(.x(x_3), .z(tmp00_3_62));
	booth__014 #(.WIDTH(WIDTH)) mul00620004(.x(x_4), .z(tmp00_4_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620005(.x(x_5), .z(tmp00_5_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620006(.x(x_6), .z(tmp00_6_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620007(.x(x_7), .z(tmp00_7_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620008(.x(x_8), .z(tmp00_8_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620009(.x(x_9), .z(tmp00_9_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620010(.x(x_10), .z(tmp00_10_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620011(.x(x_11), .z(tmp00_11_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620012(.x(x_12), .z(tmp00_12_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620013(.x(x_13), .z(tmp00_13_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620014(.x(x_14), .z(tmp00_14_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620015(.x(x_15), .z(tmp00_15_62));
	booth_0010 #(.WIDTH(WIDTH)) mul00620016(.x(x_16), .z(tmp00_16_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620017(.x(x_17), .z(tmp00_17_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620018(.x(x_18), .z(tmp00_18_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620019(.x(x_19), .z(tmp00_19_62));
	booth_0006 #(.WIDTH(WIDTH)) mul00620020(.x(x_20), .z(tmp00_20_62));
	booth_0002 #(.WIDTH(WIDTH)) mul00620021(.x(x_21), .z(tmp00_21_62));
	booth_0010 #(.WIDTH(WIDTH)) mul00620022(.x(x_22), .z(tmp00_22_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620023(.x(x_23), .z(tmp00_23_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620024(.x(x_24), .z(tmp00_24_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620025(.x(x_25), .z(tmp00_25_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620026(.x(x_26), .z(tmp00_26_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620027(.x(x_27), .z(tmp00_27_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620028(.x(x_28), .z(tmp00_28_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620029(.x(x_29), .z(tmp00_29_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620030(.x(x_30), .z(tmp00_30_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620031(.x(x_31), .z(tmp00_31_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620032(.x(x_32), .z(tmp00_32_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620033(.x(x_33), .z(tmp00_33_62));
	booth__006 #(.WIDTH(WIDTH)) mul00620034(.x(x_34), .z(tmp00_34_62));
	booth_0012 #(.WIDTH(WIDTH)) mul00620035(.x(x_35), .z(tmp00_35_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620036(.x(x_36), .z(tmp00_36_62));
	booth_0006 #(.WIDTH(WIDTH)) mul00620037(.x(x_37), .z(tmp00_37_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620038(.x(x_38), .z(tmp00_38_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620039(.x(x_39), .z(tmp00_39_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620040(.x(x_40), .z(tmp00_40_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620041(.x(x_41), .z(tmp00_41_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620042(.x(x_42), .z(tmp00_42_62));
	booth__010 #(.WIDTH(WIDTH)) mul00620043(.x(x_43), .z(tmp00_43_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620044(.x(x_44), .z(tmp00_44_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620045(.x(x_45), .z(tmp00_45_62));
	booth_0010 #(.WIDTH(WIDTH)) mul00620046(.x(x_46), .z(tmp00_46_62));
	booth_0002 #(.WIDTH(WIDTH)) mul00620047(.x(x_47), .z(tmp00_47_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620048(.x(x_48), .z(tmp00_48_62));
	booth_0006 #(.WIDTH(WIDTH)) mul00620049(.x(x_49), .z(tmp00_49_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620050(.x(x_50), .z(tmp00_50_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620051(.x(x_51), .z(tmp00_51_62));
	booth_0012 #(.WIDTH(WIDTH)) mul00620052(.x(x_52), .z(tmp00_52_62));
	booth_0002 #(.WIDTH(WIDTH)) mul00620053(.x(x_53), .z(tmp00_53_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620054(.x(x_54), .z(tmp00_54_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620055(.x(x_55), .z(tmp00_55_62));
	booth_0012 #(.WIDTH(WIDTH)) mul00620056(.x(x_56), .z(tmp00_56_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620057(.x(x_57), .z(tmp00_57_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620058(.x(x_58), .z(tmp00_58_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620059(.x(x_59), .z(tmp00_59_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620060(.x(x_60), .z(tmp00_60_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620061(.x(x_61), .z(tmp00_61_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620062(.x(x_62), .z(tmp00_62_62));
	booth_0006 #(.WIDTH(WIDTH)) mul00620063(.x(x_63), .z(tmp00_63_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620064(.x(x_64), .z(tmp00_64_62));
	booth__002 #(.WIDTH(WIDTH)) mul00620065(.x(x_65), .z(tmp00_65_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620066(.x(x_66), .z(tmp00_66_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620067(.x(x_67), .z(tmp00_67_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620068(.x(x_68), .z(tmp00_68_62));
	booth__012 #(.WIDTH(WIDTH)) mul00620069(.x(x_69), .z(tmp00_69_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620070(.x(x_70), .z(tmp00_70_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620071(.x(x_71), .z(tmp00_71_62));
	booth__002 #(.WIDTH(WIDTH)) mul00620072(.x(x_72), .z(tmp00_72_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620073(.x(x_73), .z(tmp00_73_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620074(.x(x_74), .z(tmp00_74_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620075(.x(x_75), .z(tmp00_75_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620076(.x(x_76), .z(tmp00_76_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620077(.x(x_77), .z(tmp00_77_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620078(.x(x_78), .z(tmp00_78_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620079(.x(x_79), .z(tmp00_79_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620080(.x(x_80), .z(tmp00_80_62));
	booth_0010 #(.WIDTH(WIDTH)) mul00620081(.x(x_81), .z(tmp00_81_62));
	booth__012 #(.WIDTH(WIDTH)) mul00620082(.x(x_82), .z(tmp00_82_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620083(.x(x_83), .z(tmp00_83_62));
	booth__006 #(.WIDTH(WIDTH)) mul00620084(.x(x_84), .z(tmp00_84_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620085(.x(x_85), .z(tmp00_85_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620086(.x(x_86), .z(tmp00_86_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620087(.x(x_87), .z(tmp00_87_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620088(.x(x_88), .z(tmp00_88_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620089(.x(x_89), .z(tmp00_89_62));
	booth_0012 #(.WIDTH(WIDTH)) mul00620090(.x(x_90), .z(tmp00_90_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620091(.x(x_91), .z(tmp00_91_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620092(.x(x_92), .z(tmp00_92_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620093(.x(x_93), .z(tmp00_93_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620094(.x(x_94), .z(tmp00_94_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620095(.x(x_95), .z(tmp00_95_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620096(.x(x_96), .z(tmp00_96_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620097(.x(x_97), .z(tmp00_97_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620098(.x(x_98), .z(tmp00_98_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620099(.x(x_99), .z(tmp00_99_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620100(.x(x_100), .z(tmp00_100_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620101(.x(x_101), .z(tmp00_101_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620102(.x(x_102), .z(tmp00_102_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620103(.x(x_103), .z(tmp00_103_62));
	booth__002 #(.WIDTH(WIDTH)) mul00620104(.x(x_104), .z(tmp00_104_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620105(.x(x_105), .z(tmp00_105_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620106(.x(x_106), .z(tmp00_106_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620107(.x(x_107), .z(tmp00_107_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620108(.x(x_108), .z(tmp00_108_62));
	booth__012 #(.WIDTH(WIDTH)) mul00620109(.x(x_109), .z(tmp00_109_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620110(.x(x_110), .z(tmp00_110_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620111(.x(x_111), .z(tmp00_111_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620112(.x(x_112), .z(tmp00_112_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620113(.x(x_113), .z(tmp00_113_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620114(.x(x_114), .z(tmp00_114_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620115(.x(x_115), .z(tmp00_115_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620116(.x(x_116), .z(tmp00_116_62));
	booth_0004 #(.WIDTH(WIDTH)) mul00620117(.x(x_117), .z(tmp00_117_62));
	booth_0000 #(.WIDTH(WIDTH)) mul00620118(.x(x_118), .z(tmp00_118_62));
	booth_0006 #(.WIDTH(WIDTH)) mul00620119(.x(x_119), .z(tmp00_119_62));
	booth__008 #(.WIDTH(WIDTH)) mul00620120(.x(x_120), .z(tmp00_120_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620121(.x(x_121), .z(tmp00_121_62));
	booth__002 #(.WIDTH(WIDTH)) mul00620122(.x(x_122), .z(tmp00_122_62));
	booth__004 #(.WIDTH(WIDTH)) mul00620123(.x(x_123), .z(tmp00_123_62));
	booth__010 #(.WIDTH(WIDTH)) mul00620124(.x(x_124), .z(tmp00_124_62));
	booth_0008 #(.WIDTH(WIDTH)) mul00620125(.x(x_125), .z(tmp00_125_62));
	booth_0006 #(.WIDTH(WIDTH)) mul00620126(.x(x_126), .z(tmp00_126_62));
	booth__006 #(.WIDTH(WIDTH)) mul00620127(.x(x_127), .z(tmp00_127_62));
	booth_0006 #(.WIDTH(WIDTH)) mul00630000(.x(x_0), .z(tmp00_0_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630001(.x(x_1), .z(tmp00_1_63));
	booth__010 #(.WIDTH(WIDTH)) mul00630002(.x(x_2), .z(tmp00_2_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630003(.x(x_3), .z(tmp00_3_63));
	booth__016 #(.WIDTH(WIDTH)) mul00630004(.x(x_4), .z(tmp00_4_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630005(.x(x_5), .z(tmp00_5_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630006(.x(x_6), .z(tmp00_6_63));
	booth_0010 #(.WIDTH(WIDTH)) mul00630007(.x(x_7), .z(tmp00_7_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630008(.x(x_8), .z(tmp00_8_63));
	booth_0006 #(.WIDTH(WIDTH)) mul00630009(.x(x_9), .z(tmp00_9_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630010(.x(x_10), .z(tmp00_10_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630011(.x(x_11), .z(tmp00_11_63));
	booth__008 #(.WIDTH(WIDTH)) mul00630012(.x(x_12), .z(tmp00_12_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630013(.x(x_13), .z(tmp00_13_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630014(.x(x_14), .z(tmp00_14_63));
	booth__008 #(.WIDTH(WIDTH)) mul00630015(.x(x_15), .z(tmp00_15_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630016(.x(x_16), .z(tmp00_16_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630017(.x(x_17), .z(tmp00_17_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630018(.x(x_18), .z(tmp00_18_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630019(.x(x_19), .z(tmp00_19_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630020(.x(x_20), .z(tmp00_20_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630021(.x(x_21), .z(tmp00_21_63));
	booth_0016 #(.WIDTH(WIDTH)) mul00630022(.x(x_22), .z(tmp00_22_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630023(.x(x_23), .z(tmp00_23_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630024(.x(x_24), .z(tmp00_24_63));
	booth_0012 #(.WIDTH(WIDTH)) mul00630025(.x(x_25), .z(tmp00_25_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630026(.x(x_26), .z(tmp00_26_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630027(.x(x_27), .z(tmp00_27_63));
	booth_0002 #(.WIDTH(WIDTH)) mul00630028(.x(x_28), .z(tmp00_28_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630029(.x(x_29), .z(tmp00_29_63));
	booth_0006 #(.WIDTH(WIDTH)) mul00630030(.x(x_30), .z(tmp00_30_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630031(.x(x_31), .z(tmp00_31_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630032(.x(x_32), .z(tmp00_32_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630033(.x(x_33), .z(tmp00_33_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630034(.x(x_34), .z(tmp00_34_63));
	booth_0002 #(.WIDTH(WIDTH)) mul00630035(.x(x_35), .z(tmp00_35_63));
	booth__006 #(.WIDTH(WIDTH)) mul00630036(.x(x_36), .z(tmp00_36_63));
	booth__006 #(.WIDTH(WIDTH)) mul00630037(.x(x_37), .z(tmp00_37_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630038(.x(x_38), .z(tmp00_38_63));
	booth_0016 #(.WIDTH(WIDTH)) mul00630039(.x(x_39), .z(tmp00_39_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630040(.x(x_40), .z(tmp00_40_63));
	booth__012 #(.WIDTH(WIDTH)) mul00630041(.x(x_41), .z(tmp00_41_63));
	booth__008 #(.WIDTH(WIDTH)) mul00630042(.x(x_42), .z(tmp00_42_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630043(.x(x_43), .z(tmp00_43_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630044(.x(x_44), .z(tmp00_44_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630045(.x(x_45), .z(tmp00_45_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630046(.x(x_46), .z(tmp00_46_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630047(.x(x_47), .z(tmp00_47_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630048(.x(x_48), .z(tmp00_48_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630049(.x(x_49), .z(tmp00_49_63));
	booth_0012 #(.WIDTH(WIDTH)) mul00630050(.x(x_50), .z(tmp00_50_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630051(.x(x_51), .z(tmp00_51_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630052(.x(x_52), .z(tmp00_52_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630053(.x(x_53), .z(tmp00_53_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630054(.x(x_54), .z(tmp00_54_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630055(.x(x_55), .z(tmp00_55_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630056(.x(x_56), .z(tmp00_56_63));
	booth_0002 #(.WIDTH(WIDTH)) mul00630057(.x(x_57), .z(tmp00_57_63));
	booth__008 #(.WIDTH(WIDTH)) mul00630058(.x(x_58), .z(tmp00_58_63));
	booth_0014 #(.WIDTH(WIDTH)) mul00630059(.x(x_59), .z(tmp00_59_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630060(.x(x_60), .z(tmp00_60_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630061(.x(x_61), .z(tmp00_61_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630062(.x(x_62), .z(tmp00_62_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630063(.x(x_63), .z(tmp00_63_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630064(.x(x_64), .z(tmp00_64_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630065(.x(x_65), .z(tmp00_65_63));
	booth__008 #(.WIDTH(WIDTH)) mul00630066(.x(x_66), .z(tmp00_66_63));
	booth__006 #(.WIDTH(WIDTH)) mul00630067(.x(x_67), .z(tmp00_67_63));
	booth_0012 #(.WIDTH(WIDTH)) mul00630068(.x(x_68), .z(tmp00_68_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630069(.x(x_69), .z(tmp00_69_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630070(.x(x_70), .z(tmp00_70_63));
	booth_0002 #(.WIDTH(WIDTH)) mul00630071(.x(x_71), .z(tmp00_71_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630072(.x(x_72), .z(tmp00_72_63));
	booth__008 #(.WIDTH(WIDTH)) mul00630073(.x(x_73), .z(tmp00_73_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630074(.x(x_74), .z(tmp00_74_63));
	booth_0010 #(.WIDTH(WIDTH)) mul00630075(.x(x_75), .z(tmp00_75_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630076(.x(x_76), .z(tmp00_76_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630077(.x(x_77), .z(tmp00_77_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630078(.x(x_78), .z(tmp00_78_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630079(.x(x_79), .z(tmp00_79_63));
	booth_0010 #(.WIDTH(WIDTH)) mul00630080(.x(x_80), .z(tmp00_80_63));
	booth__008 #(.WIDTH(WIDTH)) mul00630081(.x(x_81), .z(tmp00_81_63));
	booth__006 #(.WIDTH(WIDTH)) mul00630082(.x(x_82), .z(tmp00_82_63));
	booth_0006 #(.WIDTH(WIDTH)) mul00630083(.x(x_83), .z(tmp00_83_63));
	booth_0006 #(.WIDTH(WIDTH)) mul00630084(.x(x_84), .z(tmp00_84_63));
	booth_0006 #(.WIDTH(WIDTH)) mul00630085(.x(x_85), .z(tmp00_85_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630086(.x(x_86), .z(tmp00_86_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630087(.x(x_87), .z(tmp00_87_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630088(.x(x_88), .z(tmp00_88_63));
	booth_0006 #(.WIDTH(WIDTH)) mul00630089(.x(x_89), .z(tmp00_89_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630090(.x(x_90), .z(tmp00_90_63));
	booth__006 #(.WIDTH(WIDTH)) mul00630091(.x(x_91), .z(tmp00_91_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630092(.x(x_92), .z(tmp00_92_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630093(.x(x_93), .z(tmp00_93_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630094(.x(x_94), .z(tmp00_94_63));
	booth__012 #(.WIDTH(WIDTH)) mul00630095(.x(x_95), .z(tmp00_95_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630096(.x(x_96), .z(tmp00_96_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630097(.x(x_97), .z(tmp00_97_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630098(.x(x_98), .z(tmp00_98_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630099(.x(x_99), .z(tmp00_99_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630100(.x(x_100), .z(tmp00_100_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630101(.x(x_101), .z(tmp00_101_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630102(.x(x_102), .z(tmp00_102_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630103(.x(x_103), .z(tmp00_103_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630104(.x(x_104), .z(tmp00_104_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630105(.x(x_105), .z(tmp00_105_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630106(.x(x_106), .z(tmp00_106_63));
	booth__010 #(.WIDTH(WIDTH)) mul00630107(.x(x_107), .z(tmp00_107_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630108(.x(x_108), .z(tmp00_108_63));
	booth__002 #(.WIDTH(WIDTH)) mul00630109(.x(x_109), .z(tmp00_109_63));
	booth_0002 #(.WIDTH(WIDTH)) mul00630110(.x(x_110), .z(tmp00_110_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630111(.x(x_111), .z(tmp00_111_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630112(.x(x_112), .z(tmp00_112_63));
	booth_0016 #(.WIDTH(WIDTH)) mul00630113(.x(x_113), .z(tmp00_113_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630114(.x(x_114), .z(tmp00_114_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630115(.x(x_115), .z(tmp00_115_63));
	booth_0008 #(.WIDTH(WIDTH)) mul00630116(.x(x_116), .z(tmp00_116_63));
	booth_0012 #(.WIDTH(WIDTH)) mul00630117(.x(x_117), .z(tmp00_117_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630118(.x(x_118), .z(tmp00_118_63));
	booth__004 #(.WIDTH(WIDTH)) mul00630119(.x(x_119), .z(tmp00_119_63));
	booth_0012 #(.WIDTH(WIDTH)) mul00630120(.x(x_120), .z(tmp00_120_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630121(.x(x_121), .z(tmp00_121_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630122(.x(x_122), .z(tmp00_122_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630123(.x(x_123), .z(tmp00_123_63));
	booth_0004 #(.WIDTH(WIDTH)) mul00630124(.x(x_124), .z(tmp00_124_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630125(.x(x_125), .z(tmp00_125_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00630126(.x(x_126), .z(tmp00_126_63));
	booth_0006 #(.WIDTH(WIDTH)) mul00630127(.x(x_127), .z(tmp00_127_63));
	booth_0000 #(.WIDTH(WIDTH)) mul00640000(.x(x_0), .z(tmp00_0_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640001(.x(x_1), .z(tmp00_1_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640002(.x(x_2), .z(tmp00_2_64));
	booth__010 #(.WIDTH(WIDTH)) mul00640003(.x(x_3), .z(tmp00_3_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640004(.x(x_4), .z(tmp00_4_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640005(.x(x_5), .z(tmp00_5_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640006(.x(x_6), .z(tmp00_6_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640007(.x(x_7), .z(tmp00_7_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640008(.x(x_8), .z(tmp00_8_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640009(.x(x_9), .z(tmp00_9_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640010(.x(x_10), .z(tmp00_10_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640011(.x(x_11), .z(tmp00_11_64));
	booth__010 #(.WIDTH(WIDTH)) mul00640012(.x(x_12), .z(tmp00_12_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640013(.x(x_13), .z(tmp00_13_64));
	booth__004 #(.WIDTH(WIDTH)) mul00640014(.x(x_14), .z(tmp00_14_64));
	booth_0012 #(.WIDTH(WIDTH)) mul00640015(.x(x_15), .z(tmp00_15_64));
	booth__006 #(.WIDTH(WIDTH)) mul00640016(.x(x_16), .z(tmp00_16_64));
	booth__014 #(.WIDTH(WIDTH)) mul00640017(.x(x_17), .z(tmp00_17_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640018(.x(x_18), .z(tmp00_18_64));
	booth__002 #(.WIDTH(WIDTH)) mul00640019(.x(x_19), .z(tmp00_19_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640020(.x(x_20), .z(tmp00_20_64));
	booth__006 #(.WIDTH(WIDTH)) mul00640021(.x(x_21), .z(tmp00_21_64));
	booth__006 #(.WIDTH(WIDTH)) mul00640022(.x(x_22), .z(tmp00_22_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640023(.x(x_23), .z(tmp00_23_64));
	booth_0002 #(.WIDTH(WIDTH)) mul00640024(.x(x_24), .z(tmp00_24_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640025(.x(x_25), .z(tmp00_25_64));
	booth__002 #(.WIDTH(WIDTH)) mul00640026(.x(x_26), .z(tmp00_26_64));
	booth__006 #(.WIDTH(WIDTH)) mul00640027(.x(x_27), .z(tmp00_27_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640028(.x(x_28), .z(tmp00_28_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640029(.x(x_29), .z(tmp00_29_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640030(.x(x_30), .z(tmp00_30_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640031(.x(x_31), .z(tmp00_31_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640032(.x(x_32), .z(tmp00_32_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640033(.x(x_33), .z(tmp00_33_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640034(.x(x_34), .z(tmp00_34_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640035(.x(x_35), .z(tmp00_35_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640036(.x(x_36), .z(tmp00_36_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640037(.x(x_37), .z(tmp00_37_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640038(.x(x_38), .z(tmp00_38_64));
	booth__018 #(.WIDTH(WIDTH)) mul00640039(.x(x_39), .z(tmp00_39_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640040(.x(x_40), .z(tmp00_40_64));
	booth_0012 #(.WIDTH(WIDTH)) mul00640041(.x(x_41), .z(tmp00_41_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640042(.x(x_42), .z(tmp00_42_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640043(.x(x_43), .z(tmp00_43_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640044(.x(x_44), .z(tmp00_44_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640045(.x(x_45), .z(tmp00_45_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640046(.x(x_46), .z(tmp00_46_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640047(.x(x_47), .z(tmp00_47_64));
	booth__012 #(.WIDTH(WIDTH)) mul00640048(.x(x_48), .z(tmp00_48_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640049(.x(x_49), .z(tmp00_49_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640050(.x(x_50), .z(tmp00_50_64));
	booth_0002 #(.WIDTH(WIDTH)) mul00640051(.x(x_51), .z(tmp00_51_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640052(.x(x_52), .z(tmp00_52_64));
	booth__004 #(.WIDTH(WIDTH)) mul00640053(.x(x_53), .z(tmp00_53_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640054(.x(x_54), .z(tmp00_54_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640055(.x(x_55), .z(tmp00_55_64));
	booth__002 #(.WIDTH(WIDTH)) mul00640056(.x(x_56), .z(tmp00_56_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640057(.x(x_57), .z(tmp00_57_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640058(.x(x_58), .z(tmp00_58_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640059(.x(x_59), .z(tmp00_59_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640060(.x(x_60), .z(tmp00_60_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640061(.x(x_61), .z(tmp00_61_64));
	booth__002 #(.WIDTH(WIDTH)) mul00640062(.x(x_62), .z(tmp00_62_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640063(.x(x_63), .z(tmp00_63_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640064(.x(x_64), .z(tmp00_64_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640065(.x(x_65), .z(tmp00_65_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640066(.x(x_66), .z(tmp00_66_64));
	booth_0006 #(.WIDTH(WIDTH)) mul00640067(.x(x_67), .z(tmp00_67_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640068(.x(x_68), .z(tmp00_68_64));
	booth__002 #(.WIDTH(WIDTH)) mul00640069(.x(x_69), .z(tmp00_69_64));
	booth_0002 #(.WIDTH(WIDTH)) mul00640070(.x(x_70), .z(tmp00_70_64));
	booth__006 #(.WIDTH(WIDTH)) mul00640071(.x(x_71), .z(tmp00_71_64));
	booth_0010 #(.WIDTH(WIDTH)) mul00640072(.x(x_72), .z(tmp00_72_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640073(.x(x_73), .z(tmp00_73_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640074(.x(x_74), .z(tmp00_74_64));
	booth__012 #(.WIDTH(WIDTH)) mul00640075(.x(x_75), .z(tmp00_75_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640076(.x(x_76), .z(tmp00_76_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640077(.x(x_77), .z(tmp00_77_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640078(.x(x_78), .z(tmp00_78_64));
	booth__004 #(.WIDTH(WIDTH)) mul00640079(.x(x_79), .z(tmp00_79_64));
	booth_0002 #(.WIDTH(WIDTH)) mul00640080(.x(x_80), .z(tmp00_80_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640081(.x(x_81), .z(tmp00_81_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640082(.x(x_82), .z(tmp00_82_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640083(.x(x_83), .z(tmp00_83_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640084(.x(x_84), .z(tmp00_84_64));
	booth__012 #(.WIDTH(WIDTH)) mul00640085(.x(x_85), .z(tmp00_85_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640086(.x(x_86), .z(tmp00_86_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640087(.x(x_87), .z(tmp00_87_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640088(.x(x_88), .z(tmp00_88_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640089(.x(x_89), .z(tmp00_89_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640090(.x(x_90), .z(tmp00_90_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640091(.x(x_91), .z(tmp00_91_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640092(.x(x_92), .z(tmp00_92_64));
	booth__006 #(.WIDTH(WIDTH)) mul00640093(.x(x_93), .z(tmp00_93_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640094(.x(x_94), .z(tmp00_94_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640095(.x(x_95), .z(tmp00_95_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640096(.x(x_96), .z(tmp00_96_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640097(.x(x_97), .z(tmp00_97_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640098(.x(x_98), .z(tmp00_98_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640099(.x(x_99), .z(tmp00_99_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640100(.x(x_100), .z(tmp00_100_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640101(.x(x_101), .z(tmp00_101_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640102(.x(x_102), .z(tmp00_102_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640103(.x(x_103), .z(tmp00_103_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640104(.x(x_104), .z(tmp00_104_64));
	booth__006 #(.WIDTH(WIDTH)) mul00640105(.x(x_105), .z(tmp00_105_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640106(.x(x_106), .z(tmp00_106_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640107(.x(x_107), .z(tmp00_107_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640108(.x(x_108), .z(tmp00_108_64));
	booth__004 #(.WIDTH(WIDTH)) mul00640109(.x(x_109), .z(tmp00_109_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640110(.x(x_110), .z(tmp00_110_64));
	booth_0002 #(.WIDTH(WIDTH)) mul00640111(.x(x_111), .z(tmp00_111_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640112(.x(x_112), .z(tmp00_112_64));
	booth__004 #(.WIDTH(WIDTH)) mul00640113(.x(x_113), .z(tmp00_113_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640114(.x(x_114), .z(tmp00_114_64));
	booth_0002 #(.WIDTH(WIDTH)) mul00640115(.x(x_115), .z(tmp00_115_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640116(.x(x_116), .z(tmp00_116_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640117(.x(x_117), .z(tmp00_117_64));
	booth__008 #(.WIDTH(WIDTH)) mul00640118(.x(x_118), .z(tmp00_118_64));
	booth_0016 #(.WIDTH(WIDTH)) mul00640119(.x(x_119), .z(tmp00_119_64));
	booth__012 #(.WIDTH(WIDTH)) mul00640120(.x(x_120), .z(tmp00_120_64));
	booth_0008 #(.WIDTH(WIDTH)) mul00640121(.x(x_121), .z(tmp00_121_64));
	booth_0000 #(.WIDTH(WIDTH)) mul00640122(.x(x_122), .z(tmp00_122_64));
	booth__010 #(.WIDTH(WIDTH)) mul00640123(.x(x_123), .z(tmp00_123_64));
	booth__004 #(.WIDTH(WIDTH)) mul00640124(.x(x_124), .z(tmp00_124_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640125(.x(x_125), .z(tmp00_125_64));
	booth_0006 #(.WIDTH(WIDTH)) mul00640126(.x(x_126), .z(tmp00_126_64));
	booth_0004 #(.WIDTH(WIDTH)) mul00640127(.x(x_127), .z(tmp00_127_64));
	booth__004 #(.WIDTH(WIDTH)) mul00650000(.x(x_0), .z(tmp00_0_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650001(.x(x_1), .z(tmp00_1_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650002(.x(x_2), .z(tmp00_2_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650003(.x(x_3), .z(tmp00_3_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650004(.x(x_4), .z(tmp00_4_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650005(.x(x_5), .z(tmp00_5_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650006(.x(x_6), .z(tmp00_6_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650007(.x(x_7), .z(tmp00_7_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650008(.x(x_8), .z(tmp00_8_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650009(.x(x_9), .z(tmp00_9_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650010(.x(x_10), .z(tmp00_10_65));
	booth__002 #(.WIDTH(WIDTH)) mul00650011(.x(x_11), .z(tmp00_11_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650012(.x(x_12), .z(tmp00_12_65));
	booth_0010 #(.WIDTH(WIDTH)) mul00650013(.x(x_13), .z(tmp00_13_65));
	booth__010 #(.WIDTH(WIDTH)) mul00650014(.x(x_14), .z(tmp00_14_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650015(.x(x_15), .z(tmp00_15_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650016(.x(x_16), .z(tmp00_16_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650017(.x(x_17), .z(tmp00_17_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650018(.x(x_18), .z(tmp00_18_65));
	booth_0010 #(.WIDTH(WIDTH)) mul00650019(.x(x_19), .z(tmp00_19_65));
	booth__010 #(.WIDTH(WIDTH)) mul00650020(.x(x_20), .z(tmp00_20_65));
	booth_0010 #(.WIDTH(WIDTH)) mul00650021(.x(x_21), .z(tmp00_21_65));
	booth_0010 #(.WIDTH(WIDTH)) mul00650022(.x(x_22), .z(tmp00_22_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650023(.x(x_23), .z(tmp00_23_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650024(.x(x_24), .z(tmp00_24_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650025(.x(x_25), .z(tmp00_25_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650026(.x(x_26), .z(tmp00_26_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650027(.x(x_27), .z(tmp00_27_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650028(.x(x_28), .z(tmp00_28_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650029(.x(x_29), .z(tmp00_29_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650030(.x(x_30), .z(tmp00_30_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650031(.x(x_31), .z(tmp00_31_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650032(.x(x_32), .z(tmp00_32_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650033(.x(x_33), .z(tmp00_33_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650034(.x(x_34), .z(tmp00_34_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650035(.x(x_35), .z(tmp00_35_65));
	booth__006 #(.WIDTH(WIDTH)) mul00650036(.x(x_36), .z(tmp00_36_65));
	booth_0010 #(.WIDTH(WIDTH)) mul00650037(.x(x_37), .z(tmp00_37_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650038(.x(x_38), .z(tmp00_38_65));
	booth__006 #(.WIDTH(WIDTH)) mul00650039(.x(x_39), .z(tmp00_39_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650040(.x(x_40), .z(tmp00_40_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650041(.x(x_41), .z(tmp00_41_65));
	booth__010 #(.WIDTH(WIDTH)) mul00650042(.x(x_42), .z(tmp00_42_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650043(.x(x_43), .z(tmp00_43_65));
	booth_0006 #(.WIDTH(WIDTH)) mul00650044(.x(x_44), .z(tmp00_44_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650045(.x(x_45), .z(tmp00_45_65));
	booth__006 #(.WIDTH(WIDTH)) mul00650046(.x(x_46), .z(tmp00_46_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650047(.x(x_47), .z(tmp00_47_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650048(.x(x_48), .z(tmp00_48_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650049(.x(x_49), .z(tmp00_49_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650050(.x(x_50), .z(tmp00_50_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650051(.x(x_51), .z(tmp00_51_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650052(.x(x_52), .z(tmp00_52_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650053(.x(x_53), .z(tmp00_53_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650054(.x(x_54), .z(tmp00_54_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650055(.x(x_55), .z(tmp00_55_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650056(.x(x_56), .z(tmp00_56_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650057(.x(x_57), .z(tmp00_57_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650058(.x(x_58), .z(tmp00_58_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650059(.x(x_59), .z(tmp00_59_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650060(.x(x_60), .z(tmp00_60_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650061(.x(x_61), .z(tmp00_61_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650062(.x(x_62), .z(tmp00_62_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650063(.x(x_63), .z(tmp00_63_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650064(.x(x_64), .z(tmp00_64_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650065(.x(x_65), .z(tmp00_65_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650066(.x(x_66), .z(tmp00_66_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650067(.x(x_67), .z(tmp00_67_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650068(.x(x_68), .z(tmp00_68_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650069(.x(x_69), .z(tmp00_69_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650070(.x(x_70), .z(tmp00_70_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650071(.x(x_71), .z(tmp00_71_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650072(.x(x_72), .z(tmp00_72_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650073(.x(x_73), .z(tmp00_73_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650074(.x(x_74), .z(tmp00_74_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650075(.x(x_75), .z(tmp00_75_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650076(.x(x_76), .z(tmp00_76_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650077(.x(x_77), .z(tmp00_77_65));
	booth_0006 #(.WIDTH(WIDTH)) mul00650078(.x(x_78), .z(tmp00_78_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650079(.x(x_79), .z(tmp00_79_65));
	booth__010 #(.WIDTH(WIDTH)) mul00650080(.x(x_80), .z(tmp00_80_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650081(.x(x_81), .z(tmp00_81_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650082(.x(x_82), .z(tmp00_82_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650083(.x(x_83), .z(tmp00_83_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650084(.x(x_84), .z(tmp00_84_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650085(.x(x_85), .z(tmp00_85_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650086(.x(x_86), .z(tmp00_86_65));
	booth_0010 #(.WIDTH(WIDTH)) mul00650087(.x(x_87), .z(tmp00_87_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650088(.x(x_88), .z(tmp00_88_65));
	booth__006 #(.WIDTH(WIDTH)) mul00650089(.x(x_89), .z(tmp00_89_65));
	booth_0010 #(.WIDTH(WIDTH)) mul00650090(.x(x_90), .z(tmp00_90_65));
	booth_0006 #(.WIDTH(WIDTH)) mul00650091(.x(x_91), .z(tmp00_91_65));
	booth_0006 #(.WIDTH(WIDTH)) mul00650092(.x(x_92), .z(tmp00_92_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650093(.x(x_93), .z(tmp00_93_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650094(.x(x_94), .z(tmp00_94_65));
	booth__006 #(.WIDTH(WIDTH)) mul00650095(.x(x_95), .z(tmp00_95_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650096(.x(x_96), .z(tmp00_96_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650097(.x(x_97), .z(tmp00_97_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650098(.x(x_98), .z(tmp00_98_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650099(.x(x_99), .z(tmp00_99_65));
	booth__010 #(.WIDTH(WIDTH)) mul00650100(.x(x_100), .z(tmp00_100_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650101(.x(x_101), .z(tmp00_101_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650102(.x(x_102), .z(tmp00_102_65));
	booth_0002 #(.WIDTH(WIDTH)) mul00650103(.x(x_103), .z(tmp00_103_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650104(.x(x_104), .z(tmp00_104_65));
	booth_0010 #(.WIDTH(WIDTH)) mul00650105(.x(x_105), .z(tmp00_105_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650106(.x(x_106), .z(tmp00_106_65));
	booth__012 #(.WIDTH(WIDTH)) mul00650107(.x(x_107), .z(tmp00_107_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650108(.x(x_108), .z(tmp00_108_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650109(.x(x_109), .z(tmp00_109_65));
	booth__006 #(.WIDTH(WIDTH)) mul00650110(.x(x_110), .z(tmp00_110_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650111(.x(x_111), .z(tmp00_111_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650112(.x(x_112), .z(tmp00_112_65));
	booth_0006 #(.WIDTH(WIDTH)) mul00650113(.x(x_113), .z(tmp00_113_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650114(.x(x_114), .z(tmp00_114_65));
	booth__006 #(.WIDTH(WIDTH)) mul00650115(.x(x_115), .z(tmp00_115_65));
	booth__008 #(.WIDTH(WIDTH)) mul00650116(.x(x_116), .z(tmp00_116_65));
	booth_0004 #(.WIDTH(WIDTH)) mul00650117(.x(x_117), .z(tmp00_117_65));
	booth__010 #(.WIDTH(WIDTH)) mul00650118(.x(x_118), .z(tmp00_118_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650119(.x(x_119), .z(tmp00_119_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650120(.x(x_120), .z(tmp00_120_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650121(.x(x_121), .z(tmp00_121_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650122(.x(x_122), .z(tmp00_122_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650123(.x(x_123), .z(tmp00_123_65));
	booth__004 #(.WIDTH(WIDTH)) mul00650124(.x(x_124), .z(tmp00_124_65));
	booth__012 #(.WIDTH(WIDTH)) mul00650125(.x(x_125), .z(tmp00_125_65));
	booth_0008 #(.WIDTH(WIDTH)) mul00650126(.x(x_126), .z(tmp00_126_65));
	booth_0000 #(.WIDTH(WIDTH)) mul00650127(.x(x_127), .z(tmp00_127_65));
	booth__010 #(.WIDTH(WIDTH)) mul00660000(.x(x_0), .z(tmp00_0_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660001(.x(x_1), .z(tmp00_1_66));
	booth_0002 #(.WIDTH(WIDTH)) mul00660002(.x(x_2), .z(tmp00_2_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660003(.x(x_3), .z(tmp00_3_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660004(.x(x_4), .z(tmp00_4_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660005(.x(x_5), .z(tmp00_5_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660006(.x(x_6), .z(tmp00_6_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660007(.x(x_7), .z(tmp00_7_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660008(.x(x_8), .z(tmp00_8_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660009(.x(x_9), .z(tmp00_9_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660010(.x(x_10), .z(tmp00_10_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660011(.x(x_11), .z(tmp00_11_66));
	booth_0012 #(.WIDTH(WIDTH)) mul00660012(.x(x_12), .z(tmp00_12_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660013(.x(x_13), .z(tmp00_13_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660014(.x(x_14), .z(tmp00_14_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660015(.x(x_15), .z(tmp00_15_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660016(.x(x_16), .z(tmp00_16_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660017(.x(x_17), .z(tmp00_17_66));
	booth__002 #(.WIDTH(WIDTH)) mul00660018(.x(x_18), .z(tmp00_18_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660019(.x(x_19), .z(tmp00_19_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660020(.x(x_20), .z(tmp00_20_66));
	booth__012 #(.WIDTH(WIDTH)) mul00660021(.x(x_21), .z(tmp00_21_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660022(.x(x_22), .z(tmp00_22_66));
	booth__006 #(.WIDTH(WIDTH)) mul00660023(.x(x_23), .z(tmp00_23_66));
	booth_0006 #(.WIDTH(WIDTH)) mul00660024(.x(x_24), .z(tmp00_24_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660025(.x(x_25), .z(tmp00_25_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660026(.x(x_26), .z(tmp00_26_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660027(.x(x_27), .z(tmp00_27_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660028(.x(x_28), .z(tmp00_28_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660029(.x(x_29), .z(tmp00_29_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660030(.x(x_30), .z(tmp00_30_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660031(.x(x_31), .z(tmp00_31_66));
	booth__006 #(.WIDTH(WIDTH)) mul00660032(.x(x_32), .z(tmp00_32_66));
	booth_0006 #(.WIDTH(WIDTH)) mul00660033(.x(x_33), .z(tmp00_33_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660034(.x(x_34), .z(tmp00_34_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660035(.x(x_35), .z(tmp00_35_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660036(.x(x_36), .z(tmp00_36_66));
	booth_0002 #(.WIDTH(WIDTH)) mul00660037(.x(x_37), .z(tmp00_37_66));
	booth_0006 #(.WIDTH(WIDTH)) mul00660038(.x(x_38), .z(tmp00_38_66));
	booth__012 #(.WIDTH(WIDTH)) mul00660039(.x(x_39), .z(tmp00_39_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660040(.x(x_40), .z(tmp00_40_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660041(.x(x_41), .z(tmp00_41_66));
	booth_0014 #(.WIDTH(WIDTH)) mul00660042(.x(x_42), .z(tmp00_42_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660043(.x(x_43), .z(tmp00_43_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660044(.x(x_44), .z(tmp00_44_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660045(.x(x_45), .z(tmp00_45_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660046(.x(x_46), .z(tmp00_46_66));
	booth_0002 #(.WIDTH(WIDTH)) mul00660047(.x(x_47), .z(tmp00_47_66));
	booth_0002 #(.WIDTH(WIDTH)) mul00660048(.x(x_48), .z(tmp00_48_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660049(.x(x_49), .z(tmp00_49_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660050(.x(x_50), .z(tmp00_50_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660051(.x(x_51), .z(tmp00_51_66));
	booth_0012 #(.WIDTH(WIDTH)) mul00660052(.x(x_52), .z(tmp00_52_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660053(.x(x_53), .z(tmp00_53_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660054(.x(x_54), .z(tmp00_54_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660055(.x(x_55), .z(tmp00_55_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660056(.x(x_56), .z(tmp00_56_66));
	booth__002 #(.WIDTH(WIDTH)) mul00660057(.x(x_57), .z(tmp00_57_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660058(.x(x_58), .z(tmp00_58_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660059(.x(x_59), .z(tmp00_59_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660060(.x(x_60), .z(tmp00_60_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660061(.x(x_61), .z(tmp00_61_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660062(.x(x_62), .z(tmp00_62_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660063(.x(x_63), .z(tmp00_63_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660064(.x(x_64), .z(tmp00_64_66));
	booth_0002 #(.WIDTH(WIDTH)) mul00660065(.x(x_65), .z(tmp00_65_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660066(.x(x_66), .z(tmp00_66_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660067(.x(x_67), .z(tmp00_67_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660068(.x(x_68), .z(tmp00_68_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660069(.x(x_69), .z(tmp00_69_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660070(.x(x_70), .z(tmp00_70_66));
	booth__002 #(.WIDTH(WIDTH)) mul00660071(.x(x_71), .z(tmp00_71_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660072(.x(x_72), .z(tmp00_72_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660073(.x(x_73), .z(tmp00_73_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660074(.x(x_74), .z(tmp00_74_66));
	booth__006 #(.WIDTH(WIDTH)) mul00660075(.x(x_75), .z(tmp00_75_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660076(.x(x_76), .z(tmp00_76_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660077(.x(x_77), .z(tmp00_77_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660078(.x(x_78), .z(tmp00_78_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660079(.x(x_79), .z(tmp00_79_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660080(.x(x_80), .z(tmp00_80_66));
	booth_0010 #(.WIDTH(WIDTH)) mul00660081(.x(x_81), .z(tmp00_81_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660082(.x(x_82), .z(tmp00_82_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660083(.x(x_83), .z(tmp00_83_66));
	booth_0002 #(.WIDTH(WIDTH)) mul00660084(.x(x_84), .z(tmp00_84_66));
	booth_0010 #(.WIDTH(WIDTH)) mul00660085(.x(x_85), .z(tmp00_85_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660086(.x(x_86), .z(tmp00_86_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660087(.x(x_87), .z(tmp00_87_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660088(.x(x_88), .z(tmp00_88_66));
	booth_0006 #(.WIDTH(WIDTH)) mul00660089(.x(x_89), .z(tmp00_89_66));
	booth_0002 #(.WIDTH(WIDTH)) mul00660090(.x(x_90), .z(tmp00_90_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660091(.x(x_91), .z(tmp00_91_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660092(.x(x_92), .z(tmp00_92_66));
	booth__012 #(.WIDTH(WIDTH)) mul00660093(.x(x_93), .z(tmp00_93_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660094(.x(x_94), .z(tmp00_94_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660095(.x(x_95), .z(tmp00_95_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660096(.x(x_96), .z(tmp00_96_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660097(.x(x_97), .z(tmp00_97_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660098(.x(x_98), .z(tmp00_98_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660099(.x(x_99), .z(tmp00_99_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660100(.x(x_100), .z(tmp00_100_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660101(.x(x_101), .z(tmp00_101_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660102(.x(x_102), .z(tmp00_102_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660103(.x(x_103), .z(tmp00_103_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660104(.x(x_104), .z(tmp00_104_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660105(.x(x_105), .z(tmp00_105_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660106(.x(x_106), .z(tmp00_106_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660107(.x(x_107), .z(tmp00_107_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660108(.x(x_108), .z(tmp00_108_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660109(.x(x_109), .z(tmp00_109_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660110(.x(x_110), .z(tmp00_110_66));
	booth__006 #(.WIDTH(WIDTH)) mul00660111(.x(x_111), .z(tmp00_111_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660112(.x(x_112), .z(tmp00_112_66));
	booth__006 #(.WIDTH(WIDTH)) mul00660113(.x(x_113), .z(tmp00_113_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660114(.x(x_114), .z(tmp00_114_66));
	booth_0006 #(.WIDTH(WIDTH)) mul00660115(.x(x_115), .z(tmp00_115_66));
	booth_0000 #(.WIDTH(WIDTH)) mul00660116(.x(x_116), .z(tmp00_116_66));
	booth_0006 #(.WIDTH(WIDTH)) mul00660117(.x(x_117), .z(tmp00_117_66));
	booth_0010 #(.WIDTH(WIDTH)) mul00660118(.x(x_118), .z(tmp00_118_66));
	booth_0012 #(.WIDTH(WIDTH)) mul00660119(.x(x_119), .z(tmp00_119_66));
	booth__002 #(.WIDTH(WIDTH)) mul00660120(.x(x_120), .z(tmp00_120_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660121(.x(x_121), .z(tmp00_121_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660122(.x(x_122), .z(tmp00_122_66));
	booth__004 #(.WIDTH(WIDTH)) mul00660123(.x(x_123), .z(tmp00_123_66));
	booth__008 #(.WIDTH(WIDTH)) mul00660124(.x(x_124), .z(tmp00_124_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660125(.x(x_125), .z(tmp00_125_66));
	booth_0008 #(.WIDTH(WIDTH)) mul00660126(.x(x_126), .z(tmp00_126_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00660127(.x(x_127), .z(tmp00_127_66));
	booth_0004 #(.WIDTH(WIDTH)) mul00670000(.x(x_0), .z(tmp00_0_67));
	booth_0006 #(.WIDTH(WIDTH)) mul00670001(.x(x_1), .z(tmp00_1_67));
	booth__002 #(.WIDTH(WIDTH)) mul00670002(.x(x_2), .z(tmp00_2_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670003(.x(x_3), .z(tmp00_3_67));
	booth__016 #(.WIDTH(WIDTH)) mul00670004(.x(x_4), .z(tmp00_4_67));
	booth_0002 #(.WIDTH(WIDTH)) mul00670005(.x(x_5), .z(tmp00_5_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670006(.x(x_6), .z(tmp00_6_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670007(.x(x_7), .z(tmp00_7_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670008(.x(x_8), .z(tmp00_8_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670009(.x(x_9), .z(tmp00_9_67));
	booth__012 #(.WIDTH(WIDTH)) mul00670010(.x(x_10), .z(tmp00_10_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670011(.x(x_11), .z(tmp00_11_67));
	booth_0002 #(.WIDTH(WIDTH)) mul00670012(.x(x_12), .z(tmp00_12_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670013(.x(x_13), .z(tmp00_13_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670014(.x(x_14), .z(tmp00_14_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670015(.x(x_15), .z(tmp00_15_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670016(.x(x_16), .z(tmp00_16_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670017(.x(x_17), .z(tmp00_17_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670018(.x(x_18), .z(tmp00_18_67));
	booth_0010 #(.WIDTH(WIDTH)) mul00670019(.x(x_19), .z(tmp00_19_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670020(.x(x_20), .z(tmp00_20_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670021(.x(x_21), .z(tmp00_21_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670022(.x(x_22), .z(tmp00_22_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670023(.x(x_23), .z(tmp00_23_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670024(.x(x_24), .z(tmp00_24_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670025(.x(x_25), .z(tmp00_25_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670026(.x(x_26), .z(tmp00_26_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670027(.x(x_27), .z(tmp00_27_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670028(.x(x_28), .z(tmp00_28_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670029(.x(x_29), .z(tmp00_29_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670030(.x(x_30), .z(tmp00_30_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670031(.x(x_31), .z(tmp00_31_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670032(.x(x_32), .z(tmp00_32_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670033(.x(x_33), .z(tmp00_33_67));
	booth__002 #(.WIDTH(WIDTH)) mul00670034(.x(x_34), .z(tmp00_34_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670035(.x(x_35), .z(tmp00_35_67));
	booth_0006 #(.WIDTH(WIDTH)) mul00670036(.x(x_36), .z(tmp00_36_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670037(.x(x_37), .z(tmp00_37_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670038(.x(x_38), .z(tmp00_38_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670039(.x(x_39), .z(tmp00_39_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670040(.x(x_40), .z(tmp00_40_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670041(.x(x_41), .z(tmp00_41_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670042(.x(x_42), .z(tmp00_42_67));
	booth__002 #(.WIDTH(WIDTH)) mul00670043(.x(x_43), .z(tmp00_43_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670044(.x(x_44), .z(tmp00_44_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670045(.x(x_45), .z(tmp00_45_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670046(.x(x_46), .z(tmp00_46_67));
	booth_0012 #(.WIDTH(WIDTH)) mul00670047(.x(x_47), .z(tmp00_47_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670048(.x(x_48), .z(tmp00_48_67));
	booth_0016 #(.WIDTH(WIDTH)) mul00670049(.x(x_49), .z(tmp00_49_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670050(.x(x_50), .z(tmp00_50_67));
	booth__012 #(.WIDTH(WIDTH)) mul00670051(.x(x_51), .z(tmp00_51_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670052(.x(x_52), .z(tmp00_52_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670053(.x(x_53), .z(tmp00_53_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670054(.x(x_54), .z(tmp00_54_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670055(.x(x_55), .z(tmp00_55_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670056(.x(x_56), .z(tmp00_56_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670057(.x(x_57), .z(tmp00_57_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670058(.x(x_58), .z(tmp00_58_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670059(.x(x_59), .z(tmp00_59_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670060(.x(x_60), .z(tmp00_60_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670061(.x(x_61), .z(tmp00_61_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670062(.x(x_62), .z(tmp00_62_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670063(.x(x_63), .z(tmp00_63_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670064(.x(x_64), .z(tmp00_64_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670065(.x(x_65), .z(tmp00_65_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670066(.x(x_66), .z(tmp00_66_67));
	booth_0010 #(.WIDTH(WIDTH)) mul00670067(.x(x_67), .z(tmp00_67_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670068(.x(x_68), .z(tmp00_68_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670069(.x(x_69), .z(tmp00_69_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670070(.x(x_70), .z(tmp00_70_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670071(.x(x_71), .z(tmp00_71_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670072(.x(x_72), .z(tmp00_72_67));
	booth__006 #(.WIDTH(WIDTH)) mul00670073(.x(x_73), .z(tmp00_73_67));
	booth_0006 #(.WIDTH(WIDTH)) mul00670074(.x(x_74), .z(tmp00_74_67));
	booth_0012 #(.WIDTH(WIDTH)) mul00670075(.x(x_75), .z(tmp00_75_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670076(.x(x_76), .z(tmp00_76_67));
	booth_0006 #(.WIDTH(WIDTH)) mul00670077(.x(x_77), .z(tmp00_77_67));
	booth_0012 #(.WIDTH(WIDTH)) mul00670078(.x(x_78), .z(tmp00_78_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670079(.x(x_79), .z(tmp00_79_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670080(.x(x_80), .z(tmp00_80_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670081(.x(x_81), .z(tmp00_81_67));
	booth__006 #(.WIDTH(WIDTH)) mul00670082(.x(x_82), .z(tmp00_82_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670083(.x(x_83), .z(tmp00_83_67));
	booth__002 #(.WIDTH(WIDTH)) mul00670084(.x(x_84), .z(tmp00_84_67));
	booth__016 #(.WIDTH(WIDTH)) mul00670085(.x(x_85), .z(tmp00_85_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670086(.x(x_86), .z(tmp00_86_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670087(.x(x_87), .z(tmp00_87_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670088(.x(x_88), .z(tmp00_88_67));
	booth__010 #(.WIDTH(WIDTH)) mul00670089(.x(x_89), .z(tmp00_89_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670090(.x(x_90), .z(tmp00_90_67));
	booth__012 #(.WIDTH(WIDTH)) mul00670091(.x(x_91), .z(tmp00_91_67));
	booth_0012 #(.WIDTH(WIDTH)) mul00670092(.x(x_92), .z(tmp00_92_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670093(.x(x_93), .z(tmp00_93_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670094(.x(x_94), .z(tmp00_94_67));
	booth__002 #(.WIDTH(WIDTH)) mul00670095(.x(x_95), .z(tmp00_95_67));
	booth_0006 #(.WIDTH(WIDTH)) mul00670096(.x(x_96), .z(tmp00_96_67));
	booth__008 #(.WIDTH(WIDTH)) mul00670097(.x(x_97), .z(tmp00_97_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670098(.x(x_98), .z(tmp00_98_67));
	booth_0012 #(.WIDTH(WIDTH)) mul00670099(.x(x_99), .z(tmp00_99_67));
	booth_0016 #(.WIDTH(WIDTH)) mul00670100(.x(x_100), .z(tmp00_100_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670101(.x(x_101), .z(tmp00_101_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670102(.x(x_102), .z(tmp00_102_67));
	booth__006 #(.WIDTH(WIDTH)) mul00670103(.x(x_103), .z(tmp00_103_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670104(.x(x_104), .z(tmp00_104_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670105(.x(x_105), .z(tmp00_105_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670106(.x(x_106), .z(tmp00_106_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670107(.x(x_107), .z(tmp00_107_67));
	booth__012 #(.WIDTH(WIDTH)) mul00670108(.x(x_108), .z(tmp00_108_67));
	booth_0016 #(.WIDTH(WIDTH)) mul00670109(.x(x_109), .z(tmp00_109_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670110(.x(x_110), .z(tmp00_110_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670111(.x(x_111), .z(tmp00_111_67));
	booth__002 #(.WIDTH(WIDTH)) mul00670112(.x(x_112), .z(tmp00_112_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670113(.x(x_113), .z(tmp00_113_67));
	booth_0002 #(.WIDTH(WIDTH)) mul00670114(.x(x_114), .z(tmp00_114_67));
	booth__016 #(.WIDTH(WIDTH)) mul00670115(.x(x_115), .z(tmp00_115_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670116(.x(x_116), .z(tmp00_116_67));
	booth_0008 #(.WIDTH(WIDTH)) mul00670117(.x(x_117), .z(tmp00_117_67));
	booth_0004 #(.WIDTH(WIDTH)) mul00670118(.x(x_118), .z(tmp00_118_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670119(.x(x_119), .z(tmp00_119_67));
	booth__016 #(.WIDTH(WIDTH)) mul00670120(.x(x_120), .z(tmp00_120_67));
	booth__004 #(.WIDTH(WIDTH)) mul00670121(.x(x_121), .z(tmp00_121_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670122(.x(x_122), .z(tmp00_122_67));
	booth__006 #(.WIDTH(WIDTH)) mul00670123(.x(x_123), .z(tmp00_123_67));
	booth_0016 #(.WIDTH(WIDTH)) mul00670124(.x(x_124), .z(tmp00_124_67));
	booth__002 #(.WIDTH(WIDTH)) mul00670125(.x(x_125), .z(tmp00_125_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670126(.x(x_126), .z(tmp00_126_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00670127(.x(x_127), .z(tmp00_127_67));
	booth_0000 #(.WIDTH(WIDTH)) mul00680000(.x(x_0), .z(tmp00_0_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680001(.x(x_1), .z(tmp00_1_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680002(.x(x_2), .z(tmp00_2_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680003(.x(x_3), .z(tmp00_3_68));
	booth__016 #(.WIDTH(WIDTH)) mul00680004(.x(x_4), .z(tmp00_4_68));
	booth__010 #(.WIDTH(WIDTH)) mul00680005(.x(x_5), .z(tmp00_5_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680006(.x(x_6), .z(tmp00_6_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680007(.x(x_7), .z(tmp00_7_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680008(.x(x_8), .z(tmp00_8_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680009(.x(x_9), .z(tmp00_9_68));
	booth_0006 #(.WIDTH(WIDTH)) mul00680010(.x(x_10), .z(tmp00_10_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680011(.x(x_11), .z(tmp00_11_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680012(.x(x_12), .z(tmp00_12_68));
	booth_0012 #(.WIDTH(WIDTH)) mul00680013(.x(x_13), .z(tmp00_13_68));
	booth_0006 #(.WIDTH(WIDTH)) mul00680014(.x(x_14), .z(tmp00_14_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680015(.x(x_15), .z(tmp00_15_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680016(.x(x_16), .z(tmp00_16_68));
	booth_0002 #(.WIDTH(WIDTH)) mul00680017(.x(x_17), .z(tmp00_17_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680018(.x(x_18), .z(tmp00_18_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680019(.x(x_19), .z(tmp00_19_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680020(.x(x_20), .z(tmp00_20_68));
	booth_0002 #(.WIDTH(WIDTH)) mul00680021(.x(x_21), .z(tmp00_21_68));
	booth_0016 #(.WIDTH(WIDTH)) mul00680022(.x(x_22), .z(tmp00_22_68));
	booth__010 #(.WIDTH(WIDTH)) mul00680023(.x(x_23), .z(tmp00_23_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680024(.x(x_24), .z(tmp00_24_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680025(.x(x_25), .z(tmp00_25_68));
	booth_0012 #(.WIDTH(WIDTH)) mul00680026(.x(x_26), .z(tmp00_26_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680027(.x(x_27), .z(tmp00_27_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680028(.x(x_28), .z(tmp00_28_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680029(.x(x_29), .z(tmp00_29_68));
	booth_0010 #(.WIDTH(WIDTH)) mul00680030(.x(x_30), .z(tmp00_30_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680031(.x(x_31), .z(tmp00_31_68));
	booth__006 #(.WIDTH(WIDTH)) mul00680032(.x(x_32), .z(tmp00_32_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680033(.x(x_33), .z(tmp00_33_68));
	booth_0012 #(.WIDTH(WIDTH)) mul00680034(.x(x_34), .z(tmp00_34_68));
	booth_0002 #(.WIDTH(WIDTH)) mul00680035(.x(x_35), .z(tmp00_35_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680036(.x(x_36), .z(tmp00_36_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680037(.x(x_37), .z(tmp00_37_68));
	booth__016 #(.WIDTH(WIDTH)) mul00680038(.x(x_38), .z(tmp00_38_68));
	booth_0020 #(.WIDTH(WIDTH)) mul00680039(.x(x_39), .z(tmp00_39_68));
	booth_0012 #(.WIDTH(WIDTH)) mul00680040(.x(x_40), .z(tmp00_40_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680041(.x(x_41), .z(tmp00_41_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680042(.x(x_42), .z(tmp00_42_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680043(.x(x_43), .z(tmp00_43_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680044(.x(x_44), .z(tmp00_44_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680045(.x(x_45), .z(tmp00_45_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680046(.x(x_46), .z(tmp00_46_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680047(.x(x_47), .z(tmp00_47_68));
	booth_0006 #(.WIDTH(WIDTH)) mul00680048(.x(x_48), .z(tmp00_48_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680049(.x(x_49), .z(tmp00_49_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680050(.x(x_50), .z(tmp00_50_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680051(.x(x_51), .z(tmp00_51_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680052(.x(x_52), .z(tmp00_52_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680053(.x(x_53), .z(tmp00_53_68));
	booth_0012 #(.WIDTH(WIDTH)) mul00680054(.x(x_54), .z(tmp00_54_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680055(.x(x_55), .z(tmp00_55_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680056(.x(x_56), .z(tmp00_56_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680057(.x(x_57), .z(tmp00_57_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680058(.x(x_58), .z(tmp00_58_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680059(.x(x_59), .z(tmp00_59_68));
	booth__010 #(.WIDTH(WIDTH)) mul00680060(.x(x_60), .z(tmp00_60_68));
	booth_0006 #(.WIDTH(WIDTH)) mul00680061(.x(x_61), .z(tmp00_61_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680062(.x(x_62), .z(tmp00_62_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680063(.x(x_63), .z(tmp00_63_68));
	booth__006 #(.WIDTH(WIDTH)) mul00680064(.x(x_64), .z(tmp00_64_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680065(.x(x_65), .z(tmp00_65_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680066(.x(x_66), .z(tmp00_66_68));
	booth_0006 #(.WIDTH(WIDTH)) mul00680067(.x(x_67), .z(tmp00_67_68));
	booth_0016 #(.WIDTH(WIDTH)) mul00680068(.x(x_68), .z(tmp00_68_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680069(.x(x_69), .z(tmp00_69_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680070(.x(x_70), .z(tmp00_70_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680071(.x(x_71), .z(tmp00_71_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680072(.x(x_72), .z(tmp00_72_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680073(.x(x_73), .z(tmp00_73_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680074(.x(x_74), .z(tmp00_74_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680075(.x(x_75), .z(tmp00_75_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680076(.x(x_76), .z(tmp00_76_68));
	booth_0010 #(.WIDTH(WIDTH)) mul00680077(.x(x_77), .z(tmp00_77_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680078(.x(x_78), .z(tmp00_78_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680079(.x(x_79), .z(tmp00_79_68));
	booth_0012 #(.WIDTH(WIDTH)) mul00680080(.x(x_80), .z(tmp00_80_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680081(.x(x_81), .z(tmp00_81_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680082(.x(x_82), .z(tmp00_82_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680083(.x(x_83), .z(tmp00_83_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680084(.x(x_84), .z(tmp00_84_68));
	booth_0014 #(.WIDTH(WIDTH)) mul00680085(.x(x_85), .z(tmp00_85_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680086(.x(x_86), .z(tmp00_86_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680087(.x(x_87), .z(tmp00_87_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680088(.x(x_88), .z(tmp00_88_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680089(.x(x_89), .z(tmp00_89_68));
	booth_0012 #(.WIDTH(WIDTH)) mul00680090(.x(x_90), .z(tmp00_90_68));
	booth_0010 #(.WIDTH(WIDTH)) mul00680091(.x(x_91), .z(tmp00_91_68));
	booth_0016 #(.WIDTH(WIDTH)) mul00680092(.x(x_92), .z(tmp00_92_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680093(.x(x_93), .z(tmp00_93_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680094(.x(x_94), .z(tmp00_94_68));
	booth__012 #(.WIDTH(WIDTH)) mul00680095(.x(x_95), .z(tmp00_95_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680096(.x(x_96), .z(tmp00_96_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680097(.x(x_97), .z(tmp00_97_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680098(.x(x_98), .z(tmp00_98_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680099(.x(x_99), .z(tmp00_99_68));
	booth_0012 #(.WIDTH(WIDTH)) mul00680100(.x(x_100), .z(tmp00_100_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680101(.x(x_101), .z(tmp00_101_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680102(.x(x_102), .z(tmp00_102_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680103(.x(x_103), .z(tmp00_103_68));
	booth__006 #(.WIDTH(WIDTH)) mul00680104(.x(x_104), .z(tmp00_104_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680105(.x(x_105), .z(tmp00_105_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680106(.x(x_106), .z(tmp00_106_68));
	booth__012 #(.WIDTH(WIDTH)) mul00680107(.x(x_107), .z(tmp00_107_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680108(.x(x_108), .z(tmp00_108_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680109(.x(x_109), .z(tmp00_109_68));
	booth__004 #(.WIDTH(WIDTH)) mul00680110(.x(x_110), .z(tmp00_110_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680111(.x(x_111), .z(tmp00_111_68));
	booth_0010 #(.WIDTH(WIDTH)) mul00680112(.x(x_112), .z(tmp00_112_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680113(.x(x_113), .z(tmp00_113_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680114(.x(x_114), .z(tmp00_114_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680115(.x(x_115), .z(tmp00_115_68));
	booth__002 #(.WIDTH(WIDTH)) mul00680116(.x(x_116), .z(tmp00_116_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680117(.x(x_117), .z(tmp00_117_68));
	booth__010 #(.WIDTH(WIDTH)) mul00680118(.x(x_118), .z(tmp00_118_68));
	booth__012 #(.WIDTH(WIDTH)) mul00680119(.x(x_119), .z(tmp00_119_68));
	booth_0016 #(.WIDTH(WIDTH)) mul00680120(.x(x_120), .z(tmp00_120_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680121(.x(x_121), .z(tmp00_121_68));
	booth__008 #(.WIDTH(WIDTH)) mul00680122(.x(x_122), .z(tmp00_122_68));
	booth_0008 #(.WIDTH(WIDTH)) mul00680123(.x(x_123), .z(tmp00_123_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680124(.x(x_124), .z(tmp00_124_68));
	booth_0004 #(.WIDTH(WIDTH)) mul00680125(.x(x_125), .z(tmp00_125_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680126(.x(x_126), .z(tmp00_126_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00680127(.x(x_127), .z(tmp00_127_68));
	booth_0000 #(.WIDTH(WIDTH)) mul00690000(.x(x_0), .z(tmp00_0_69));
	booth_0010 #(.WIDTH(WIDTH)) mul00690001(.x(x_1), .z(tmp00_1_69));
	booth_0002 #(.WIDTH(WIDTH)) mul00690002(.x(x_2), .z(tmp00_2_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690003(.x(x_3), .z(tmp00_3_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690004(.x(x_4), .z(tmp00_4_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690005(.x(x_5), .z(tmp00_5_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690006(.x(x_6), .z(tmp00_6_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690007(.x(x_7), .z(tmp00_7_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690008(.x(x_8), .z(tmp00_8_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690009(.x(x_9), .z(tmp00_9_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690010(.x(x_10), .z(tmp00_10_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690011(.x(x_11), .z(tmp00_11_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690012(.x(x_12), .z(tmp00_12_69));
	booth__002 #(.WIDTH(WIDTH)) mul00690013(.x(x_13), .z(tmp00_13_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690014(.x(x_14), .z(tmp00_14_69));
	booth__002 #(.WIDTH(WIDTH)) mul00690015(.x(x_15), .z(tmp00_15_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690016(.x(x_16), .z(tmp00_16_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690017(.x(x_17), .z(tmp00_17_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690018(.x(x_18), .z(tmp00_18_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690019(.x(x_19), .z(tmp00_19_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690020(.x(x_20), .z(tmp00_20_69));
	booth_0002 #(.WIDTH(WIDTH)) mul00690021(.x(x_21), .z(tmp00_21_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690022(.x(x_22), .z(tmp00_22_69));
	booth__002 #(.WIDTH(WIDTH)) mul00690023(.x(x_23), .z(tmp00_23_69));
	booth_0002 #(.WIDTH(WIDTH)) mul00690024(.x(x_24), .z(tmp00_24_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690025(.x(x_25), .z(tmp00_25_69));
	booth_0010 #(.WIDTH(WIDTH)) mul00690026(.x(x_26), .z(tmp00_26_69));
	booth_0002 #(.WIDTH(WIDTH)) mul00690027(.x(x_27), .z(tmp00_27_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690028(.x(x_28), .z(tmp00_28_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690029(.x(x_29), .z(tmp00_29_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690030(.x(x_30), .z(tmp00_30_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690031(.x(x_31), .z(tmp00_31_69));
	booth__006 #(.WIDTH(WIDTH)) mul00690032(.x(x_32), .z(tmp00_32_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690033(.x(x_33), .z(tmp00_33_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690034(.x(x_34), .z(tmp00_34_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690035(.x(x_35), .z(tmp00_35_69));
	booth_0006 #(.WIDTH(WIDTH)) mul00690036(.x(x_36), .z(tmp00_36_69));
	booth_0006 #(.WIDTH(WIDTH)) mul00690037(.x(x_37), .z(tmp00_37_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690038(.x(x_38), .z(tmp00_38_69));
	booth_0010 #(.WIDTH(WIDTH)) mul00690039(.x(x_39), .z(tmp00_39_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690040(.x(x_40), .z(tmp00_40_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690041(.x(x_41), .z(tmp00_41_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690042(.x(x_42), .z(tmp00_42_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690043(.x(x_43), .z(tmp00_43_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690044(.x(x_44), .z(tmp00_44_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690045(.x(x_45), .z(tmp00_45_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690046(.x(x_46), .z(tmp00_46_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690047(.x(x_47), .z(tmp00_47_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690048(.x(x_48), .z(tmp00_48_69));
	booth__002 #(.WIDTH(WIDTH)) mul00690049(.x(x_49), .z(tmp00_49_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690050(.x(x_50), .z(tmp00_50_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690051(.x(x_51), .z(tmp00_51_69));
	booth_0006 #(.WIDTH(WIDTH)) mul00690052(.x(x_52), .z(tmp00_52_69));
	booth__002 #(.WIDTH(WIDTH)) mul00690053(.x(x_53), .z(tmp00_53_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690054(.x(x_54), .z(tmp00_54_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690055(.x(x_55), .z(tmp00_55_69));
	booth_0010 #(.WIDTH(WIDTH)) mul00690056(.x(x_56), .z(tmp00_56_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690057(.x(x_57), .z(tmp00_57_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690058(.x(x_58), .z(tmp00_58_69));
	booth__006 #(.WIDTH(WIDTH)) mul00690059(.x(x_59), .z(tmp00_59_69));
	booth__006 #(.WIDTH(WIDTH)) mul00690060(.x(x_60), .z(tmp00_60_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690061(.x(x_61), .z(tmp00_61_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690062(.x(x_62), .z(tmp00_62_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690063(.x(x_63), .z(tmp00_63_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690064(.x(x_64), .z(tmp00_64_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690065(.x(x_65), .z(tmp00_65_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690066(.x(x_66), .z(tmp00_66_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690067(.x(x_67), .z(tmp00_67_69));
	booth_0006 #(.WIDTH(WIDTH)) mul00690068(.x(x_68), .z(tmp00_68_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690069(.x(x_69), .z(tmp00_69_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690070(.x(x_70), .z(tmp00_70_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690071(.x(x_71), .z(tmp00_71_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690072(.x(x_72), .z(tmp00_72_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690073(.x(x_73), .z(tmp00_73_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690074(.x(x_74), .z(tmp00_74_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690075(.x(x_75), .z(tmp00_75_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690076(.x(x_76), .z(tmp00_76_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690077(.x(x_77), .z(tmp00_77_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690078(.x(x_78), .z(tmp00_78_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690079(.x(x_79), .z(tmp00_79_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690080(.x(x_80), .z(tmp00_80_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690081(.x(x_81), .z(tmp00_81_69));
	booth__012 #(.WIDTH(WIDTH)) mul00690082(.x(x_82), .z(tmp00_82_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690083(.x(x_83), .z(tmp00_83_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690084(.x(x_84), .z(tmp00_84_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690085(.x(x_85), .z(tmp00_85_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690086(.x(x_86), .z(tmp00_86_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690087(.x(x_87), .z(tmp00_87_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690088(.x(x_88), .z(tmp00_88_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690089(.x(x_89), .z(tmp00_89_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690090(.x(x_90), .z(tmp00_90_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690091(.x(x_91), .z(tmp00_91_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690092(.x(x_92), .z(tmp00_92_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690093(.x(x_93), .z(tmp00_93_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690094(.x(x_94), .z(tmp00_94_69));
	booth_0010 #(.WIDTH(WIDTH)) mul00690095(.x(x_95), .z(tmp00_95_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690096(.x(x_96), .z(tmp00_96_69));
	booth__006 #(.WIDTH(WIDTH)) mul00690097(.x(x_97), .z(tmp00_97_69));
	booth__006 #(.WIDTH(WIDTH)) mul00690098(.x(x_98), .z(tmp00_98_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690099(.x(x_99), .z(tmp00_99_69));
	booth_0002 #(.WIDTH(WIDTH)) mul00690100(.x(x_100), .z(tmp00_100_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690101(.x(x_101), .z(tmp00_101_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690102(.x(x_102), .z(tmp00_102_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690103(.x(x_103), .z(tmp00_103_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690104(.x(x_104), .z(tmp00_104_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690105(.x(x_105), .z(tmp00_105_69));
	booth__006 #(.WIDTH(WIDTH)) mul00690106(.x(x_106), .z(tmp00_106_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690107(.x(x_107), .z(tmp00_107_69));
	booth_0002 #(.WIDTH(WIDTH)) mul00690108(.x(x_108), .z(tmp00_108_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690109(.x(x_109), .z(tmp00_109_69));
	booth_0012 #(.WIDTH(WIDTH)) mul00690110(.x(x_110), .z(tmp00_110_69));
	booth__002 #(.WIDTH(WIDTH)) mul00690111(.x(x_111), .z(tmp00_111_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690112(.x(x_112), .z(tmp00_112_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690113(.x(x_113), .z(tmp00_113_69));
	booth__002 #(.WIDTH(WIDTH)) mul00690114(.x(x_114), .z(tmp00_114_69));
	booth_0006 #(.WIDTH(WIDTH)) mul00690115(.x(x_115), .z(tmp00_115_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690116(.x(x_116), .z(tmp00_116_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690117(.x(x_117), .z(tmp00_117_69));
	booth__012 #(.WIDTH(WIDTH)) mul00690118(.x(x_118), .z(tmp00_118_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690119(.x(x_119), .z(tmp00_119_69));
	booth__008 #(.WIDTH(WIDTH)) mul00690120(.x(x_120), .z(tmp00_120_69));
	booth__004 #(.WIDTH(WIDTH)) mul00690121(.x(x_121), .z(tmp00_121_69));
	booth_0010 #(.WIDTH(WIDTH)) mul00690122(.x(x_122), .z(tmp00_122_69));
	booth_0008 #(.WIDTH(WIDTH)) mul00690123(.x(x_123), .z(tmp00_123_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690124(.x(x_124), .z(tmp00_124_69));
	booth_0000 #(.WIDTH(WIDTH)) mul00690125(.x(x_125), .z(tmp00_125_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00690126(.x(x_126), .z(tmp00_126_69));
	booth__010 #(.WIDTH(WIDTH)) mul00690127(.x(x_127), .z(tmp00_127_69));
	booth_0004 #(.WIDTH(WIDTH)) mul00700000(.x(x_0), .z(tmp00_0_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700001(.x(x_1), .z(tmp00_1_70));
	booth_0012 #(.WIDTH(WIDTH)) mul00700002(.x(x_2), .z(tmp00_2_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700003(.x(x_3), .z(tmp00_3_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700004(.x(x_4), .z(tmp00_4_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700005(.x(x_5), .z(tmp00_5_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700006(.x(x_6), .z(tmp00_6_70));
	booth_0010 #(.WIDTH(WIDTH)) mul00700007(.x(x_7), .z(tmp00_7_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700008(.x(x_8), .z(tmp00_8_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700009(.x(x_9), .z(tmp00_9_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700010(.x(x_10), .z(tmp00_10_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700011(.x(x_11), .z(tmp00_11_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700012(.x(x_12), .z(tmp00_12_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700013(.x(x_13), .z(tmp00_13_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700014(.x(x_14), .z(tmp00_14_70));
	booth_0012 #(.WIDTH(WIDTH)) mul00700015(.x(x_15), .z(tmp00_15_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700016(.x(x_16), .z(tmp00_16_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700017(.x(x_17), .z(tmp00_17_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700018(.x(x_18), .z(tmp00_18_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700019(.x(x_19), .z(tmp00_19_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700020(.x(x_20), .z(tmp00_20_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700021(.x(x_21), .z(tmp00_21_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700022(.x(x_22), .z(tmp00_22_70));
	booth__006 #(.WIDTH(WIDTH)) mul00700023(.x(x_23), .z(tmp00_23_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700024(.x(x_24), .z(tmp00_24_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700025(.x(x_25), .z(tmp00_25_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700026(.x(x_26), .z(tmp00_26_70));
	booth_0012 #(.WIDTH(WIDTH)) mul00700027(.x(x_27), .z(tmp00_27_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700028(.x(x_28), .z(tmp00_28_70));
	booth__002 #(.WIDTH(WIDTH)) mul00700029(.x(x_29), .z(tmp00_29_70));
	booth__006 #(.WIDTH(WIDTH)) mul00700030(.x(x_30), .z(tmp00_30_70));
	booth_0002 #(.WIDTH(WIDTH)) mul00700031(.x(x_31), .z(tmp00_31_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700032(.x(x_32), .z(tmp00_32_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700033(.x(x_33), .z(tmp00_33_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700034(.x(x_34), .z(tmp00_34_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700035(.x(x_35), .z(tmp00_35_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700036(.x(x_36), .z(tmp00_36_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700037(.x(x_37), .z(tmp00_37_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700038(.x(x_38), .z(tmp00_38_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700039(.x(x_39), .z(tmp00_39_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700040(.x(x_40), .z(tmp00_40_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700041(.x(x_41), .z(tmp00_41_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700042(.x(x_42), .z(tmp00_42_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700043(.x(x_43), .z(tmp00_43_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700044(.x(x_44), .z(tmp00_44_70));
	booth_0006 #(.WIDTH(WIDTH)) mul00700045(.x(x_45), .z(tmp00_45_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700046(.x(x_46), .z(tmp00_46_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700047(.x(x_47), .z(tmp00_47_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700048(.x(x_48), .z(tmp00_48_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700049(.x(x_49), .z(tmp00_49_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700050(.x(x_50), .z(tmp00_50_70));
	booth_0006 #(.WIDTH(WIDTH)) mul00700051(.x(x_51), .z(tmp00_51_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700052(.x(x_52), .z(tmp00_52_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700053(.x(x_53), .z(tmp00_53_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700054(.x(x_54), .z(tmp00_54_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700055(.x(x_55), .z(tmp00_55_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700056(.x(x_56), .z(tmp00_56_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700057(.x(x_57), .z(tmp00_57_70));
	booth__012 #(.WIDTH(WIDTH)) mul00700058(.x(x_58), .z(tmp00_58_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700059(.x(x_59), .z(tmp00_59_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700060(.x(x_60), .z(tmp00_60_70));
	booth__002 #(.WIDTH(WIDTH)) mul00700061(.x(x_61), .z(tmp00_61_70));
	booth__006 #(.WIDTH(WIDTH)) mul00700062(.x(x_62), .z(tmp00_62_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700063(.x(x_63), .z(tmp00_63_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700064(.x(x_64), .z(tmp00_64_70));
	booth_0010 #(.WIDTH(WIDTH)) mul00700065(.x(x_65), .z(tmp00_65_70));
	booth__002 #(.WIDTH(WIDTH)) mul00700066(.x(x_66), .z(tmp00_66_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700067(.x(x_67), .z(tmp00_67_70));
	booth_0006 #(.WIDTH(WIDTH)) mul00700068(.x(x_68), .z(tmp00_68_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700069(.x(x_69), .z(tmp00_69_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700070(.x(x_70), .z(tmp00_70_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700071(.x(x_71), .z(tmp00_71_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700072(.x(x_72), .z(tmp00_72_70));
	booth_0010 #(.WIDTH(WIDTH)) mul00700073(.x(x_73), .z(tmp00_73_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700074(.x(x_74), .z(tmp00_74_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700075(.x(x_75), .z(tmp00_75_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700076(.x(x_76), .z(tmp00_76_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700077(.x(x_77), .z(tmp00_77_70));
	booth_0010 #(.WIDTH(WIDTH)) mul00700078(.x(x_78), .z(tmp00_78_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700079(.x(x_79), .z(tmp00_79_70));
	booth__010 #(.WIDTH(WIDTH)) mul00700080(.x(x_80), .z(tmp00_80_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700081(.x(x_81), .z(tmp00_81_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700082(.x(x_82), .z(tmp00_82_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700083(.x(x_83), .z(tmp00_83_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700084(.x(x_84), .z(tmp00_84_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700085(.x(x_85), .z(tmp00_85_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700086(.x(x_86), .z(tmp00_86_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700087(.x(x_87), .z(tmp00_87_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700088(.x(x_88), .z(tmp00_88_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700089(.x(x_89), .z(tmp00_89_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700090(.x(x_90), .z(tmp00_90_70));
	booth_0010 #(.WIDTH(WIDTH)) mul00700091(.x(x_91), .z(tmp00_91_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700092(.x(x_92), .z(tmp00_92_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700093(.x(x_93), .z(tmp00_93_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700094(.x(x_94), .z(tmp00_94_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700095(.x(x_95), .z(tmp00_95_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700096(.x(x_96), .z(tmp00_96_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700097(.x(x_97), .z(tmp00_97_70));
	booth_0004 #(.WIDTH(WIDTH)) mul00700098(.x(x_98), .z(tmp00_98_70));
	booth__002 #(.WIDTH(WIDTH)) mul00700099(.x(x_99), .z(tmp00_99_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700100(.x(x_100), .z(tmp00_100_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700101(.x(x_101), .z(tmp00_101_70));
	booth_0006 #(.WIDTH(WIDTH)) mul00700102(.x(x_102), .z(tmp00_102_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700103(.x(x_103), .z(tmp00_103_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700104(.x(x_104), .z(tmp00_104_70));
	booth__002 #(.WIDTH(WIDTH)) mul00700105(.x(x_105), .z(tmp00_105_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700106(.x(x_106), .z(tmp00_106_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700107(.x(x_107), .z(tmp00_107_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700108(.x(x_108), .z(tmp00_108_70));
	booth_0002 #(.WIDTH(WIDTH)) mul00700109(.x(x_109), .z(tmp00_109_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700110(.x(x_110), .z(tmp00_110_70));
	booth__012 #(.WIDTH(WIDTH)) mul00700111(.x(x_111), .z(tmp00_111_70));
	booth__006 #(.WIDTH(WIDTH)) mul00700112(.x(x_112), .z(tmp00_112_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700113(.x(x_113), .z(tmp00_113_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700114(.x(x_114), .z(tmp00_114_70));
	booth__010 #(.WIDTH(WIDTH)) mul00700115(.x(x_115), .z(tmp00_115_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700116(.x(x_116), .z(tmp00_116_70));
	booth_0010 #(.WIDTH(WIDTH)) mul00700117(.x(x_117), .z(tmp00_117_70));
	booth__004 #(.WIDTH(WIDTH)) mul00700118(.x(x_118), .z(tmp00_118_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700119(.x(x_119), .z(tmp00_119_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700120(.x(x_120), .z(tmp00_120_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700121(.x(x_121), .z(tmp00_121_70));
	booth__006 #(.WIDTH(WIDTH)) mul00700122(.x(x_122), .z(tmp00_122_70));
	booth__008 #(.WIDTH(WIDTH)) mul00700123(.x(x_123), .z(tmp00_123_70));
	booth_0008 #(.WIDTH(WIDTH)) mul00700124(.x(x_124), .z(tmp00_124_70));
	booth_0002 #(.WIDTH(WIDTH)) mul00700125(.x(x_125), .z(tmp00_125_70));
	booth_0000 #(.WIDTH(WIDTH)) mul00700126(.x(x_126), .z(tmp00_126_70));
	booth__010 #(.WIDTH(WIDTH)) mul00700127(.x(x_127), .z(tmp00_127_70));
	booth__008 #(.WIDTH(WIDTH)) mul00710000(.x(x_0), .z(tmp00_0_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710001(.x(x_1), .z(tmp00_1_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710002(.x(x_2), .z(tmp00_2_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710003(.x(x_3), .z(tmp00_3_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710004(.x(x_4), .z(tmp00_4_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710005(.x(x_5), .z(tmp00_5_71));
	booth_0012 #(.WIDTH(WIDTH)) mul00710006(.x(x_6), .z(tmp00_6_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710007(.x(x_7), .z(tmp00_7_71));
	booth_0002 #(.WIDTH(WIDTH)) mul00710008(.x(x_8), .z(tmp00_8_71));
	booth_0010 #(.WIDTH(WIDTH)) mul00710009(.x(x_9), .z(tmp00_9_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710010(.x(x_10), .z(tmp00_10_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710011(.x(x_11), .z(tmp00_11_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710012(.x(x_12), .z(tmp00_12_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710013(.x(x_13), .z(tmp00_13_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710014(.x(x_14), .z(tmp00_14_71));
	booth_0012 #(.WIDTH(WIDTH)) mul00710015(.x(x_15), .z(tmp00_15_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710016(.x(x_16), .z(tmp00_16_71));
	booth__002 #(.WIDTH(WIDTH)) mul00710017(.x(x_17), .z(tmp00_17_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710018(.x(x_18), .z(tmp00_18_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710019(.x(x_19), .z(tmp00_19_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710020(.x(x_20), .z(tmp00_20_71));
	booth__006 #(.WIDTH(WIDTH)) mul00710021(.x(x_21), .z(tmp00_21_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710022(.x(x_22), .z(tmp00_22_71));
	booth_0016 #(.WIDTH(WIDTH)) mul00710023(.x(x_23), .z(tmp00_23_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710024(.x(x_24), .z(tmp00_24_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710025(.x(x_25), .z(tmp00_25_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710026(.x(x_26), .z(tmp00_26_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710027(.x(x_27), .z(tmp00_27_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710028(.x(x_28), .z(tmp00_28_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710029(.x(x_29), .z(tmp00_29_71));
	booth__006 #(.WIDTH(WIDTH)) mul00710030(.x(x_30), .z(tmp00_30_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710031(.x(x_31), .z(tmp00_31_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710032(.x(x_32), .z(tmp00_32_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710033(.x(x_33), .z(tmp00_33_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710034(.x(x_34), .z(tmp00_34_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710035(.x(x_35), .z(tmp00_35_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710036(.x(x_36), .z(tmp00_36_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710037(.x(x_37), .z(tmp00_37_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710038(.x(x_38), .z(tmp00_38_71));
	booth__016 #(.WIDTH(WIDTH)) mul00710039(.x(x_39), .z(tmp00_39_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710040(.x(x_40), .z(tmp00_40_71));
	booth_0002 #(.WIDTH(WIDTH)) mul00710041(.x(x_41), .z(tmp00_41_71));
	booth__012 #(.WIDTH(WIDTH)) mul00710042(.x(x_42), .z(tmp00_42_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710043(.x(x_43), .z(tmp00_43_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710044(.x(x_44), .z(tmp00_44_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710045(.x(x_45), .z(tmp00_45_71));
	booth__012 #(.WIDTH(WIDTH)) mul00710046(.x(x_46), .z(tmp00_46_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710047(.x(x_47), .z(tmp00_47_71));
	booth__006 #(.WIDTH(WIDTH)) mul00710048(.x(x_48), .z(tmp00_48_71));
	booth__006 #(.WIDTH(WIDTH)) mul00710049(.x(x_49), .z(tmp00_49_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710050(.x(x_50), .z(tmp00_50_71));
	booth__012 #(.WIDTH(WIDTH)) mul00710051(.x(x_51), .z(tmp00_51_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710052(.x(x_52), .z(tmp00_52_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710053(.x(x_53), .z(tmp00_53_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710054(.x(x_54), .z(tmp00_54_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710055(.x(x_55), .z(tmp00_55_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710056(.x(x_56), .z(tmp00_56_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710057(.x(x_57), .z(tmp00_57_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710058(.x(x_58), .z(tmp00_58_71));
	booth_0002 #(.WIDTH(WIDTH)) mul00710059(.x(x_59), .z(tmp00_59_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710060(.x(x_60), .z(tmp00_60_71));
	booth__006 #(.WIDTH(WIDTH)) mul00710061(.x(x_61), .z(tmp00_61_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710062(.x(x_62), .z(tmp00_62_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710063(.x(x_63), .z(tmp00_63_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710064(.x(x_64), .z(tmp00_64_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710065(.x(x_65), .z(tmp00_65_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710066(.x(x_66), .z(tmp00_66_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710067(.x(x_67), .z(tmp00_67_71));
	booth__010 #(.WIDTH(WIDTH)) mul00710068(.x(x_68), .z(tmp00_68_71));
	booth_0012 #(.WIDTH(WIDTH)) mul00710069(.x(x_69), .z(tmp00_69_71));
	booth__006 #(.WIDTH(WIDTH)) mul00710070(.x(x_70), .z(tmp00_70_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710071(.x(x_71), .z(tmp00_71_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710072(.x(x_72), .z(tmp00_72_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710073(.x(x_73), .z(tmp00_73_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710074(.x(x_74), .z(tmp00_74_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710075(.x(x_75), .z(tmp00_75_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710076(.x(x_76), .z(tmp00_76_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710077(.x(x_77), .z(tmp00_77_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710078(.x(x_78), .z(tmp00_78_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710079(.x(x_79), .z(tmp00_79_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710080(.x(x_80), .z(tmp00_80_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710081(.x(x_81), .z(tmp00_81_71));
	booth_0010 #(.WIDTH(WIDTH)) mul00710082(.x(x_82), .z(tmp00_82_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710083(.x(x_83), .z(tmp00_83_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710084(.x(x_84), .z(tmp00_84_71));
	booth__012 #(.WIDTH(WIDTH)) mul00710085(.x(x_85), .z(tmp00_85_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710086(.x(x_86), .z(tmp00_86_71));
	booth_0016 #(.WIDTH(WIDTH)) mul00710087(.x(x_87), .z(tmp00_87_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710088(.x(x_88), .z(tmp00_88_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710089(.x(x_89), .z(tmp00_89_71));
	booth__016 #(.WIDTH(WIDTH)) mul00710090(.x(x_90), .z(tmp00_90_71));
	booth__012 #(.WIDTH(WIDTH)) mul00710091(.x(x_91), .z(tmp00_91_71));
	booth_0006 #(.WIDTH(WIDTH)) mul00710092(.x(x_92), .z(tmp00_92_71));
	booth__006 #(.WIDTH(WIDTH)) mul00710093(.x(x_93), .z(tmp00_93_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710094(.x(x_94), .z(tmp00_94_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710095(.x(x_95), .z(tmp00_95_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710096(.x(x_96), .z(tmp00_96_71));
	booth__006 #(.WIDTH(WIDTH)) mul00710097(.x(x_97), .z(tmp00_97_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710098(.x(x_98), .z(tmp00_98_71));
	booth_0012 #(.WIDTH(WIDTH)) mul00710099(.x(x_99), .z(tmp00_99_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710100(.x(x_100), .z(tmp00_100_71));
	booth__010 #(.WIDTH(WIDTH)) mul00710101(.x(x_101), .z(tmp00_101_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710102(.x(x_102), .z(tmp00_102_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710103(.x(x_103), .z(tmp00_103_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710104(.x(x_104), .z(tmp00_104_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710105(.x(x_105), .z(tmp00_105_71));
	booth_0006 #(.WIDTH(WIDTH)) mul00710106(.x(x_106), .z(tmp00_106_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710107(.x(x_107), .z(tmp00_107_71));
	booth_0004 #(.WIDTH(WIDTH)) mul00710108(.x(x_108), .z(tmp00_108_71));
	booth_0012 #(.WIDTH(WIDTH)) mul00710109(.x(x_109), .z(tmp00_109_71));
	booth_0014 #(.WIDTH(WIDTH)) mul00710110(.x(x_110), .z(tmp00_110_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710111(.x(x_111), .z(tmp00_111_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710112(.x(x_112), .z(tmp00_112_71));
	booth_0016 #(.WIDTH(WIDTH)) mul00710113(.x(x_113), .z(tmp00_113_71));
	booth_0010 #(.WIDTH(WIDTH)) mul00710114(.x(x_114), .z(tmp00_114_71));
	booth_0012 #(.WIDTH(WIDTH)) mul00710115(.x(x_115), .z(tmp00_115_71));
	booth__012 #(.WIDTH(WIDTH)) mul00710116(.x(x_116), .z(tmp00_116_71));
	booth_0008 #(.WIDTH(WIDTH)) mul00710117(.x(x_117), .z(tmp00_117_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710118(.x(x_118), .z(tmp00_118_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710119(.x(x_119), .z(tmp00_119_71));
	booth_0016 #(.WIDTH(WIDTH)) mul00710120(.x(x_120), .z(tmp00_120_71));
	booth_0016 #(.WIDTH(WIDTH)) mul00710121(.x(x_121), .z(tmp00_121_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710122(.x(x_122), .z(tmp00_122_71));
	booth__010 #(.WIDTH(WIDTH)) mul00710123(.x(x_123), .z(tmp00_123_71));
	booth_0000 #(.WIDTH(WIDTH)) mul00710124(.x(x_124), .z(tmp00_124_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710125(.x(x_125), .z(tmp00_125_71));
	booth__008 #(.WIDTH(WIDTH)) mul00710126(.x(x_126), .z(tmp00_126_71));
	booth__004 #(.WIDTH(WIDTH)) mul00710127(.x(x_127), .z(tmp00_127_71));
	booth_0002 #(.WIDTH(WIDTH)) mul00720000(.x(x_0), .z(tmp00_0_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720001(.x(x_1), .z(tmp00_1_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720002(.x(x_2), .z(tmp00_2_72));
	booth__002 #(.WIDTH(WIDTH)) mul00720003(.x(x_3), .z(tmp00_3_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720004(.x(x_4), .z(tmp00_4_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720005(.x(x_5), .z(tmp00_5_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720006(.x(x_6), .z(tmp00_6_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720007(.x(x_7), .z(tmp00_7_72));
	booth_0010 #(.WIDTH(WIDTH)) mul00720008(.x(x_8), .z(tmp00_8_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720009(.x(x_9), .z(tmp00_9_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720010(.x(x_10), .z(tmp00_10_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720011(.x(x_11), .z(tmp00_11_72));
	booth__002 #(.WIDTH(WIDTH)) mul00720012(.x(x_12), .z(tmp00_12_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720013(.x(x_13), .z(tmp00_13_72));
	booth_0012 #(.WIDTH(WIDTH)) mul00720014(.x(x_14), .z(tmp00_14_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720015(.x(x_15), .z(tmp00_15_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720016(.x(x_16), .z(tmp00_16_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720017(.x(x_17), .z(tmp00_17_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720018(.x(x_18), .z(tmp00_18_72));
	booth__016 #(.WIDTH(WIDTH)) mul00720019(.x(x_19), .z(tmp00_19_72));
	booth_0006 #(.WIDTH(WIDTH)) mul00720020(.x(x_20), .z(tmp00_20_72));
	booth__010 #(.WIDTH(WIDTH)) mul00720021(.x(x_21), .z(tmp00_21_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720022(.x(x_22), .z(tmp00_22_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720023(.x(x_23), .z(tmp00_23_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720024(.x(x_24), .z(tmp00_24_72));
	booth_0012 #(.WIDTH(WIDTH)) mul00720025(.x(x_25), .z(tmp00_25_72));
	booth__010 #(.WIDTH(WIDTH)) mul00720026(.x(x_26), .z(tmp00_26_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720027(.x(x_27), .z(tmp00_27_72));
	booth_0016 #(.WIDTH(WIDTH)) mul00720028(.x(x_28), .z(tmp00_28_72));
	booth_0002 #(.WIDTH(WIDTH)) mul00720029(.x(x_29), .z(tmp00_29_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720030(.x(x_30), .z(tmp00_30_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720031(.x(x_31), .z(tmp00_31_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720032(.x(x_32), .z(tmp00_32_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720033(.x(x_33), .z(tmp00_33_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720034(.x(x_34), .z(tmp00_34_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720035(.x(x_35), .z(tmp00_35_72));
	booth_0010 #(.WIDTH(WIDTH)) mul00720036(.x(x_36), .z(tmp00_36_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720037(.x(x_37), .z(tmp00_37_72));
	booth_0020 #(.WIDTH(WIDTH)) mul00720038(.x(x_38), .z(tmp00_38_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720039(.x(x_39), .z(tmp00_39_72));
	booth__016 #(.WIDTH(WIDTH)) mul00720040(.x(x_40), .z(tmp00_40_72));
	booth_0016 #(.WIDTH(WIDTH)) mul00720041(.x(x_41), .z(tmp00_41_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720042(.x(x_42), .z(tmp00_42_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720043(.x(x_43), .z(tmp00_43_72));
	booth_0012 #(.WIDTH(WIDTH)) mul00720044(.x(x_44), .z(tmp00_44_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720045(.x(x_45), .z(tmp00_45_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720046(.x(x_46), .z(tmp00_46_72));
	booth__012 #(.WIDTH(WIDTH)) mul00720047(.x(x_47), .z(tmp00_47_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720048(.x(x_48), .z(tmp00_48_72));
	booth_0002 #(.WIDTH(WIDTH)) mul00720049(.x(x_49), .z(tmp00_49_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720050(.x(x_50), .z(tmp00_50_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720051(.x(x_51), .z(tmp00_51_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720052(.x(x_52), .z(tmp00_52_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720053(.x(x_53), .z(tmp00_53_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720054(.x(x_54), .z(tmp00_54_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720055(.x(x_55), .z(tmp00_55_72));
	booth_0012 #(.WIDTH(WIDTH)) mul00720056(.x(x_56), .z(tmp00_56_72));
	booth__012 #(.WIDTH(WIDTH)) mul00720057(.x(x_57), .z(tmp00_57_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720058(.x(x_58), .z(tmp00_58_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720059(.x(x_59), .z(tmp00_59_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720060(.x(x_60), .z(tmp00_60_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720061(.x(x_61), .z(tmp00_61_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720062(.x(x_62), .z(tmp00_62_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720063(.x(x_63), .z(tmp00_63_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720064(.x(x_64), .z(tmp00_64_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720065(.x(x_65), .z(tmp00_65_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720066(.x(x_66), .z(tmp00_66_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720067(.x(x_67), .z(tmp00_67_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720068(.x(x_68), .z(tmp00_68_72));
	booth_0002 #(.WIDTH(WIDTH)) mul00720069(.x(x_69), .z(tmp00_69_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720070(.x(x_70), .z(tmp00_70_72));
	booth_0006 #(.WIDTH(WIDTH)) mul00720071(.x(x_71), .z(tmp00_71_72));
	booth__016 #(.WIDTH(WIDTH)) mul00720072(.x(x_72), .z(tmp00_72_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720073(.x(x_73), .z(tmp00_73_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720074(.x(x_74), .z(tmp00_74_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720075(.x(x_75), .z(tmp00_75_72));
	booth__006 #(.WIDTH(WIDTH)) mul00720076(.x(x_76), .z(tmp00_76_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720077(.x(x_77), .z(tmp00_77_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720078(.x(x_78), .z(tmp00_78_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720079(.x(x_79), .z(tmp00_79_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720080(.x(x_80), .z(tmp00_80_72));
	booth_0014 #(.WIDTH(WIDTH)) mul00720081(.x(x_81), .z(tmp00_81_72));
	booth_0006 #(.WIDTH(WIDTH)) mul00720082(.x(x_82), .z(tmp00_82_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720083(.x(x_83), .z(tmp00_83_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720084(.x(x_84), .z(tmp00_84_72));
	booth__012 #(.WIDTH(WIDTH)) mul00720085(.x(x_85), .z(tmp00_85_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720086(.x(x_86), .z(tmp00_86_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720087(.x(x_87), .z(tmp00_87_72));
	booth_0010 #(.WIDTH(WIDTH)) mul00720088(.x(x_88), .z(tmp00_88_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720089(.x(x_89), .z(tmp00_89_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720090(.x(x_90), .z(tmp00_90_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720091(.x(x_91), .z(tmp00_91_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720092(.x(x_92), .z(tmp00_92_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720093(.x(x_93), .z(tmp00_93_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720094(.x(x_94), .z(tmp00_94_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720095(.x(x_95), .z(tmp00_95_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720096(.x(x_96), .z(tmp00_96_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720097(.x(x_97), .z(tmp00_97_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720098(.x(x_98), .z(tmp00_98_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720099(.x(x_99), .z(tmp00_99_72));
	booth__012 #(.WIDTH(WIDTH)) mul00720100(.x(x_100), .z(tmp00_100_72));
	booth_0010 #(.WIDTH(WIDTH)) mul00720101(.x(x_101), .z(tmp00_101_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720102(.x(x_102), .z(tmp00_102_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720103(.x(x_103), .z(tmp00_103_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720104(.x(x_104), .z(tmp00_104_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720105(.x(x_105), .z(tmp00_105_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720106(.x(x_106), .z(tmp00_106_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720107(.x(x_107), .z(tmp00_107_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720108(.x(x_108), .z(tmp00_108_72));
	booth__016 #(.WIDTH(WIDTH)) mul00720109(.x(x_109), .z(tmp00_109_72));
	booth_0012 #(.WIDTH(WIDTH)) mul00720110(.x(x_110), .z(tmp00_110_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720111(.x(x_111), .z(tmp00_111_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720112(.x(x_112), .z(tmp00_112_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720113(.x(x_113), .z(tmp00_113_72));
	booth__016 #(.WIDTH(WIDTH)) mul00720114(.x(x_114), .z(tmp00_114_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720115(.x(x_115), .z(tmp00_115_72));
	booth_0004 #(.WIDTH(WIDTH)) mul00720116(.x(x_116), .z(tmp00_116_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720117(.x(x_117), .z(tmp00_117_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720118(.x(x_118), .z(tmp00_118_72));
	booth_0020 #(.WIDTH(WIDTH)) mul00720119(.x(x_119), .z(tmp00_119_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720120(.x(x_120), .z(tmp00_120_72));
	booth__004 #(.WIDTH(WIDTH)) mul00720121(.x(x_121), .z(tmp00_121_72));
	booth__010 #(.WIDTH(WIDTH)) mul00720122(.x(x_122), .z(tmp00_122_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00720123(.x(x_123), .z(tmp00_123_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720124(.x(x_124), .z(tmp00_124_72));
	booth__008 #(.WIDTH(WIDTH)) mul00720125(.x(x_125), .z(tmp00_125_72));
	booth_0016 #(.WIDTH(WIDTH)) mul00720126(.x(x_126), .z(tmp00_126_72));
	booth_0008 #(.WIDTH(WIDTH)) mul00720127(.x(x_127), .z(tmp00_127_72));
	booth_0000 #(.WIDTH(WIDTH)) mul00730000(.x(x_0), .z(tmp00_0_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730001(.x(x_1), .z(tmp00_1_73));
	booth__006 #(.WIDTH(WIDTH)) mul00730002(.x(x_2), .z(tmp00_2_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730003(.x(x_3), .z(tmp00_3_73));
	booth_0010 #(.WIDTH(WIDTH)) mul00730004(.x(x_4), .z(tmp00_4_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730005(.x(x_5), .z(tmp00_5_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730006(.x(x_6), .z(tmp00_6_73));
	booth__002 #(.WIDTH(WIDTH)) mul00730007(.x(x_7), .z(tmp00_7_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730008(.x(x_8), .z(tmp00_8_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730009(.x(x_9), .z(tmp00_9_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730010(.x(x_10), .z(tmp00_10_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730011(.x(x_11), .z(tmp00_11_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730012(.x(x_12), .z(tmp00_12_73));
	booth_0012 #(.WIDTH(WIDTH)) mul00730013(.x(x_13), .z(tmp00_13_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730014(.x(x_14), .z(tmp00_14_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730015(.x(x_15), .z(tmp00_15_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730016(.x(x_16), .z(tmp00_16_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730017(.x(x_17), .z(tmp00_17_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730018(.x(x_18), .z(tmp00_18_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730019(.x(x_19), .z(tmp00_19_73));
	booth_0006 #(.WIDTH(WIDTH)) mul00730020(.x(x_20), .z(tmp00_20_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730021(.x(x_21), .z(tmp00_21_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730022(.x(x_22), .z(tmp00_22_73));
	booth_0012 #(.WIDTH(WIDTH)) mul00730023(.x(x_23), .z(tmp00_23_73));
	booth_0010 #(.WIDTH(WIDTH)) mul00730024(.x(x_24), .z(tmp00_24_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730025(.x(x_25), .z(tmp00_25_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730026(.x(x_26), .z(tmp00_26_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730027(.x(x_27), .z(tmp00_27_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730028(.x(x_28), .z(tmp00_28_73));
	booth__002 #(.WIDTH(WIDTH)) mul00730029(.x(x_29), .z(tmp00_29_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730030(.x(x_30), .z(tmp00_30_73));
	booth__006 #(.WIDTH(WIDTH)) mul00730031(.x(x_31), .z(tmp00_31_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730032(.x(x_32), .z(tmp00_32_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730033(.x(x_33), .z(tmp00_33_73));
	booth_0006 #(.WIDTH(WIDTH)) mul00730034(.x(x_34), .z(tmp00_34_73));
	booth__006 #(.WIDTH(WIDTH)) mul00730035(.x(x_35), .z(tmp00_35_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730036(.x(x_36), .z(tmp00_36_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730037(.x(x_37), .z(tmp00_37_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730038(.x(x_38), .z(tmp00_38_73));
	booth__006 #(.WIDTH(WIDTH)) mul00730039(.x(x_39), .z(tmp00_39_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730040(.x(x_40), .z(tmp00_40_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730041(.x(x_41), .z(tmp00_41_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730042(.x(x_42), .z(tmp00_42_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730043(.x(x_43), .z(tmp00_43_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730044(.x(x_44), .z(tmp00_44_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730045(.x(x_45), .z(tmp00_45_73));
	booth__006 #(.WIDTH(WIDTH)) mul00730046(.x(x_46), .z(tmp00_46_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730047(.x(x_47), .z(tmp00_47_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730048(.x(x_48), .z(tmp00_48_73));
	booth__012 #(.WIDTH(WIDTH)) mul00730049(.x(x_49), .z(tmp00_49_73));
	booth__004 #(.WIDTH(WIDTH)) mul00730050(.x(x_50), .z(tmp00_50_73));
	booth__004 #(.WIDTH(WIDTH)) mul00730051(.x(x_51), .z(tmp00_51_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730052(.x(x_52), .z(tmp00_52_73));
	booth__004 #(.WIDTH(WIDTH)) mul00730053(.x(x_53), .z(tmp00_53_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730054(.x(x_54), .z(tmp00_54_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730055(.x(x_55), .z(tmp00_55_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730056(.x(x_56), .z(tmp00_56_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730057(.x(x_57), .z(tmp00_57_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730058(.x(x_58), .z(tmp00_58_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730059(.x(x_59), .z(tmp00_59_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730060(.x(x_60), .z(tmp00_60_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730061(.x(x_61), .z(tmp00_61_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730062(.x(x_62), .z(tmp00_62_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730063(.x(x_63), .z(tmp00_63_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730064(.x(x_64), .z(tmp00_64_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730065(.x(x_65), .z(tmp00_65_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730066(.x(x_66), .z(tmp00_66_73));
	booth__006 #(.WIDTH(WIDTH)) mul00730067(.x(x_67), .z(tmp00_67_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730068(.x(x_68), .z(tmp00_68_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730069(.x(x_69), .z(tmp00_69_73));
	booth_0010 #(.WIDTH(WIDTH)) mul00730070(.x(x_70), .z(tmp00_70_73));
	booth__012 #(.WIDTH(WIDTH)) mul00730071(.x(x_71), .z(tmp00_71_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730072(.x(x_72), .z(tmp00_72_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730073(.x(x_73), .z(tmp00_73_73));
	booth__004 #(.WIDTH(WIDTH)) mul00730074(.x(x_74), .z(tmp00_74_73));
	booth__012 #(.WIDTH(WIDTH)) mul00730075(.x(x_75), .z(tmp00_75_73));
	booth__002 #(.WIDTH(WIDTH)) mul00730076(.x(x_76), .z(tmp00_76_73));
	booth_0010 #(.WIDTH(WIDTH)) mul00730077(.x(x_77), .z(tmp00_77_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730078(.x(x_78), .z(tmp00_78_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730079(.x(x_79), .z(tmp00_79_73));
	booth__016 #(.WIDTH(WIDTH)) mul00730080(.x(x_80), .z(tmp00_80_73));
	booth_0010 #(.WIDTH(WIDTH)) mul00730081(.x(x_81), .z(tmp00_81_73));
	booth_0014 #(.WIDTH(WIDTH)) mul00730082(.x(x_82), .z(tmp00_82_73));
	booth_0006 #(.WIDTH(WIDTH)) mul00730083(.x(x_83), .z(tmp00_83_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730084(.x(x_84), .z(tmp00_84_73));
	booth_0012 #(.WIDTH(WIDTH)) mul00730085(.x(x_85), .z(tmp00_85_73));
	booth_0006 #(.WIDTH(WIDTH)) mul00730086(.x(x_86), .z(tmp00_86_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730087(.x(x_87), .z(tmp00_87_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730088(.x(x_88), .z(tmp00_88_73));
	booth_0010 #(.WIDTH(WIDTH)) mul00730089(.x(x_89), .z(tmp00_89_73));
	booth_0010 #(.WIDTH(WIDTH)) mul00730090(.x(x_90), .z(tmp00_90_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730091(.x(x_91), .z(tmp00_91_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730092(.x(x_92), .z(tmp00_92_73));
	booth__004 #(.WIDTH(WIDTH)) mul00730093(.x(x_93), .z(tmp00_93_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730094(.x(x_94), .z(tmp00_94_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730095(.x(x_95), .z(tmp00_95_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730096(.x(x_96), .z(tmp00_96_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730097(.x(x_97), .z(tmp00_97_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730098(.x(x_98), .z(tmp00_98_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730099(.x(x_99), .z(tmp00_99_73));
	booth_0006 #(.WIDTH(WIDTH)) mul00730100(.x(x_100), .z(tmp00_100_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730101(.x(x_101), .z(tmp00_101_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730102(.x(x_102), .z(tmp00_102_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730103(.x(x_103), .z(tmp00_103_73));
	booth_0012 #(.WIDTH(WIDTH)) mul00730104(.x(x_104), .z(tmp00_104_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730105(.x(x_105), .z(tmp00_105_73));
	booth__010 #(.WIDTH(WIDTH)) mul00730106(.x(x_106), .z(tmp00_106_73));
	booth_0004 #(.WIDTH(WIDTH)) mul00730107(.x(x_107), .z(tmp00_107_73));
	booth_0008 #(.WIDTH(WIDTH)) mul00730108(.x(x_108), .z(tmp00_108_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730109(.x(x_109), .z(tmp00_109_73));
	booth_0016 #(.WIDTH(WIDTH)) mul00730110(.x(x_110), .z(tmp00_110_73));
	booth__006 #(.WIDTH(WIDTH)) mul00730111(.x(x_111), .z(tmp00_111_73));
	booth_0012 #(.WIDTH(WIDTH)) mul00730112(.x(x_112), .z(tmp00_112_73));
	booth__002 #(.WIDTH(WIDTH)) mul00730113(.x(x_113), .z(tmp00_113_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730114(.x(x_114), .z(tmp00_114_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730115(.x(x_115), .z(tmp00_115_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730116(.x(x_116), .z(tmp00_116_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730117(.x(x_117), .z(tmp00_117_73));
	booth__004 #(.WIDTH(WIDTH)) mul00730118(.x(x_118), .z(tmp00_118_73));
	booth_0012 #(.WIDTH(WIDTH)) mul00730119(.x(x_119), .z(tmp00_119_73));
	booth_0020 #(.WIDTH(WIDTH)) mul00730120(.x(x_120), .z(tmp00_120_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730121(.x(x_121), .z(tmp00_121_73));
	booth__004 #(.WIDTH(WIDTH)) mul00730122(.x(x_122), .z(tmp00_122_73));
	booth__008 #(.WIDTH(WIDTH)) mul00730123(.x(x_123), .z(tmp00_123_73));
	booth_0002 #(.WIDTH(WIDTH)) mul00730124(.x(x_124), .z(tmp00_124_73));
	booth_0000 #(.WIDTH(WIDTH)) mul00730125(.x(x_125), .z(tmp00_125_73));
	booth__014 #(.WIDTH(WIDTH)) mul00730126(.x(x_126), .z(tmp00_126_73));
	booth__004 #(.WIDTH(WIDTH)) mul00730127(.x(x_127), .z(tmp00_127_73));
	booth_0010 #(.WIDTH(WIDTH)) mul00740000(.x(x_0), .z(tmp00_0_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740001(.x(x_1), .z(tmp00_1_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740002(.x(x_2), .z(tmp00_2_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740003(.x(x_3), .z(tmp00_3_74));
	booth__012 #(.WIDTH(WIDTH)) mul00740004(.x(x_4), .z(tmp00_4_74));
	booth__006 #(.WIDTH(WIDTH)) mul00740005(.x(x_5), .z(tmp00_5_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740006(.x(x_6), .z(tmp00_6_74));
	booth__006 #(.WIDTH(WIDTH)) mul00740007(.x(x_7), .z(tmp00_7_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740008(.x(x_8), .z(tmp00_8_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740009(.x(x_9), .z(tmp00_9_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740010(.x(x_10), .z(tmp00_10_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740011(.x(x_11), .z(tmp00_11_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740012(.x(x_12), .z(tmp00_12_74));
	booth__010 #(.WIDTH(WIDTH)) mul00740013(.x(x_13), .z(tmp00_13_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740014(.x(x_14), .z(tmp00_14_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740015(.x(x_15), .z(tmp00_15_74));
	booth_0002 #(.WIDTH(WIDTH)) mul00740016(.x(x_16), .z(tmp00_16_74));
	booth_0002 #(.WIDTH(WIDTH)) mul00740017(.x(x_17), .z(tmp00_17_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740018(.x(x_18), .z(tmp00_18_74));
	booth_0002 #(.WIDTH(WIDTH)) mul00740019(.x(x_19), .z(tmp00_19_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740020(.x(x_20), .z(tmp00_20_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740021(.x(x_21), .z(tmp00_21_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740022(.x(x_22), .z(tmp00_22_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740023(.x(x_23), .z(tmp00_23_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740024(.x(x_24), .z(tmp00_24_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740025(.x(x_25), .z(tmp00_25_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740026(.x(x_26), .z(tmp00_26_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740027(.x(x_27), .z(tmp00_27_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740028(.x(x_28), .z(tmp00_28_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740029(.x(x_29), .z(tmp00_29_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740030(.x(x_30), .z(tmp00_30_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740031(.x(x_31), .z(tmp00_31_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740032(.x(x_32), .z(tmp00_32_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740033(.x(x_33), .z(tmp00_33_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740034(.x(x_34), .z(tmp00_34_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740035(.x(x_35), .z(tmp00_35_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740036(.x(x_36), .z(tmp00_36_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740037(.x(x_37), .z(tmp00_37_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740038(.x(x_38), .z(tmp00_38_74));
	booth_0006 #(.WIDTH(WIDTH)) mul00740039(.x(x_39), .z(tmp00_39_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740040(.x(x_40), .z(tmp00_40_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740041(.x(x_41), .z(tmp00_41_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740042(.x(x_42), .z(tmp00_42_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740043(.x(x_43), .z(tmp00_43_74));
	booth__010 #(.WIDTH(WIDTH)) mul00740044(.x(x_44), .z(tmp00_44_74));
	booth_0012 #(.WIDTH(WIDTH)) mul00740045(.x(x_45), .z(tmp00_45_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740046(.x(x_46), .z(tmp00_46_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740047(.x(x_47), .z(tmp00_47_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740048(.x(x_48), .z(tmp00_48_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740049(.x(x_49), .z(tmp00_49_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740050(.x(x_50), .z(tmp00_50_74));
	booth__006 #(.WIDTH(WIDTH)) mul00740051(.x(x_51), .z(tmp00_51_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740052(.x(x_52), .z(tmp00_52_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740053(.x(x_53), .z(tmp00_53_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740054(.x(x_54), .z(tmp00_54_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740055(.x(x_55), .z(tmp00_55_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740056(.x(x_56), .z(tmp00_56_74));
	booth__010 #(.WIDTH(WIDTH)) mul00740057(.x(x_57), .z(tmp00_57_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740058(.x(x_58), .z(tmp00_58_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740059(.x(x_59), .z(tmp00_59_74));
	booth_0006 #(.WIDTH(WIDTH)) mul00740060(.x(x_60), .z(tmp00_60_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740061(.x(x_61), .z(tmp00_61_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740062(.x(x_62), .z(tmp00_62_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740063(.x(x_63), .z(tmp00_63_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740064(.x(x_64), .z(tmp00_64_74));
	booth_0012 #(.WIDTH(WIDTH)) mul00740065(.x(x_65), .z(tmp00_65_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740066(.x(x_66), .z(tmp00_66_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740067(.x(x_67), .z(tmp00_67_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740068(.x(x_68), .z(tmp00_68_74));
	booth__010 #(.WIDTH(WIDTH)) mul00740069(.x(x_69), .z(tmp00_69_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740070(.x(x_70), .z(tmp00_70_74));
	booth_0002 #(.WIDTH(WIDTH)) mul00740071(.x(x_71), .z(tmp00_71_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740072(.x(x_72), .z(tmp00_72_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740073(.x(x_73), .z(tmp00_73_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740074(.x(x_74), .z(tmp00_74_74));
	booth_0006 #(.WIDTH(WIDTH)) mul00740075(.x(x_75), .z(tmp00_75_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740076(.x(x_76), .z(tmp00_76_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740077(.x(x_77), .z(tmp00_77_74));
	booth__012 #(.WIDTH(WIDTH)) mul00740078(.x(x_78), .z(tmp00_78_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740079(.x(x_79), .z(tmp00_79_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740080(.x(x_80), .z(tmp00_80_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740081(.x(x_81), .z(tmp00_81_74));
	booth__010 #(.WIDTH(WIDTH)) mul00740082(.x(x_82), .z(tmp00_82_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740083(.x(x_83), .z(tmp00_83_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740084(.x(x_84), .z(tmp00_84_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740085(.x(x_85), .z(tmp00_85_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740086(.x(x_86), .z(tmp00_86_74));
	booth_0002 #(.WIDTH(WIDTH)) mul00740087(.x(x_87), .z(tmp00_87_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740088(.x(x_88), .z(tmp00_88_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740089(.x(x_89), .z(tmp00_89_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740090(.x(x_90), .z(tmp00_90_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740091(.x(x_91), .z(tmp00_91_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740092(.x(x_92), .z(tmp00_92_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740093(.x(x_93), .z(tmp00_93_74));
	booth_0002 #(.WIDTH(WIDTH)) mul00740094(.x(x_94), .z(tmp00_94_74));
	booth_0012 #(.WIDTH(WIDTH)) mul00740095(.x(x_95), .z(tmp00_95_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740096(.x(x_96), .z(tmp00_96_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740097(.x(x_97), .z(tmp00_97_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740098(.x(x_98), .z(tmp00_98_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740099(.x(x_99), .z(tmp00_99_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740100(.x(x_100), .z(tmp00_100_74));
	booth_0002 #(.WIDTH(WIDTH)) mul00740101(.x(x_101), .z(tmp00_101_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740102(.x(x_102), .z(tmp00_102_74));
	booth__006 #(.WIDTH(WIDTH)) mul00740103(.x(x_103), .z(tmp00_103_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740104(.x(x_104), .z(tmp00_104_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740105(.x(x_105), .z(tmp00_105_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740106(.x(x_106), .z(tmp00_106_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740107(.x(x_107), .z(tmp00_107_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740108(.x(x_108), .z(tmp00_108_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740109(.x(x_109), .z(tmp00_109_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740110(.x(x_110), .z(tmp00_110_74));
	booth_0010 #(.WIDTH(WIDTH)) mul00740111(.x(x_111), .z(tmp00_111_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740112(.x(x_112), .z(tmp00_112_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740113(.x(x_113), .z(tmp00_113_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740114(.x(x_114), .z(tmp00_114_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740115(.x(x_115), .z(tmp00_115_74));
	booth_0008 #(.WIDTH(WIDTH)) mul00740116(.x(x_116), .z(tmp00_116_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740117(.x(x_117), .z(tmp00_117_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740118(.x(x_118), .z(tmp00_118_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740119(.x(x_119), .z(tmp00_119_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740120(.x(x_120), .z(tmp00_120_74));
	booth_0004 #(.WIDTH(WIDTH)) mul00740121(.x(x_121), .z(tmp00_121_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740122(.x(x_122), .z(tmp00_122_74));
	booth__002 #(.WIDTH(WIDTH)) mul00740123(.x(x_123), .z(tmp00_123_74));
	booth_0000 #(.WIDTH(WIDTH)) mul00740124(.x(x_124), .z(tmp00_124_74));
	booth__004 #(.WIDTH(WIDTH)) mul00740125(.x(x_125), .z(tmp00_125_74));
	booth__010 #(.WIDTH(WIDTH)) mul00740126(.x(x_126), .z(tmp00_126_74));
	booth__008 #(.WIDTH(WIDTH)) mul00740127(.x(x_127), .z(tmp00_127_74));
	booth__008 #(.WIDTH(WIDTH)) mul00750000(.x(x_0), .z(tmp00_0_75));
	booth__006 #(.WIDTH(WIDTH)) mul00750001(.x(x_1), .z(tmp00_1_75));
	booth_0012 #(.WIDTH(WIDTH)) mul00750002(.x(x_2), .z(tmp00_2_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750003(.x(x_3), .z(tmp00_3_75));
	booth__002 #(.WIDTH(WIDTH)) mul00750004(.x(x_4), .z(tmp00_4_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750005(.x(x_5), .z(tmp00_5_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750006(.x(x_6), .z(tmp00_6_75));
	booth_0010 #(.WIDTH(WIDTH)) mul00750007(.x(x_7), .z(tmp00_7_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750008(.x(x_8), .z(tmp00_8_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750009(.x(x_9), .z(tmp00_9_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750010(.x(x_10), .z(tmp00_10_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750011(.x(x_11), .z(tmp00_11_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750012(.x(x_12), .z(tmp00_12_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750013(.x(x_13), .z(tmp00_13_75));
	booth_0002 #(.WIDTH(WIDTH)) mul00750014(.x(x_14), .z(tmp00_14_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750015(.x(x_15), .z(tmp00_15_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750016(.x(x_16), .z(tmp00_16_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750017(.x(x_17), .z(tmp00_17_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750018(.x(x_18), .z(tmp00_18_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750019(.x(x_19), .z(tmp00_19_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750020(.x(x_20), .z(tmp00_20_75));
	booth__006 #(.WIDTH(WIDTH)) mul00750021(.x(x_21), .z(tmp00_21_75));
	booth__002 #(.WIDTH(WIDTH)) mul00750022(.x(x_22), .z(tmp00_22_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750023(.x(x_23), .z(tmp00_23_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750024(.x(x_24), .z(tmp00_24_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750025(.x(x_25), .z(tmp00_25_75));
	booth_0010 #(.WIDTH(WIDTH)) mul00750026(.x(x_26), .z(tmp00_26_75));
	booth__010 #(.WIDTH(WIDTH)) mul00750027(.x(x_27), .z(tmp00_27_75));
	booth_0006 #(.WIDTH(WIDTH)) mul00750028(.x(x_28), .z(tmp00_28_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750029(.x(x_29), .z(tmp00_29_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750030(.x(x_30), .z(tmp00_30_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750031(.x(x_31), .z(tmp00_31_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750032(.x(x_32), .z(tmp00_32_75));
	booth_0006 #(.WIDTH(WIDTH)) mul00750033(.x(x_33), .z(tmp00_33_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750034(.x(x_34), .z(tmp00_34_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750035(.x(x_35), .z(tmp00_35_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750036(.x(x_36), .z(tmp00_36_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750037(.x(x_37), .z(tmp00_37_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750038(.x(x_38), .z(tmp00_38_75));
	booth__006 #(.WIDTH(WIDTH)) mul00750039(.x(x_39), .z(tmp00_39_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750040(.x(x_40), .z(tmp00_40_75));
	booth_0002 #(.WIDTH(WIDTH)) mul00750041(.x(x_41), .z(tmp00_41_75));
	booth_0012 #(.WIDTH(WIDTH)) mul00750042(.x(x_42), .z(tmp00_42_75));
	booth__002 #(.WIDTH(WIDTH)) mul00750043(.x(x_43), .z(tmp00_43_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750044(.x(x_44), .z(tmp00_44_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750045(.x(x_45), .z(tmp00_45_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750046(.x(x_46), .z(tmp00_46_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750047(.x(x_47), .z(tmp00_47_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750048(.x(x_48), .z(tmp00_48_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750049(.x(x_49), .z(tmp00_49_75));
	booth__002 #(.WIDTH(WIDTH)) mul00750050(.x(x_50), .z(tmp00_50_75));
	booth_0002 #(.WIDTH(WIDTH)) mul00750051(.x(x_51), .z(tmp00_51_75));
	booth_0002 #(.WIDTH(WIDTH)) mul00750052(.x(x_52), .z(tmp00_52_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750053(.x(x_53), .z(tmp00_53_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750054(.x(x_54), .z(tmp00_54_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750055(.x(x_55), .z(tmp00_55_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750056(.x(x_56), .z(tmp00_56_75));
	booth_0002 #(.WIDTH(WIDTH)) mul00750057(.x(x_57), .z(tmp00_57_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750058(.x(x_58), .z(tmp00_58_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750059(.x(x_59), .z(tmp00_59_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750060(.x(x_60), .z(tmp00_60_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750061(.x(x_61), .z(tmp00_61_75));
	booth__010 #(.WIDTH(WIDTH)) mul00750062(.x(x_62), .z(tmp00_62_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750063(.x(x_63), .z(tmp00_63_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750064(.x(x_64), .z(tmp00_64_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750065(.x(x_65), .z(tmp00_65_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750066(.x(x_66), .z(tmp00_66_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750067(.x(x_67), .z(tmp00_67_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750068(.x(x_68), .z(tmp00_68_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750069(.x(x_69), .z(tmp00_69_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750070(.x(x_70), .z(tmp00_70_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750071(.x(x_71), .z(tmp00_71_75));
	booth_0006 #(.WIDTH(WIDTH)) mul00750072(.x(x_72), .z(tmp00_72_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750073(.x(x_73), .z(tmp00_73_75));
	booth_0010 #(.WIDTH(WIDTH)) mul00750074(.x(x_74), .z(tmp00_74_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750075(.x(x_75), .z(tmp00_75_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750076(.x(x_76), .z(tmp00_76_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750077(.x(x_77), .z(tmp00_77_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750078(.x(x_78), .z(tmp00_78_75));
	booth__006 #(.WIDTH(WIDTH)) mul00750079(.x(x_79), .z(tmp00_79_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750080(.x(x_80), .z(tmp00_80_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750081(.x(x_81), .z(tmp00_81_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750082(.x(x_82), .z(tmp00_82_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750083(.x(x_83), .z(tmp00_83_75));
	booth_0010 #(.WIDTH(WIDTH)) mul00750084(.x(x_84), .z(tmp00_84_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750085(.x(x_85), .z(tmp00_85_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750086(.x(x_86), .z(tmp00_86_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750087(.x(x_87), .z(tmp00_87_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750088(.x(x_88), .z(tmp00_88_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750089(.x(x_89), .z(tmp00_89_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750090(.x(x_90), .z(tmp00_90_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750091(.x(x_91), .z(tmp00_91_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750092(.x(x_92), .z(tmp00_92_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750093(.x(x_93), .z(tmp00_93_75));
	booth__006 #(.WIDTH(WIDTH)) mul00750094(.x(x_94), .z(tmp00_94_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750095(.x(x_95), .z(tmp00_95_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750096(.x(x_96), .z(tmp00_96_75));
	booth_0010 #(.WIDTH(WIDTH)) mul00750097(.x(x_97), .z(tmp00_97_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750098(.x(x_98), .z(tmp00_98_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750099(.x(x_99), .z(tmp00_99_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750100(.x(x_100), .z(tmp00_100_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750101(.x(x_101), .z(tmp00_101_75));
	booth__010 #(.WIDTH(WIDTH)) mul00750102(.x(x_102), .z(tmp00_102_75));
	booth_0010 #(.WIDTH(WIDTH)) mul00750103(.x(x_103), .z(tmp00_103_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750104(.x(x_104), .z(tmp00_104_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750105(.x(x_105), .z(tmp00_105_75));
	booth__006 #(.WIDTH(WIDTH)) mul00750106(.x(x_106), .z(tmp00_106_75));
	booth_0010 #(.WIDTH(WIDTH)) mul00750107(.x(x_107), .z(tmp00_107_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750108(.x(x_108), .z(tmp00_108_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750109(.x(x_109), .z(tmp00_109_75));
	booth_0002 #(.WIDTH(WIDTH)) mul00750110(.x(x_110), .z(tmp00_110_75));
	booth__012 #(.WIDTH(WIDTH)) mul00750111(.x(x_111), .z(tmp00_111_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750112(.x(x_112), .z(tmp00_112_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750113(.x(x_113), .z(tmp00_113_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750114(.x(x_114), .z(tmp00_114_75));
	booth_0002 #(.WIDTH(WIDTH)) mul00750115(.x(x_115), .z(tmp00_115_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750116(.x(x_116), .z(tmp00_116_75));
	booth_0008 #(.WIDTH(WIDTH)) mul00750117(.x(x_117), .z(tmp00_117_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750118(.x(x_118), .z(tmp00_118_75));
	booth_0010 #(.WIDTH(WIDTH)) mul00750119(.x(x_119), .z(tmp00_119_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750120(.x(x_120), .z(tmp00_120_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750121(.x(x_121), .z(tmp00_121_75));
	booth_0004 #(.WIDTH(WIDTH)) mul00750122(.x(x_122), .z(tmp00_122_75));
	booth_0006 #(.WIDTH(WIDTH)) mul00750123(.x(x_123), .z(tmp00_123_75));
	booth__008 #(.WIDTH(WIDTH)) mul00750124(.x(x_124), .z(tmp00_124_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750125(.x(x_125), .z(tmp00_125_75));
	booth__004 #(.WIDTH(WIDTH)) mul00750126(.x(x_126), .z(tmp00_126_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00750127(.x(x_127), .z(tmp00_127_75));
	booth_0000 #(.WIDTH(WIDTH)) mul00760000(.x(x_0), .z(tmp00_0_76));
	booth_0006 #(.WIDTH(WIDTH)) mul00760001(.x(x_1), .z(tmp00_1_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760002(.x(x_2), .z(tmp00_2_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760003(.x(x_3), .z(tmp00_3_76));
	booth__014 #(.WIDTH(WIDTH)) mul00760004(.x(x_4), .z(tmp00_4_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760005(.x(x_5), .z(tmp00_5_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760006(.x(x_6), .z(tmp00_6_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760007(.x(x_7), .z(tmp00_7_76));
	booth_0002 #(.WIDTH(WIDTH)) mul00760008(.x(x_8), .z(tmp00_8_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760009(.x(x_9), .z(tmp00_9_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760010(.x(x_10), .z(tmp00_10_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760011(.x(x_11), .z(tmp00_11_76));
	booth__010 #(.WIDTH(WIDTH)) mul00760012(.x(x_12), .z(tmp00_12_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760013(.x(x_13), .z(tmp00_13_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760014(.x(x_14), .z(tmp00_14_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760015(.x(x_15), .z(tmp00_15_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760016(.x(x_16), .z(tmp00_16_76));
	booth_0006 #(.WIDTH(WIDTH)) mul00760017(.x(x_17), .z(tmp00_17_76));
	booth__006 #(.WIDTH(WIDTH)) mul00760018(.x(x_18), .z(tmp00_18_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760019(.x(x_19), .z(tmp00_19_76));
	booth__012 #(.WIDTH(WIDTH)) mul00760020(.x(x_20), .z(tmp00_20_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760021(.x(x_21), .z(tmp00_21_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760022(.x(x_22), .z(tmp00_22_76));
	booth_0006 #(.WIDTH(WIDTH)) mul00760023(.x(x_23), .z(tmp00_23_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760024(.x(x_24), .z(tmp00_24_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760025(.x(x_25), .z(tmp00_25_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760026(.x(x_26), .z(tmp00_26_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760027(.x(x_27), .z(tmp00_27_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760028(.x(x_28), .z(tmp00_28_76));
	booth_0002 #(.WIDTH(WIDTH)) mul00760029(.x(x_29), .z(tmp00_29_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760030(.x(x_30), .z(tmp00_30_76));
	booth__012 #(.WIDTH(WIDTH)) mul00760031(.x(x_31), .z(tmp00_31_76));
	booth_0010 #(.WIDTH(WIDTH)) mul00760032(.x(x_32), .z(tmp00_32_76));
	booth_0010 #(.WIDTH(WIDTH)) mul00760033(.x(x_33), .z(tmp00_33_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760034(.x(x_34), .z(tmp00_34_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760035(.x(x_35), .z(tmp00_35_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760036(.x(x_36), .z(tmp00_36_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760037(.x(x_37), .z(tmp00_37_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760038(.x(x_38), .z(tmp00_38_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760039(.x(x_39), .z(tmp00_39_76));
	booth_0002 #(.WIDTH(WIDTH)) mul00760040(.x(x_40), .z(tmp00_40_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760041(.x(x_41), .z(tmp00_41_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760042(.x(x_42), .z(tmp00_42_76));
	booth_0002 #(.WIDTH(WIDTH)) mul00760043(.x(x_43), .z(tmp00_43_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760044(.x(x_44), .z(tmp00_44_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760045(.x(x_45), .z(tmp00_45_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760046(.x(x_46), .z(tmp00_46_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760047(.x(x_47), .z(tmp00_47_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760048(.x(x_48), .z(tmp00_48_76));
	booth_0012 #(.WIDTH(WIDTH)) mul00760049(.x(x_49), .z(tmp00_49_76));
	booth_0002 #(.WIDTH(WIDTH)) mul00760050(.x(x_50), .z(tmp00_50_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760051(.x(x_51), .z(tmp00_51_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760052(.x(x_52), .z(tmp00_52_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760053(.x(x_53), .z(tmp00_53_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760054(.x(x_54), .z(tmp00_54_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760055(.x(x_55), .z(tmp00_55_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760056(.x(x_56), .z(tmp00_56_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760057(.x(x_57), .z(tmp00_57_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760058(.x(x_58), .z(tmp00_58_76));
	booth_0016 #(.WIDTH(WIDTH)) mul00760059(.x(x_59), .z(tmp00_59_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760060(.x(x_60), .z(tmp00_60_76));
	booth_0006 #(.WIDTH(WIDTH)) mul00760061(.x(x_61), .z(tmp00_61_76));
	booth__006 #(.WIDTH(WIDTH)) mul00760062(.x(x_62), .z(tmp00_62_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760063(.x(x_63), .z(tmp00_63_76));
	booth__010 #(.WIDTH(WIDTH)) mul00760064(.x(x_64), .z(tmp00_64_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760065(.x(x_65), .z(tmp00_65_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760066(.x(x_66), .z(tmp00_66_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760067(.x(x_67), .z(tmp00_67_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760068(.x(x_68), .z(tmp00_68_76));
	booth__002 #(.WIDTH(WIDTH)) mul00760069(.x(x_69), .z(tmp00_69_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760070(.x(x_70), .z(tmp00_70_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760071(.x(x_71), .z(tmp00_71_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760072(.x(x_72), .z(tmp00_72_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760073(.x(x_73), .z(tmp00_73_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760074(.x(x_74), .z(tmp00_74_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760075(.x(x_75), .z(tmp00_75_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760076(.x(x_76), .z(tmp00_76_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760077(.x(x_77), .z(tmp00_77_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760078(.x(x_78), .z(tmp00_78_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760079(.x(x_79), .z(tmp00_79_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760080(.x(x_80), .z(tmp00_80_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760081(.x(x_81), .z(tmp00_81_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760082(.x(x_82), .z(tmp00_82_76));
	booth_0002 #(.WIDTH(WIDTH)) mul00760083(.x(x_83), .z(tmp00_83_76));
	booth__006 #(.WIDTH(WIDTH)) mul00760084(.x(x_84), .z(tmp00_84_76));
	booth__012 #(.WIDTH(WIDTH)) mul00760085(.x(x_85), .z(tmp00_85_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760086(.x(x_86), .z(tmp00_86_76));
	booth__002 #(.WIDTH(WIDTH)) mul00760087(.x(x_87), .z(tmp00_87_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760088(.x(x_88), .z(tmp00_88_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760089(.x(x_89), .z(tmp00_89_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760090(.x(x_90), .z(tmp00_90_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760091(.x(x_91), .z(tmp00_91_76));
	booth_0006 #(.WIDTH(WIDTH)) mul00760092(.x(x_92), .z(tmp00_92_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760093(.x(x_93), .z(tmp00_93_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760094(.x(x_94), .z(tmp00_94_76));
	booth__012 #(.WIDTH(WIDTH)) mul00760095(.x(x_95), .z(tmp00_95_76));
	booth_0010 #(.WIDTH(WIDTH)) mul00760096(.x(x_96), .z(tmp00_96_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760097(.x(x_97), .z(tmp00_97_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760098(.x(x_98), .z(tmp00_98_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760099(.x(x_99), .z(tmp00_99_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760100(.x(x_100), .z(tmp00_100_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760101(.x(x_101), .z(tmp00_101_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760102(.x(x_102), .z(tmp00_102_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760103(.x(x_103), .z(tmp00_103_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760104(.x(x_104), .z(tmp00_104_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760105(.x(x_105), .z(tmp00_105_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760106(.x(x_106), .z(tmp00_106_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760107(.x(x_107), .z(tmp00_107_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760108(.x(x_108), .z(tmp00_108_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760109(.x(x_109), .z(tmp00_109_76));
	booth__008 #(.WIDTH(WIDTH)) mul00760110(.x(x_110), .z(tmp00_110_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760111(.x(x_111), .z(tmp00_111_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760112(.x(x_112), .z(tmp00_112_76));
	booth_0008 #(.WIDTH(WIDTH)) mul00760113(.x(x_113), .z(tmp00_113_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760114(.x(x_114), .z(tmp00_114_76));
	booth_0006 #(.WIDTH(WIDTH)) mul00760115(.x(x_115), .z(tmp00_115_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760116(.x(x_116), .z(tmp00_116_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760117(.x(x_117), .z(tmp00_117_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760118(.x(x_118), .z(tmp00_118_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760119(.x(x_119), .z(tmp00_119_76));
	booth__002 #(.WIDTH(WIDTH)) mul00760120(.x(x_120), .z(tmp00_120_76));
	booth_0014 #(.WIDTH(WIDTH)) mul00760121(.x(x_121), .z(tmp00_121_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760122(.x(x_122), .z(tmp00_122_76));
	booth__004 #(.WIDTH(WIDTH)) mul00760123(.x(x_123), .z(tmp00_123_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00760124(.x(x_124), .z(tmp00_124_76));
	booth_0006 #(.WIDTH(WIDTH)) mul00760125(.x(x_125), .z(tmp00_125_76));
	booth_0002 #(.WIDTH(WIDTH)) mul00760126(.x(x_126), .z(tmp00_126_76));
	booth_0000 #(.WIDTH(WIDTH)) mul00760127(.x(x_127), .z(tmp00_127_76));
	booth_0004 #(.WIDTH(WIDTH)) mul00770000(.x(x_0), .z(tmp00_0_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770001(.x(x_1), .z(tmp00_1_77));
	booth_0002 #(.WIDTH(WIDTH)) mul00770002(.x(x_2), .z(tmp00_2_77));
	booth_0006 #(.WIDTH(WIDTH)) mul00770003(.x(x_3), .z(tmp00_3_77));
	booth_0006 #(.WIDTH(WIDTH)) mul00770004(.x(x_4), .z(tmp00_4_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770005(.x(x_5), .z(tmp00_5_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770006(.x(x_6), .z(tmp00_6_77));
	booth__004 #(.WIDTH(WIDTH)) mul00770007(.x(x_7), .z(tmp00_7_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770008(.x(x_8), .z(tmp00_8_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770009(.x(x_9), .z(tmp00_9_77));
	booth__004 #(.WIDTH(WIDTH)) mul00770010(.x(x_10), .z(tmp00_10_77));
	booth__010 #(.WIDTH(WIDTH)) mul00770011(.x(x_11), .z(tmp00_11_77));
	booth__010 #(.WIDTH(WIDTH)) mul00770012(.x(x_12), .z(tmp00_12_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770013(.x(x_13), .z(tmp00_13_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770014(.x(x_14), .z(tmp00_14_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770015(.x(x_15), .z(tmp00_15_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770016(.x(x_16), .z(tmp00_16_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770017(.x(x_17), .z(tmp00_17_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770018(.x(x_18), .z(tmp00_18_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770019(.x(x_19), .z(tmp00_19_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770020(.x(x_20), .z(tmp00_20_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770021(.x(x_21), .z(tmp00_21_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770022(.x(x_22), .z(tmp00_22_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770023(.x(x_23), .z(tmp00_23_77));
	booth_0008 #(.WIDTH(WIDTH)) mul00770024(.x(x_24), .z(tmp00_24_77));
	booth_0002 #(.WIDTH(WIDTH)) mul00770025(.x(x_25), .z(tmp00_25_77));
	booth_0010 #(.WIDTH(WIDTH)) mul00770026(.x(x_26), .z(tmp00_26_77));
	booth__006 #(.WIDTH(WIDTH)) mul00770027(.x(x_27), .z(tmp00_27_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770028(.x(x_28), .z(tmp00_28_77));
	booth_0006 #(.WIDTH(WIDTH)) mul00770029(.x(x_29), .z(tmp00_29_77));
	booth__002 #(.WIDTH(WIDTH)) mul00770030(.x(x_30), .z(tmp00_30_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770031(.x(x_31), .z(tmp00_31_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770032(.x(x_32), .z(tmp00_32_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770033(.x(x_33), .z(tmp00_33_77));
	booth__012 #(.WIDTH(WIDTH)) mul00770034(.x(x_34), .z(tmp00_34_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770035(.x(x_35), .z(tmp00_35_77));
	booth_0006 #(.WIDTH(WIDTH)) mul00770036(.x(x_36), .z(tmp00_36_77));
	booth__004 #(.WIDTH(WIDTH)) mul00770037(.x(x_37), .z(tmp00_37_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770038(.x(x_38), .z(tmp00_38_77));
	booth_0008 #(.WIDTH(WIDTH)) mul00770039(.x(x_39), .z(tmp00_39_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770040(.x(x_40), .z(tmp00_40_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770041(.x(x_41), .z(tmp00_41_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770042(.x(x_42), .z(tmp00_42_77));
	booth_0002 #(.WIDTH(WIDTH)) mul00770043(.x(x_43), .z(tmp00_43_77));
	booth_0008 #(.WIDTH(WIDTH)) mul00770044(.x(x_44), .z(tmp00_44_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770045(.x(x_45), .z(tmp00_45_77));
	booth_0016 #(.WIDTH(WIDTH)) mul00770046(.x(x_46), .z(tmp00_46_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770047(.x(x_47), .z(tmp00_47_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770048(.x(x_48), .z(tmp00_48_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770049(.x(x_49), .z(tmp00_49_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770050(.x(x_50), .z(tmp00_50_77));
	booth_0010 #(.WIDTH(WIDTH)) mul00770051(.x(x_51), .z(tmp00_51_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770052(.x(x_52), .z(tmp00_52_77));
	booth_0010 #(.WIDTH(WIDTH)) mul00770053(.x(x_53), .z(tmp00_53_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770054(.x(x_54), .z(tmp00_54_77));
	booth_0008 #(.WIDTH(WIDTH)) mul00770055(.x(x_55), .z(tmp00_55_77));
	booth_0016 #(.WIDTH(WIDTH)) mul00770056(.x(x_56), .z(tmp00_56_77));
	booth__006 #(.WIDTH(WIDTH)) mul00770057(.x(x_57), .z(tmp00_57_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770058(.x(x_58), .z(tmp00_58_77));
	booth__004 #(.WIDTH(WIDTH)) mul00770059(.x(x_59), .z(tmp00_59_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770060(.x(x_60), .z(tmp00_60_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770061(.x(x_61), .z(tmp00_61_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770062(.x(x_62), .z(tmp00_62_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770063(.x(x_63), .z(tmp00_63_77));
	booth__010 #(.WIDTH(WIDTH)) mul00770064(.x(x_64), .z(tmp00_64_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770065(.x(x_65), .z(tmp00_65_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770066(.x(x_66), .z(tmp00_66_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770067(.x(x_67), .z(tmp00_67_77));
	booth_0010 #(.WIDTH(WIDTH)) mul00770068(.x(x_68), .z(tmp00_68_77));
	booth__014 #(.WIDTH(WIDTH)) mul00770069(.x(x_69), .z(tmp00_69_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770070(.x(x_70), .z(tmp00_70_77));
	booth_0006 #(.WIDTH(WIDTH)) mul00770071(.x(x_71), .z(tmp00_71_77));
	booth__012 #(.WIDTH(WIDTH)) mul00770072(.x(x_72), .z(tmp00_72_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770073(.x(x_73), .z(tmp00_73_77));
	booth_0002 #(.WIDTH(WIDTH)) mul00770074(.x(x_74), .z(tmp00_74_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770075(.x(x_75), .z(tmp00_75_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770076(.x(x_76), .z(tmp00_76_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770077(.x(x_77), .z(tmp00_77_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770078(.x(x_78), .z(tmp00_78_77));
	booth__006 #(.WIDTH(WIDTH)) mul00770079(.x(x_79), .z(tmp00_79_77));
	booth__006 #(.WIDTH(WIDTH)) mul00770080(.x(x_80), .z(tmp00_80_77));
	booth_0008 #(.WIDTH(WIDTH)) mul00770081(.x(x_81), .z(tmp00_81_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770082(.x(x_82), .z(tmp00_82_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770083(.x(x_83), .z(tmp00_83_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770084(.x(x_84), .z(tmp00_84_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770085(.x(x_85), .z(tmp00_85_77));
	booth__004 #(.WIDTH(WIDTH)) mul00770086(.x(x_86), .z(tmp00_86_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770087(.x(x_87), .z(tmp00_87_77));
	booth__004 #(.WIDTH(WIDTH)) mul00770088(.x(x_88), .z(tmp00_88_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770089(.x(x_89), .z(tmp00_89_77));
	booth_0016 #(.WIDTH(WIDTH)) mul00770090(.x(x_90), .z(tmp00_90_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770091(.x(x_91), .z(tmp00_91_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770092(.x(x_92), .z(tmp00_92_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770093(.x(x_93), .z(tmp00_93_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770094(.x(x_94), .z(tmp00_94_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770095(.x(x_95), .z(tmp00_95_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770096(.x(x_96), .z(tmp00_96_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770097(.x(x_97), .z(tmp00_97_77));
	booth__012 #(.WIDTH(WIDTH)) mul00770098(.x(x_98), .z(tmp00_98_77));
	booth_0008 #(.WIDTH(WIDTH)) mul00770099(.x(x_99), .z(tmp00_99_77));
	booth_0010 #(.WIDTH(WIDTH)) mul00770100(.x(x_100), .z(tmp00_100_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770101(.x(x_101), .z(tmp00_101_77));
	booth__010 #(.WIDTH(WIDTH)) mul00770102(.x(x_102), .z(tmp00_102_77));
	booth_0002 #(.WIDTH(WIDTH)) mul00770103(.x(x_103), .z(tmp00_103_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770104(.x(x_104), .z(tmp00_104_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770105(.x(x_105), .z(tmp00_105_77));
	booth_0008 #(.WIDTH(WIDTH)) mul00770106(.x(x_106), .z(tmp00_106_77));
	booth__006 #(.WIDTH(WIDTH)) mul00770107(.x(x_107), .z(tmp00_107_77));
	booth_0010 #(.WIDTH(WIDTH)) mul00770108(.x(x_108), .z(tmp00_108_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770109(.x(x_109), .z(tmp00_109_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770110(.x(x_110), .z(tmp00_110_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770111(.x(x_111), .z(tmp00_111_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770112(.x(x_112), .z(tmp00_112_77));
	booth__002 #(.WIDTH(WIDTH)) mul00770113(.x(x_113), .z(tmp00_113_77));
	booth_0006 #(.WIDTH(WIDTH)) mul00770114(.x(x_114), .z(tmp00_114_77));
	booth__006 #(.WIDTH(WIDTH)) mul00770115(.x(x_115), .z(tmp00_115_77));
	booth_0002 #(.WIDTH(WIDTH)) mul00770116(.x(x_116), .z(tmp00_116_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770117(.x(x_117), .z(tmp00_117_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770118(.x(x_118), .z(tmp00_118_77));
	booth_0012 #(.WIDTH(WIDTH)) mul00770119(.x(x_119), .z(tmp00_119_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770120(.x(x_120), .z(tmp00_120_77));
	booth__016 #(.WIDTH(WIDTH)) mul00770121(.x(x_121), .z(tmp00_121_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770122(.x(x_122), .z(tmp00_122_77));
	booth__008 #(.WIDTH(WIDTH)) mul00770123(.x(x_123), .z(tmp00_123_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770124(.x(x_124), .z(tmp00_124_77));
	booth__004 #(.WIDTH(WIDTH)) mul00770125(.x(x_125), .z(tmp00_125_77));
	booth_0000 #(.WIDTH(WIDTH)) mul00770126(.x(x_126), .z(tmp00_126_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00770127(.x(x_127), .z(tmp00_127_77));
	booth_0004 #(.WIDTH(WIDTH)) mul00780000(.x(x_0), .z(tmp00_0_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780001(.x(x_1), .z(tmp00_1_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780002(.x(x_2), .z(tmp00_2_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780003(.x(x_3), .z(tmp00_3_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780004(.x(x_4), .z(tmp00_4_78));
	booth_0010 #(.WIDTH(WIDTH)) mul00780005(.x(x_5), .z(tmp00_5_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780006(.x(x_6), .z(tmp00_6_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780007(.x(x_7), .z(tmp00_7_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780008(.x(x_8), .z(tmp00_8_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780009(.x(x_9), .z(tmp00_9_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780010(.x(x_10), .z(tmp00_10_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780011(.x(x_11), .z(tmp00_11_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780012(.x(x_12), .z(tmp00_12_78));
	booth_0010 #(.WIDTH(WIDTH)) mul00780013(.x(x_13), .z(tmp00_13_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780014(.x(x_14), .z(tmp00_14_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780015(.x(x_15), .z(tmp00_15_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780016(.x(x_16), .z(tmp00_16_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780017(.x(x_17), .z(tmp00_17_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780018(.x(x_18), .z(tmp00_18_78));
	booth_0012 #(.WIDTH(WIDTH)) mul00780019(.x(x_19), .z(tmp00_19_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780020(.x(x_20), .z(tmp00_20_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780021(.x(x_21), .z(tmp00_21_78));
	booth_0002 #(.WIDTH(WIDTH)) mul00780022(.x(x_22), .z(tmp00_22_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780023(.x(x_23), .z(tmp00_23_78));
	booth_0012 #(.WIDTH(WIDTH)) mul00780024(.x(x_24), .z(tmp00_24_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780025(.x(x_25), .z(tmp00_25_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780026(.x(x_26), .z(tmp00_26_78));
	booth_0010 #(.WIDTH(WIDTH)) mul00780027(.x(x_27), .z(tmp00_27_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780028(.x(x_28), .z(tmp00_28_78));
	booth_0006 #(.WIDTH(WIDTH)) mul00780029(.x(x_29), .z(tmp00_29_78));
	booth__006 #(.WIDTH(WIDTH)) mul00780030(.x(x_30), .z(tmp00_30_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780031(.x(x_31), .z(tmp00_31_78));
	booth_0012 #(.WIDTH(WIDTH)) mul00780032(.x(x_32), .z(tmp00_32_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780033(.x(x_33), .z(tmp00_33_78));
	booth__010 #(.WIDTH(WIDTH)) mul00780034(.x(x_34), .z(tmp00_34_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780035(.x(x_35), .z(tmp00_35_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780036(.x(x_36), .z(tmp00_36_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780037(.x(x_37), .z(tmp00_37_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780038(.x(x_38), .z(tmp00_38_78));
	booth_0018 #(.WIDTH(WIDTH)) mul00780039(.x(x_39), .z(tmp00_39_78));
	booth_0012 #(.WIDTH(WIDTH)) mul00780040(.x(x_40), .z(tmp00_40_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780041(.x(x_41), .z(tmp00_41_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780042(.x(x_42), .z(tmp00_42_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780043(.x(x_43), .z(tmp00_43_78));
	booth__016 #(.WIDTH(WIDTH)) mul00780044(.x(x_44), .z(tmp00_44_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780045(.x(x_45), .z(tmp00_45_78));
	booth_0012 #(.WIDTH(WIDTH)) mul00780046(.x(x_46), .z(tmp00_46_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780047(.x(x_47), .z(tmp00_47_78));
	booth_0010 #(.WIDTH(WIDTH)) mul00780048(.x(x_48), .z(tmp00_48_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780049(.x(x_49), .z(tmp00_49_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780050(.x(x_50), .z(tmp00_50_78));
	booth_0010 #(.WIDTH(WIDTH)) mul00780051(.x(x_51), .z(tmp00_51_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780052(.x(x_52), .z(tmp00_52_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780053(.x(x_53), .z(tmp00_53_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780054(.x(x_54), .z(tmp00_54_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780055(.x(x_55), .z(tmp00_55_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780056(.x(x_56), .z(tmp00_56_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780057(.x(x_57), .z(tmp00_57_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780058(.x(x_58), .z(tmp00_58_78));
	booth_0016 #(.WIDTH(WIDTH)) mul00780059(.x(x_59), .z(tmp00_59_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780060(.x(x_60), .z(tmp00_60_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780061(.x(x_61), .z(tmp00_61_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780062(.x(x_62), .z(tmp00_62_78));
	booth_0002 #(.WIDTH(WIDTH)) mul00780063(.x(x_63), .z(tmp00_63_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780064(.x(x_64), .z(tmp00_64_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780065(.x(x_65), .z(tmp00_65_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780066(.x(x_66), .z(tmp00_66_78));
	booth__010 #(.WIDTH(WIDTH)) mul00780067(.x(x_67), .z(tmp00_67_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780068(.x(x_68), .z(tmp00_68_78));
	booth_0010 #(.WIDTH(WIDTH)) mul00780069(.x(x_69), .z(tmp00_69_78));
	booth__010 #(.WIDTH(WIDTH)) mul00780070(.x(x_70), .z(tmp00_70_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780071(.x(x_71), .z(tmp00_71_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780072(.x(x_72), .z(tmp00_72_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780073(.x(x_73), .z(tmp00_73_78));
	booth__010 #(.WIDTH(WIDTH)) mul00780074(.x(x_74), .z(tmp00_74_78));
	booth_0002 #(.WIDTH(WIDTH)) mul00780075(.x(x_75), .z(tmp00_75_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780076(.x(x_76), .z(tmp00_76_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780077(.x(x_77), .z(tmp00_77_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780078(.x(x_78), .z(tmp00_78_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780079(.x(x_79), .z(tmp00_79_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780080(.x(x_80), .z(tmp00_80_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780081(.x(x_81), .z(tmp00_81_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780082(.x(x_82), .z(tmp00_82_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780083(.x(x_83), .z(tmp00_83_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780084(.x(x_84), .z(tmp00_84_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780085(.x(x_85), .z(tmp00_85_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780086(.x(x_86), .z(tmp00_86_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780087(.x(x_87), .z(tmp00_87_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780088(.x(x_88), .z(tmp00_88_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780089(.x(x_89), .z(tmp00_89_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780090(.x(x_90), .z(tmp00_90_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780091(.x(x_91), .z(tmp00_91_78));
	booth__012 #(.WIDTH(WIDTH)) mul00780092(.x(x_92), .z(tmp00_92_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780093(.x(x_93), .z(tmp00_93_78));
	booth_0012 #(.WIDTH(WIDTH)) mul00780094(.x(x_94), .z(tmp00_94_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780095(.x(x_95), .z(tmp00_95_78));
	booth_0016 #(.WIDTH(WIDTH)) mul00780096(.x(x_96), .z(tmp00_96_78));
	booth_0006 #(.WIDTH(WIDTH)) mul00780097(.x(x_97), .z(tmp00_97_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780098(.x(x_98), .z(tmp00_98_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780099(.x(x_99), .z(tmp00_99_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780100(.x(x_100), .z(tmp00_100_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780101(.x(x_101), .z(tmp00_101_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780102(.x(x_102), .z(tmp00_102_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780103(.x(x_103), .z(tmp00_103_78));
	booth__002 #(.WIDTH(WIDTH)) mul00780104(.x(x_104), .z(tmp00_104_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780105(.x(x_105), .z(tmp00_105_78));
	booth_0002 #(.WIDTH(WIDTH)) mul00780106(.x(x_106), .z(tmp00_106_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780107(.x(x_107), .z(tmp00_107_78));
	booth__012 #(.WIDTH(WIDTH)) mul00780108(.x(x_108), .z(tmp00_108_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780109(.x(x_109), .z(tmp00_109_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780110(.x(x_110), .z(tmp00_110_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780111(.x(x_111), .z(tmp00_111_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780112(.x(x_112), .z(tmp00_112_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780113(.x(x_113), .z(tmp00_113_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780114(.x(x_114), .z(tmp00_114_78));
	booth__008 #(.WIDTH(WIDTH)) mul00780115(.x(x_115), .z(tmp00_115_78));
	booth_0012 #(.WIDTH(WIDTH)) mul00780116(.x(x_116), .z(tmp00_116_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780117(.x(x_117), .z(tmp00_117_78));
	booth__004 #(.WIDTH(WIDTH)) mul00780118(.x(x_118), .z(tmp00_118_78));
	booth__016 #(.WIDTH(WIDTH)) mul00780119(.x(x_119), .z(tmp00_119_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780120(.x(x_120), .z(tmp00_120_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780121(.x(x_121), .z(tmp00_121_78));
	booth_0002 #(.WIDTH(WIDTH)) mul00780122(.x(x_122), .z(tmp00_122_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780123(.x(x_123), .z(tmp00_123_78));
	booth_0016 #(.WIDTH(WIDTH)) mul00780124(.x(x_124), .z(tmp00_124_78));
	booth_0008 #(.WIDTH(WIDTH)) mul00780125(.x(x_125), .z(tmp00_125_78));
	booth_0004 #(.WIDTH(WIDTH)) mul00780126(.x(x_126), .z(tmp00_126_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00780127(.x(x_127), .z(tmp00_127_78));
	booth_0000 #(.WIDTH(WIDTH)) mul00790000(.x(x_0), .z(tmp00_0_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790001(.x(x_1), .z(tmp00_1_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790002(.x(x_2), .z(tmp00_2_79));
	booth_0010 #(.WIDTH(WIDTH)) mul00790003(.x(x_3), .z(tmp00_3_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790004(.x(x_4), .z(tmp00_4_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790005(.x(x_5), .z(tmp00_5_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790006(.x(x_6), .z(tmp00_6_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790007(.x(x_7), .z(tmp00_7_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790008(.x(x_8), .z(tmp00_8_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790009(.x(x_9), .z(tmp00_9_79));
	booth_0002 #(.WIDTH(WIDTH)) mul00790010(.x(x_10), .z(tmp00_10_79));
	booth_0010 #(.WIDTH(WIDTH)) mul00790011(.x(x_11), .z(tmp00_11_79));
	booth_0002 #(.WIDTH(WIDTH)) mul00790012(.x(x_12), .z(tmp00_12_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790013(.x(x_13), .z(tmp00_13_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790014(.x(x_14), .z(tmp00_14_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790015(.x(x_15), .z(tmp00_15_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790016(.x(x_16), .z(tmp00_16_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790017(.x(x_17), .z(tmp00_17_79));
	booth__006 #(.WIDTH(WIDTH)) mul00790018(.x(x_18), .z(tmp00_18_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790019(.x(x_19), .z(tmp00_19_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790020(.x(x_20), .z(tmp00_20_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790021(.x(x_21), .z(tmp00_21_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790022(.x(x_22), .z(tmp00_22_79));
	booth_0006 #(.WIDTH(WIDTH)) mul00790023(.x(x_23), .z(tmp00_23_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790024(.x(x_24), .z(tmp00_24_79));
	booth_0006 #(.WIDTH(WIDTH)) mul00790025(.x(x_25), .z(tmp00_25_79));
	booth__006 #(.WIDTH(WIDTH)) mul00790026(.x(x_26), .z(tmp00_26_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790027(.x(x_27), .z(tmp00_27_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790028(.x(x_28), .z(tmp00_28_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790029(.x(x_29), .z(tmp00_29_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790030(.x(x_30), .z(tmp00_30_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790031(.x(x_31), .z(tmp00_31_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790032(.x(x_32), .z(tmp00_32_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790033(.x(x_33), .z(tmp00_33_79));
	booth_0010 #(.WIDTH(WIDTH)) mul00790034(.x(x_34), .z(tmp00_34_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790035(.x(x_35), .z(tmp00_35_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790036(.x(x_36), .z(tmp00_36_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790037(.x(x_37), .z(tmp00_37_79));
	booth_0002 #(.WIDTH(WIDTH)) mul00790038(.x(x_38), .z(tmp00_38_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790039(.x(x_39), .z(tmp00_39_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790040(.x(x_40), .z(tmp00_40_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790041(.x(x_41), .z(tmp00_41_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790042(.x(x_42), .z(tmp00_42_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790043(.x(x_43), .z(tmp00_43_79));
	booth__010 #(.WIDTH(WIDTH)) mul00790044(.x(x_44), .z(tmp00_44_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790045(.x(x_45), .z(tmp00_45_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790046(.x(x_46), .z(tmp00_46_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790047(.x(x_47), .z(tmp00_47_79));
	booth_0010 #(.WIDTH(WIDTH)) mul00790048(.x(x_48), .z(tmp00_48_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790049(.x(x_49), .z(tmp00_49_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790050(.x(x_50), .z(tmp00_50_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790051(.x(x_51), .z(tmp00_51_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790052(.x(x_52), .z(tmp00_52_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790053(.x(x_53), .z(tmp00_53_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790054(.x(x_54), .z(tmp00_54_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790055(.x(x_55), .z(tmp00_55_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790056(.x(x_56), .z(tmp00_56_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790057(.x(x_57), .z(tmp00_57_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790058(.x(x_58), .z(tmp00_58_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790059(.x(x_59), .z(tmp00_59_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790060(.x(x_60), .z(tmp00_60_79));
	booth__010 #(.WIDTH(WIDTH)) mul00790061(.x(x_61), .z(tmp00_61_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790062(.x(x_62), .z(tmp00_62_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790063(.x(x_63), .z(tmp00_63_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790064(.x(x_64), .z(tmp00_64_79));
	booth__006 #(.WIDTH(WIDTH)) mul00790065(.x(x_65), .z(tmp00_65_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790066(.x(x_66), .z(tmp00_66_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790067(.x(x_67), .z(tmp00_67_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790068(.x(x_68), .z(tmp00_68_79));
	booth__006 #(.WIDTH(WIDTH)) mul00790069(.x(x_69), .z(tmp00_69_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790070(.x(x_70), .z(tmp00_70_79));
	booth_0010 #(.WIDTH(WIDTH)) mul00790071(.x(x_71), .z(tmp00_71_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790072(.x(x_72), .z(tmp00_72_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790073(.x(x_73), .z(tmp00_73_79));
	booth__006 #(.WIDTH(WIDTH)) mul00790074(.x(x_74), .z(tmp00_74_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790075(.x(x_75), .z(tmp00_75_79));
	booth__012 #(.WIDTH(WIDTH)) mul00790076(.x(x_76), .z(tmp00_76_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790077(.x(x_77), .z(tmp00_77_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790078(.x(x_78), .z(tmp00_78_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790079(.x(x_79), .z(tmp00_79_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790080(.x(x_80), .z(tmp00_80_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790081(.x(x_81), .z(tmp00_81_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790082(.x(x_82), .z(tmp00_82_79));
	booth_0006 #(.WIDTH(WIDTH)) mul00790083(.x(x_83), .z(tmp00_83_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790084(.x(x_84), .z(tmp00_84_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790085(.x(x_85), .z(tmp00_85_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790086(.x(x_86), .z(tmp00_86_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790087(.x(x_87), .z(tmp00_87_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790088(.x(x_88), .z(tmp00_88_79));
	booth__006 #(.WIDTH(WIDTH)) mul00790089(.x(x_89), .z(tmp00_89_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790090(.x(x_90), .z(tmp00_90_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790091(.x(x_91), .z(tmp00_91_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790092(.x(x_92), .z(tmp00_92_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790093(.x(x_93), .z(tmp00_93_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790094(.x(x_94), .z(tmp00_94_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790095(.x(x_95), .z(tmp00_95_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790096(.x(x_96), .z(tmp00_96_79));
	booth__010 #(.WIDTH(WIDTH)) mul00790097(.x(x_97), .z(tmp00_97_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790098(.x(x_98), .z(tmp00_98_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790099(.x(x_99), .z(tmp00_99_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790100(.x(x_100), .z(tmp00_100_79));
	booth__002 #(.WIDTH(WIDTH)) mul00790101(.x(x_101), .z(tmp00_101_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790102(.x(x_102), .z(tmp00_102_79));
	booth__006 #(.WIDTH(WIDTH)) mul00790103(.x(x_103), .z(tmp00_103_79));
	booth_0010 #(.WIDTH(WIDTH)) mul00790104(.x(x_104), .z(tmp00_104_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790105(.x(x_105), .z(tmp00_105_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790106(.x(x_106), .z(tmp00_106_79));
	booth_0006 #(.WIDTH(WIDTH)) mul00790107(.x(x_107), .z(tmp00_107_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790108(.x(x_108), .z(tmp00_108_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790109(.x(x_109), .z(tmp00_109_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790110(.x(x_110), .z(tmp00_110_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790111(.x(x_111), .z(tmp00_111_79));
	booth_0006 #(.WIDTH(WIDTH)) mul00790112(.x(x_112), .z(tmp00_112_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790113(.x(x_113), .z(tmp00_113_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790114(.x(x_114), .z(tmp00_114_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790115(.x(x_115), .z(tmp00_115_79));
	booth_0006 #(.WIDTH(WIDTH)) mul00790116(.x(x_116), .z(tmp00_116_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790117(.x(x_117), .z(tmp00_117_79));
	booth_0008 #(.WIDTH(WIDTH)) mul00790118(.x(x_118), .z(tmp00_118_79));
	booth_0000 #(.WIDTH(WIDTH)) mul00790119(.x(x_119), .z(tmp00_119_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790120(.x(x_120), .z(tmp00_120_79));
	booth_0006 #(.WIDTH(WIDTH)) mul00790121(.x(x_121), .z(tmp00_121_79));
	booth__004 #(.WIDTH(WIDTH)) mul00790122(.x(x_122), .z(tmp00_122_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790123(.x(x_123), .z(tmp00_123_79));
	booth__008 #(.WIDTH(WIDTH)) mul00790124(.x(x_124), .z(tmp00_124_79));
	booth_0010 #(.WIDTH(WIDTH)) mul00790125(.x(x_125), .z(tmp00_125_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790126(.x(x_126), .z(tmp00_126_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00790127(.x(x_127), .z(tmp00_127_79));
	booth_0004 #(.WIDTH(WIDTH)) mul00800000(.x(x_0), .z(tmp00_0_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800001(.x(x_1), .z(tmp00_1_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800002(.x(x_2), .z(tmp00_2_80));
	booth__008 #(.WIDTH(WIDTH)) mul00800003(.x(x_3), .z(tmp00_3_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800004(.x(x_4), .z(tmp00_4_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800005(.x(x_5), .z(tmp00_5_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800006(.x(x_6), .z(tmp00_6_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800007(.x(x_7), .z(tmp00_7_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800008(.x(x_8), .z(tmp00_8_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800009(.x(x_9), .z(tmp00_9_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800010(.x(x_10), .z(tmp00_10_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800011(.x(x_11), .z(tmp00_11_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800012(.x(x_12), .z(tmp00_12_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800013(.x(x_13), .z(tmp00_13_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800014(.x(x_14), .z(tmp00_14_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800015(.x(x_15), .z(tmp00_15_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800016(.x(x_16), .z(tmp00_16_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800017(.x(x_17), .z(tmp00_17_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800018(.x(x_18), .z(tmp00_18_80));
	booth_0010 #(.WIDTH(WIDTH)) mul00800019(.x(x_19), .z(tmp00_19_80));
	booth_0012 #(.WIDTH(WIDTH)) mul00800020(.x(x_20), .z(tmp00_20_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800021(.x(x_21), .z(tmp00_21_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800022(.x(x_22), .z(tmp00_22_80));
	booth__008 #(.WIDTH(WIDTH)) mul00800023(.x(x_23), .z(tmp00_23_80));
	booth_0006 #(.WIDTH(WIDTH)) mul00800024(.x(x_24), .z(tmp00_24_80));
	booth__002 #(.WIDTH(WIDTH)) mul00800025(.x(x_25), .z(tmp00_25_80));
	booth_0010 #(.WIDTH(WIDTH)) mul00800026(.x(x_26), .z(tmp00_26_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800027(.x(x_27), .z(tmp00_27_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800028(.x(x_28), .z(tmp00_28_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800029(.x(x_29), .z(tmp00_29_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800030(.x(x_30), .z(tmp00_30_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800031(.x(x_31), .z(tmp00_31_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800032(.x(x_32), .z(tmp00_32_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800033(.x(x_33), .z(tmp00_33_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800034(.x(x_34), .z(tmp00_34_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800035(.x(x_35), .z(tmp00_35_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800036(.x(x_36), .z(tmp00_36_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800037(.x(x_37), .z(tmp00_37_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800038(.x(x_38), .z(tmp00_38_80));
	booth__008 #(.WIDTH(WIDTH)) mul00800039(.x(x_39), .z(tmp00_39_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800040(.x(x_40), .z(tmp00_40_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800041(.x(x_41), .z(tmp00_41_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800042(.x(x_42), .z(tmp00_42_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800043(.x(x_43), .z(tmp00_43_80));
	booth__008 #(.WIDTH(WIDTH)) mul00800044(.x(x_44), .z(tmp00_44_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800045(.x(x_45), .z(tmp00_45_80));
	booth__008 #(.WIDTH(WIDTH)) mul00800046(.x(x_46), .z(tmp00_46_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800047(.x(x_47), .z(tmp00_47_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800048(.x(x_48), .z(tmp00_48_80));
	booth__008 #(.WIDTH(WIDTH)) mul00800049(.x(x_49), .z(tmp00_49_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800050(.x(x_50), .z(tmp00_50_80));
	booth__002 #(.WIDTH(WIDTH)) mul00800051(.x(x_51), .z(tmp00_51_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800052(.x(x_52), .z(tmp00_52_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800053(.x(x_53), .z(tmp00_53_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800054(.x(x_54), .z(tmp00_54_80));
	booth_0012 #(.WIDTH(WIDTH)) mul00800055(.x(x_55), .z(tmp00_55_80));
	booth_0010 #(.WIDTH(WIDTH)) mul00800056(.x(x_56), .z(tmp00_56_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800057(.x(x_57), .z(tmp00_57_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800058(.x(x_58), .z(tmp00_58_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800059(.x(x_59), .z(tmp00_59_80));
	booth_0006 #(.WIDTH(WIDTH)) mul00800060(.x(x_60), .z(tmp00_60_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800061(.x(x_61), .z(tmp00_61_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800062(.x(x_62), .z(tmp00_62_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800063(.x(x_63), .z(tmp00_63_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800064(.x(x_64), .z(tmp00_64_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800065(.x(x_65), .z(tmp00_65_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800066(.x(x_66), .z(tmp00_66_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800067(.x(x_67), .z(tmp00_67_80));
	booth_0012 #(.WIDTH(WIDTH)) mul00800068(.x(x_68), .z(tmp00_68_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800069(.x(x_69), .z(tmp00_69_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800070(.x(x_70), .z(tmp00_70_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800071(.x(x_71), .z(tmp00_71_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800072(.x(x_72), .z(tmp00_72_80));
	booth__008 #(.WIDTH(WIDTH)) mul00800073(.x(x_73), .z(tmp00_73_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800074(.x(x_74), .z(tmp00_74_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800075(.x(x_75), .z(tmp00_75_80));
	booth__012 #(.WIDTH(WIDTH)) mul00800076(.x(x_76), .z(tmp00_76_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800077(.x(x_77), .z(tmp00_77_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800078(.x(x_78), .z(tmp00_78_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800079(.x(x_79), .z(tmp00_79_80));
	booth_0006 #(.WIDTH(WIDTH)) mul00800080(.x(x_80), .z(tmp00_80_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800081(.x(x_81), .z(tmp00_81_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800082(.x(x_82), .z(tmp00_82_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800083(.x(x_83), .z(tmp00_83_80));
	booth__010 #(.WIDTH(WIDTH)) mul00800084(.x(x_84), .z(tmp00_84_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800085(.x(x_85), .z(tmp00_85_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800086(.x(x_86), .z(tmp00_86_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800087(.x(x_87), .z(tmp00_87_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800088(.x(x_88), .z(tmp00_88_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800089(.x(x_89), .z(tmp00_89_80));
	booth_0012 #(.WIDTH(WIDTH)) mul00800090(.x(x_90), .z(tmp00_90_80));
	booth_0012 #(.WIDTH(WIDTH)) mul00800091(.x(x_91), .z(tmp00_91_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800092(.x(x_92), .z(tmp00_92_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800093(.x(x_93), .z(tmp00_93_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800094(.x(x_94), .z(tmp00_94_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800095(.x(x_95), .z(tmp00_95_80));
	booth__012 #(.WIDTH(WIDTH)) mul00800096(.x(x_96), .z(tmp00_96_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800097(.x(x_97), .z(tmp00_97_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800098(.x(x_98), .z(tmp00_98_80));
	booth__002 #(.WIDTH(WIDTH)) mul00800099(.x(x_99), .z(tmp00_99_80));
	booth__002 #(.WIDTH(WIDTH)) mul00800100(.x(x_100), .z(tmp00_100_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800101(.x(x_101), .z(tmp00_101_80));
	booth_0002 #(.WIDTH(WIDTH)) mul00800102(.x(x_102), .z(tmp00_102_80));
	booth__010 #(.WIDTH(WIDTH)) mul00800103(.x(x_103), .z(tmp00_103_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800104(.x(x_104), .z(tmp00_104_80));
	booth__006 #(.WIDTH(WIDTH)) mul00800105(.x(x_105), .z(tmp00_105_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800106(.x(x_106), .z(tmp00_106_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800107(.x(x_107), .z(tmp00_107_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800108(.x(x_108), .z(tmp00_108_80));
	booth__010 #(.WIDTH(WIDTH)) mul00800109(.x(x_109), .z(tmp00_109_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800110(.x(x_110), .z(tmp00_110_80));
	booth__002 #(.WIDTH(WIDTH)) mul00800111(.x(x_111), .z(tmp00_111_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800112(.x(x_112), .z(tmp00_112_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800113(.x(x_113), .z(tmp00_113_80));
	booth__010 #(.WIDTH(WIDTH)) mul00800114(.x(x_114), .z(tmp00_114_80));
	booth_0014 #(.WIDTH(WIDTH)) mul00800115(.x(x_115), .z(tmp00_115_80));
	booth_0006 #(.WIDTH(WIDTH)) mul00800116(.x(x_116), .z(tmp00_116_80));
	booth__002 #(.WIDTH(WIDTH)) mul00800117(.x(x_117), .z(tmp00_117_80));
	booth_0004 #(.WIDTH(WIDTH)) mul00800118(.x(x_118), .z(tmp00_118_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800119(.x(x_119), .z(tmp00_119_80));
	booth_0000 #(.WIDTH(WIDTH)) mul00800120(.x(x_120), .z(tmp00_120_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800121(.x(x_121), .z(tmp00_121_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800122(.x(x_122), .z(tmp00_122_80));
	booth__004 #(.WIDTH(WIDTH)) mul00800123(.x(x_123), .z(tmp00_123_80));
	booth__012 #(.WIDTH(WIDTH)) mul00800124(.x(x_124), .z(tmp00_124_80));
	booth_0006 #(.WIDTH(WIDTH)) mul00800125(.x(x_125), .z(tmp00_125_80));
	booth_0010 #(.WIDTH(WIDTH)) mul00800126(.x(x_126), .z(tmp00_126_80));
	booth_0008 #(.WIDTH(WIDTH)) mul00800127(.x(x_127), .z(tmp00_127_80));
	booth__004 #(.WIDTH(WIDTH)) mul00810000(.x(x_0), .z(tmp00_0_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810001(.x(x_1), .z(tmp00_1_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810002(.x(x_2), .z(tmp00_2_81));
	booth__002 #(.WIDTH(WIDTH)) mul00810003(.x(x_3), .z(tmp00_3_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810004(.x(x_4), .z(tmp00_4_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810005(.x(x_5), .z(tmp00_5_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810006(.x(x_6), .z(tmp00_6_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810007(.x(x_7), .z(tmp00_7_81));
	booth__010 #(.WIDTH(WIDTH)) mul00810008(.x(x_8), .z(tmp00_8_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810009(.x(x_9), .z(tmp00_9_81));
	booth__006 #(.WIDTH(WIDTH)) mul00810010(.x(x_10), .z(tmp00_10_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810011(.x(x_11), .z(tmp00_11_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810012(.x(x_12), .z(tmp00_12_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810013(.x(x_13), .z(tmp00_13_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810014(.x(x_14), .z(tmp00_14_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810015(.x(x_15), .z(tmp00_15_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810016(.x(x_16), .z(tmp00_16_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810017(.x(x_17), .z(tmp00_17_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810018(.x(x_18), .z(tmp00_18_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810019(.x(x_19), .z(tmp00_19_81));
	booth_0002 #(.WIDTH(WIDTH)) mul00810020(.x(x_20), .z(tmp00_20_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810021(.x(x_21), .z(tmp00_21_81));
	booth__010 #(.WIDTH(WIDTH)) mul00810022(.x(x_22), .z(tmp00_22_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810023(.x(x_23), .z(tmp00_23_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810024(.x(x_24), .z(tmp00_24_81));
	booth_0002 #(.WIDTH(WIDTH)) mul00810025(.x(x_25), .z(tmp00_25_81));
	booth__006 #(.WIDTH(WIDTH)) mul00810026(.x(x_26), .z(tmp00_26_81));
	booth__002 #(.WIDTH(WIDTH)) mul00810027(.x(x_27), .z(tmp00_27_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810028(.x(x_28), .z(tmp00_28_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810029(.x(x_29), .z(tmp00_29_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810030(.x(x_30), .z(tmp00_30_81));
	booth__006 #(.WIDTH(WIDTH)) mul00810031(.x(x_31), .z(tmp00_31_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810032(.x(x_32), .z(tmp00_32_81));
	booth_0006 #(.WIDTH(WIDTH)) mul00810033(.x(x_33), .z(tmp00_33_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810034(.x(x_34), .z(tmp00_34_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810035(.x(x_35), .z(tmp00_35_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810036(.x(x_36), .z(tmp00_36_81));
	booth__006 #(.WIDTH(WIDTH)) mul00810037(.x(x_37), .z(tmp00_37_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810038(.x(x_38), .z(tmp00_38_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810039(.x(x_39), .z(tmp00_39_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810040(.x(x_40), .z(tmp00_40_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810041(.x(x_41), .z(tmp00_41_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810042(.x(x_42), .z(tmp00_42_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810043(.x(x_43), .z(tmp00_43_81));
	booth__010 #(.WIDTH(WIDTH)) mul00810044(.x(x_44), .z(tmp00_44_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810045(.x(x_45), .z(tmp00_45_81));
	booth__010 #(.WIDTH(WIDTH)) mul00810046(.x(x_46), .z(tmp00_46_81));
	booth__006 #(.WIDTH(WIDTH)) mul00810047(.x(x_47), .z(tmp00_47_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810048(.x(x_48), .z(tmp00_48_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810049(.x(x_49), .z(tmp00_49_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810050(.x(x_50), .z(tmp00_50_81));
	booth__010 #(.WIDTH(WIDTH)) mul00810051(.x(x_51), .z(tmp00_51_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810052(.x(x_52), .z(tmp00_52_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810053(.x(x_53), .z(tmp00_53_81));
	booth__002 #(.WIDTH(WIDTH)) mul00810054(.x(x_54), .z(tmp00_54_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810055(.x(x_55), .z(tmp00_55_81));
	booth__002 #(.WIDTH(WIDTH)) mul00810056(.x(x_56), .z(tmp00_56_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810057(.x(x_57), .z(tmp00_57_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810058(.x(x_58), .z(tmp00_58_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810059(.x(x_59), .z(tmp00_59_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810060(.x(x_60), .z(tmp00_60_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810061(.x(x_61), .z(tmp00_61_81));
	booth_0012 #(.WIDTH(WIDTH)) mul00810062(.x(x_62), .z(tmp00_62_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810063(.x(x_63), .z(tmp00_63_81));
	booth__002 #(.WIDTH(WIDTH)) mul00810064(.x(x_64), .z(tmp00_64_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810065(.x(x_65), .z(tmp00_65_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810066(.x(x_66), .z(tmp00_66_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810067(.x(x_67), .z(tmp00_67_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810068(.x(x_68), .z(tmp00_68_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810069(.x(x_69), .z(tmp00_69_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810070(.x(x_70), .z(tmp00_70_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810071(.x(x_71), .z(tmp00_71_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810072(.x(x_72), .z(tmp00_72_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810073(.x(x_73), .z(tmp00_73_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810074(.x(x_74), .z(tmp00_74_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810075(.x(x_75), .z(tmp00_75_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810076(.x(x_76), .z(tmp00_76_81));
	booth_0010 #(.WIDTH(WIDTH)) mul00810077(.x(x_77), .z(tmp00_77_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810078(.x(x_78), .z(tmp00_78_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810079(.x(x_79), .z(tmp00_79_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810080(.x(x_80), .z(tmp00_80_81));
	booth_0006 #(.WIDTH(WIDTH)) mul00810081(.x(x_81), .z(tmp00_81_81));
	booth_0006 #(.WIDTH(WIDTH)) mul00810082(.x(x_82), .z(tmp00_82_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810083(.x(x_83), .z(tmp00_83_81));
	booth__002 #(.WIDTH(WIDTH)) mul00810084(.x(x_84), .z(tmp00_84_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810085(.x(x_85), .z(tmp00_85_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810086(.x(x_86), .z(tmp00_86_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810087(.x(x_87), .z(tmp00_87_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810088(.x(x_88), .z(tmp00_88_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810089(.x(x_89), .z(tmp00_89_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810090(.x(x_90), .z(tmp00_90_81));
	booth_0006 #(.WIDTH(WIDTH)) mul00810091(.x(x_91), .z(tmp00_91_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810092(.x(x_92), .z(tmp00_92_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810093(.x(x_93), .z(tmp00_93_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810094(.x(x_94), .z(tmp00_94_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810095(.x(x_95), .z(tmp00_95_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810096(.x(x_96), .z(tmp00_96_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810097(.x(x_97), .z(tmp00_97_81));
	booth__006 #(.WIDTH(WIDTH)) mul00810098(.x(x_98), .z(tmp00_98_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810099(.x(x_99), .z(tmp00_99_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810100(.x(x_100), .z(tmp00_100_81));
	booth__012 #(.WIDTH(WIDTH)) mul00810101(.x(x_101), .z(tmp00_101_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810102(.x(x_102), .z(tmp00_102_81));
	booth_0010 #(.WIDTH(WIDTH)) mul00810103(.x(x_103), .z(tmp00_103_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810104(.x(x_104), .z(tmp00_104_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810105(.x(x_105), .z(tmp00_105_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810106(.x(x_106), .z(tmp00_106_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810107(.x(x_107), .z(tmp00_107_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810108(.x(x_108), .z(tmp00_108_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810109(.x(x_109), .z(tmp00_109_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810110(.x(x_110), .z(tmp00_110_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810111(.x(x_111), .z(tmp00_111_81));
	booth__006 #(.WIDTH(WIDTH)) mul00810112(.x(x_112), .z(tmp00_112_81));
	booth_0002 #(.WIDTH(WIDTH)) mul00810113(.x(x_113), .z(tmp00_113_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810114(.x(x_114), .z(tmp00_114_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810115(.x(x_115), .z(tmp00_115_81));
	booth__006 #(.WIDTH(WIDTH)) mul00810116(.x(x_116), .z(tmp00_116_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810117(.x(x_117), .z(tmp00_117_81));
	booth_0002 #(.WIDTH(WIDTH)) mul00810118(.x(x_118), .z(tmp00_118_81));
	booth_0002 #(.WIDTH(WIDTH)) mul00810119(.x(x_119), .z(tmp00_119_81));
	booth__008 #(.WIDTH(WIDTH)) mul00810120(.x(x_120), .z(tmp00_120_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810121(.x(x_121), .z(tmp00_121_81));
	booth__010 #(.WIDTH(WIDTH)) mul00810122(.x(x_122), .z(tmp00_122_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00810123(.x(x_123), .z(tmp00_123_81));
	booth__004 #(.WIDTH(WIDTH)) mul00810124(.x(x_124), .z(tmp00_124_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810125(.x(x_125), .z(tmp00_125_81));
	booth_0008 #(.WIDTH(WIDTH)) mul00810126(.x(x_126), .z(tmp00_126_81));
	booth_0004 #(.WIDTH(WIDTH)) mul00810127(.x(x_127), .z(tmp00_127_81));
	booth_0000 #(.WIDTH(WIDTH)) mul00820000(.x(x_0), .z(tmp00_0_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820001(.x(x_1), .z(tmp00_1_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820002(.x(x_2), .z(tmp00_2_82));
	booth_0006 #(.WIDTH(WIDTH)) mul00820003(.x(x_3), .z(tmp00_3_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820004(.x(x_4), .z(tmp00_4_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820005(.x(x_5), .z(tmp00_5_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820006(.x(x_6), .z(tmp00_6_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820007(.x(x_7), .z(tmp00_7_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820008(.x(x_8), .z(tmp00_8_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820009(.x(x_9), .z(tmp00_9_82));
	booth__002 #(.WIDTH(WIDTH)) mul00820010(.x(x_10), .z(tmp00_10_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820011(.x(x_11), .z(tmp00_11_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820012(.x(x_12), .z(tmp00_12_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820013(.x(x_13), .z(tmp00_13_82));
	booth_0010 #(.WIDTH(WIDTH)) mul00820014(.x(x_14), .z(tmp00_14_82));
	booth__012 #(.WIDTH(WIDTH)) mul00820015(.x(x_15), .z(tmp00_15_82));
	booth_0002 #(.WIDTH(WIDTH)) mul00820016(.x(x_16), .z(tmp00_16_82));
	booth_0012 #(.WIDTH(WIDTH)) mul00820017(.x(x_17), .z(tmp00_17_82));
	booth__006 #(.WIDTH(WIDTH)) mul00820018(.x(x_18), .z(tmp00_18_82));
	booth_0012 #(.WIDTH(WIDTH)) mul00820019(.x(x_19), .z(tmp00_19_82));
	booth_0006 #(.WIDTH(WIDTH)) mul00820020(.x(x_20), .z(tmp00_20_82));
	booth_0006 #(.WIDTH(WIDTH)) mul00820021(.x(x_21), .z(tmp00_21_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820022(.x(x_22), .z(tmp00_22_82));
	booth__002 #(.WIDTH(WIDTH)) mul00820023(.x(x_23), .z(tmp00_23_82));
	booth_0012 #(.WIDTH(WIDTH)) mul00820024(.x(x_24), .z(tmp00_24_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820025(.x(x_25), .z(tmp00_25_82));
	booth_0004 #(.WIDTH(WIDTH)) mul00820026(.x(x_26), .z(tmp00_26_82));
	booth__002 #(.WIDTH(WIDTH)) mul00820027(.x(x_27), .z(tmp00_27_82));
	booth_0006 #(.WIDTH(WIDTH)) mul00820028(.x(x_28), .z(tmp00_28_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820029(.x(x_29), .z(tmp00_29_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820030(.x(x_30), .z(tmp00_30_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820031(.x(x_31), .z(tmp00_31_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820032(.x(x_32), .z(tmp00_32_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820033(.x(x_33), .z(tmp00_33_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820034(.x(x_34), .z(tmp00_34_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820035(.x(x_35), .z(tmp00_35_82));
	booth__012 #(.WIDTH(WIDTH)) mul00820036(.x(x_36), .z(tmp00_36_82));
	booth_0004 #(.WIDTH(WIDTH)) mul00820037(.x(x_37), .z(tmp00_37_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820038(.x(x_38), .z(tmp00_38_82));
	booth_0014 #(.WIDTH(WIDTH)) mul00820039(.x(x_39), .z(tmp00_39_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820040(.x(x_40), .z(tmp00_40_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820041(.x(x_41), .z(tmp00_41_82));
	booth_0010 #(.WIDTH(WIDTH)) mul00820042(.x(x_42), .z(tmp00_42_82));
	booth_0014 #(.WIDTH(WIDTH)) mul00820043(.x(x_43), .z(tmp00_43_82));
	booth__012 #(.WIDTH(WIDTH)) mul00820044(.x(x_44), .z(tmp00_44_82));
	booth_0004 #(.WIDTH(WIDTH)) mul00820045(.x(x_45), .z(tmp00_45_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820046(.x(x_46), .z(tmp00_46_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820047(.x(x_47), .z(tmp00_47_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820048(.x(x_48), .z(tmp00_48_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820049(.x(x_49), .z(tmp00_49_82));
	booth_0010 #(.WIDTH(WIDTH)) mul00820050(.x(x_50), .z(tmp00_50_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820051(.x(x_51), .z(tmp00_51_82));
	booth_0012 #(.WIDTH(WIDTH)) mul00820052(.x(x_52), .z(tmp00_52_82));
	booth_0012 #(.WIDTH(WIDTH)) mul00820053(.x(x_53), .z(tmp00_53_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820054(.x(x_54), .z(tmp00_54_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820055(.x(x_55), .z(tmp00_55_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820056(.x(x_56), .z(tmp00_56_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820057(.x(x_57), .z(tmp00_57_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820058(.x(x_58), .z(tmp00_58_82));
	booth_0012 #(.WIDTH(WIDTH)) mul00820059(.x(x_59), .z(tmp00_59_82));
	booth__012 #(.WIDTH(WIDTH)) mul00820060(.x(x_60), .z(tmp00_60_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820061(.x(x_61), .z(tmp00_61_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820062(.x(x_62), .z(tmp00_62_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820063(.x(x_63), .z(tmp00_63_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820064(.x(x_64), .z(tmp00_64_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820065(.x(x_65), .z(tmp00_65_82));
	booth__002 #(.WIDTH(WIDTH)) mul00820066(.x(x_66), .z(tmp00_66_82));
	booth__006 #(.WIDTH(WIDTH)) mul00820067(.x(x_67), .z(tmp00_67_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820068(.x(x_68), .z(tmp00_68_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820069(.x(x_69), .z(tmp00_69_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820070(.x(x_70), .z(tmp00_70_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820071(.x(x_71), .z(tmp00_71_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820072(.x(x_72), .z(tmp00_72_82));
	booth__012 #(.WIDTH(WIDTH)) mul00820073(.x(x_73), .z(tmp00_73_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820074(.x(x_74), .z(tmp00_74_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820075(.x(x_75), .z(tmp00_75_82));
	booth__006 #(.WIDTH(WIDTH)) mul00820076(.x(x_76), .z(tmp00_76_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820077(.x(x_77), .z(tmp00_77_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820078(.x(x_78), .z(tmp00_78_82));
	booth_0006 #(.WIDTH(WIDTH)) mul00820079(.x(x_79), .z(tmp00_79_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820080(.x(x_80), .z(tmp00_80_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820081(.x(x_81), .z(tmp00_81_82));
	booth__012 #(.WIDTH(WIDTH)) mul00820082(.x(x_82), .z(tmp00_82_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820083(.x(x_83), .z(tmp00_83_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820084(.x(x_84), .z(tmp00_84_82));
	booth_0002 #(.WIDTH(WIDTH)) mul00820085(.x(x_85), .z(tmp00_85_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820086(.x(x_86), .z(tmp00_86_82));
	booth__002 #(.WIDTH(WIDTH)) mul00820087(.x(x_87), .z(tmp00_87_82));
	booth_0010 #(.WIDTH(WIDTH)) mul00820088(.x(x_88), .z(tmp00_88_82));
	booth__002 #(.WIDTH(WIDTH)) mul00820089(.x(x_89), .z(tmp00_89_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820090(.x(x_90), .z(tmp00_90_82));
	booth_0016 #(.WIDTH(WIDTH)) mul00820091(.x(x_91), .z(tmp00_91_82));
	booth_0006 #(.WIDTH(WIDTH)) mul00820092(.x(x_92), .z(tmp00_92_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820093(.x(x_93), .z(tmp00_93_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820094(.x(x_94), .z(tmp00_94_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820095(.x(x_95), .z(tmp00_95_82));
	booth_0006 #(.WIDTH(WIDTH)) mul00820096(.x(x_96), .z(tmp00_96_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820097(.x(x_97), .z(tmp00_97_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820098(.x(x_98), .z(tmp00_98_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820099(.x(x_99), .z(tmp00_99_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820100(.x(x_100), .z(tmp00_100_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820101(.x(x_101), .z(tmp00_101_82));
	booth_0004 #(.WIDTH(WIDTH)) mul00820102(.x(x_102), .z(tmp00_102_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820103(.x(x_103), .z(tmp00_103_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820104(.x(x_104), .z(tmp00_104_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820105(.x(x_105), .z(tmp00_105_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820106(.x(x_106), .z(tmp00_106_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820107(.x(x_107), .z(tmp00_107_82));
	booth_0004 #(.WIDTH(WIDTH)) mul00820108(.x(x_108), .z(tmp00_108_82));
	booth_0010 #(.WIDTH(WIDTH)) mul00820109(.x(x_109), .z(tmp00_109_82));
	booth_0004 #(.WIDTH(WIDTH)) mul00820110(.x(x_110), .z(tmp00_110_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820111(.x(x_111), .z(tmp00_111_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820112(.x(x_112), .z(tmp00_112_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820113(.x(x_113), .z(tmp00_113_82));
	booth__008 #(.WIDTH(WIDTH)) mul00820114(.x(x_114), .z(tmp00_114_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820115(.x(x_115), .z(tmp00_115_82));
	booth__010 #(.WIDTH(WIDTH)) mul00820116(.x(x_116), .z(tmp00_116_82));
	booth__002 #(.WIDTH(WIDTH)) mul00820117(.x(x_117), .z(tmp00_117_82));
	booth__010 #(.WIDTH(WIDTH)) mul00820118(.x(x_118), .z(tmp00_118_82));
	booth__016 #(.WIDTH(WIDTH)) mul00820119(.x(x_119), .z(tmp00_119_82));
	booth__002 #(.WIDTH(WIDTH)) mul00820120(.x(x_120), .z(tmp00_120_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820121(.x(x_121), .z(tmp00_121_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820122(.x(x_122), .z(tmp00_122_82));
	booth__004 #(.WIDTH(WIDTH)) mul00820123(.x(x_123), .z(tmp00_123_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820124(.x(x_124), .z(tmp00_124_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820125(.x(x_125), .z(tmp00_125_82));
	booth_0000 #(.WIDTH(WIDTH)) mul00820126(.x(x_126), .z(tmp00_126_82));
	booth_0008 #(.WIDTH(WIDTH)) mul00820127(.x(x_127), .z(tmp00_127_82));
	booth_0004 #(.WIDTH(WIDTH)) mul00830000(.x(x_0), .z(tmp00_0_83));
	booth__012 #(.WIDTH(WIDTH)) mul00830001(.x(x_1), .z(tmp00_1_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830002(.x(x_2), .z(tmp00_2_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830003(.x(x_3), .z(tmp00_3_83));
	booth_0016 #(.WIDTH(WIDTH)) mul00830004(.x(x_4), .z(tmp00_4_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830005(.x(x_5), .z(tmp00_5_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830006(.x(x_6), .z(tmp00_6_83));
	booth_0012 #(.WIDTH(WIDTH)) mul00830007(.x(x_7), .z(tmp00_7_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830008(.x(x_8), .z(tmp00_8_83));
	booth__010 #(.WIDTH(WIDTH)) mul00830009(.x(x_9), .z(tmp00_9_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830010(.x(x_10), .z(tmp00_10_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830011(.x(x_11), .z(tmp00_11_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830012(.x(x_12), .z(tmp00_12_83));
	booth__010 #(.WIDTH(WIDTH)) mul00830013(.x(x_13), .z(tmp00_13_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830014(.x(x_14), .z(tmp00_14_83));
	booth_0006 #(.WIDTH(WIDTH)) mul00830015(.x(x_15), .z(tmp00_15_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830016(.x(x_16), .z(tmp00_16_83));
	booth_0012 #(.WIDTH(WIDTH)) mul00830017(.x(x_17), .z(tmp00_17_83));
	booth_0002 #(.WIDTH(WIDTH)) mul00830018(.x(x_18), .z(tmp00_18_83));
	booth__002 #(.WIDTH(WIDTH)) mul00830019(.x(x_19), .z(tmp00_19_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830020(.x(x_20), .z(tmp00_20_83));
	booth__006 #(.WIDTH(WIDTH)) mul00830021(.x(x_21), .z(tmp00_21_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830022(.x(x_22), .z(tmp00_22_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830023(.x(x_23), .z(tmp00_23_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830024(.x(x_24), .z(tmp00_24_83));
	booth__012 #(.WIDTH(WIDTH)) mul00830025(.x(x_25), .z(tmp00_25_83));
	booth__012 #(.WIDTH(WIDTH)) mul00830026(.x(x_26), .z(tmp00_26_83));
	booth__012 #(.WIDTH(WIDTH)) mul00830027(.x(x_27), .z(tmp00_27_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830028(.x(x_28), .z(tmp00_28_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830029(.x(x_29), .z(tmp00_29_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830030(.x(x_30), .z(tmp00_30_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830031(.x(x_31), .z(tmp00_31_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830032(.x(x_32), .z(tmp00_32_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830033(.x(x_33), .z(tmp00_33_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830034(.x(x_34), .z(tmp00_34_83));
	booth_0010 #(.WIDTH(WIDTH)) mul00830035(.x(x_35), .z(tmp00_35_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830036(.x(x_36), .z(tmp00_36_83));
	booth__002 #(.WIDTH(WIDTH)) mul00830037(.x(x_37), .z(tmp00_37_83));
	booth_0012 #(.WIDTH(WIDTH)) mul00830038(.x(x_38), .z(tmp00_38_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830039(.x(x_39), .z(tmp00_39_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830040(.x(x_40), .z(tmp00_40_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830041(.x(x_41), .z(tmp00_41_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830042(.x(x_42), .z(tmp00_42_83));
	booth__006 #(.WIDTH(WIDTH)) mul00830043(.x(x_43), .z(tmp00_43_83));
	booth_0012 #(.WIDTH(WIDTH)) mul00830044(.x(x_44), .z(tmp00_44_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830045(.x(x_45), .z(tmp00_45_83));
	booth__014 #(.WIDTH(WIDTH)) mul00830046(.x(x_46), .z(tmp00_46_83));
	booth_0012 #(.WIDTH(WIDTH)) mul00830047(.x(x_47), .z(tmp00_47_83));
	booth_0012 #(.WIDTH(WIDTH)) mul00830048(.x(x_48), .z(tmp00_48_83));
	booth_0006 #(.WIDTH(WIDTH)) mul00830049(.x(x_49), .z(tmp00_49_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830050(.x(x_50), .z(tmp00_50_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830051(.x(x_51), .z(tmp00_51_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830052(.x(x_52), .z(tmp00_52_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830053(.x(x_53), .z(tmp00_53_83));
	booth_0012 #(.WIDTH(WIDTH)) mul00830054(.x(x_54), .z(tmp00_54_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830055(.x(x_55), .z(tmp00_55_83));
	booth__020 #(.WIDTH(WIDTH)) mul00830056(.x(x_56), .z(tmp00_56_83));
	booth__006 #(.WIDTH(WIDTH)) mul00830057(.x(x_57), .z(tmp00_57_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830058(.x(x_58), .z(tmp00_58_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830059(.x(x_59), .z(tmp00_59_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830060(.x(x_60), .z(tmp00_60_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830061(.x(x_61), .z(tmp00_61_83));
	booth_0006 #(.WIDTH(WIDTH)) mul00830062(.x(x_62), .z(tmp00_62_83));
	booth__012 #(.WIDTH(WIDTH)) mul00830063(.x(x_63), .z(tmp00_63_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830064(.x(x_64), .z(tmp00_64_83));
	booth_0006 #(.WIDTH(WIDTH)) mul00830065(.x(x_65), .z(tmp00_65_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830066(.x(x_66), .z(tmp00_66_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830067(.x(x_67), .z(tmp00_67_83));
	booth_0002 #(.WIDTH(WIDTH)) mul00830068(.x(x_68), .z(tmp00_68_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830069(.x(x_69), .z(tmp00_69_83));
	booth_0010 #(.WIDTH(WIDTH)) mul00830070(.x(x_70), .z(tmp00_70_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830071(.x(x_71), .z(tmp00_71_83));
	booth__010 #(.WIDTH(WIDTH)) mul00830072(.x(x_72), .z(tmp00_72_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830073(.x(x_73), .z(tmp00_73_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830074(.x(x_74), .z(tmp00_74_83));
	booth_0010 #(.WIDTH(WIDTH)) mul00830075(.x(x_75), .z(tmp00_75_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830076(.x(x_76), .z(tmp00_76_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830077(.x(x_77), .z(tmp00_77_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830078(.x(x_78), .z(tmp00_78_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830079(.x(x_79), .z(tmp00_79_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830080(.x(x_80), .z(tmp00_80_83));
	booth_0006 #(.WIDTH(WIDTH)) mul00830081(.x(x_81), .z(tmp00_81_83));
	booth_0016 #(.WIDTH(WIDTH)) mul00830082(.x(x_82), .z(tmp00_82_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830083(.x(x_83), .z(tmp00_83_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830084(.x(x_84), .z(tmp00_84_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830085(.x(x_85), .z(tmp00_85_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830086(.x(x_86), .z(tmp00_86_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830087(.x(x_87), .z(tmp00_87_83));
	booth__002 #(.WIDTH(WIDTH)) mul00830088(.x(x_88), .z(tmp00_88_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830089(.x(x_89), .z(tmp00_89_83));
	booth__016 #(.WIDTH(WIDTH)) mul00830090(.x(x_90), .z(tmp00_90_83));
	booth_0016 #(.WIDTH(WIDTH)) mul00830091(.x(x_91), .z(tmp00_91_83));
	booth_0014 #(.WIDTH(WIDTH)) mul00830092(.x(x_92), .z(tmp00_92_83));
	booth__010 #(.WIDTH(WIDTH)) mul00830093(.x(x_93), .z(tmp00_93_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830094(.x(x_94), .z(tmp00_94_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830095(.x(x_95), .z(tmp00_95_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830096(.x(x_96), .z(tmp00_96_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830097(.x(x_97), .z(tmp00_97_83));
	booth_0002 #(.WIDTH(WIDTH)) mul00830098(.x(x_98), .z(tmp00_98_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830099(.x(x_99), .z(tmp00_99_83));
	booth__010 #(.WIDTH(WIDTH)) mul00830100(.x(x_100), .z(tmp00_100_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830101(.x(x_101), .z(tmp00_101_83));
	booth_0014 #(.WIDTH(WIDTH)) mul00830102(.x(x_102), .z(tmp00_102_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830103(.x(x_103), .z(tmp00_103_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830104(.x(x_104), .z(tmp00_104_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830105(.x(x_105), .z(tmp00_105_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830106(.x(x_106), .z(tmp00_106_83));
	booth_0002 #(.WIDTH(WIDTH)) mul00830107(.x(x_107), .z(tmp00_107_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830108(.x(x_108), .z(tmp00_108_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830109(.x(x_109), .z(tmp00_109_83));
	booth_0006 #(.WIDTH(WIDTH)) mul00830110(.x(x_110), .z(tmp00_110_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830111(.x(x_111), .z(tmp00_111_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830112(.x(x_112), .z(tmp00_112_83));
	booth_0012 #(.WIDTH(WIDTH)) mul00830113(.x(x_113), .z(tmp00_113_83));
	booth__012 #(.WIDTH(WIDTH)) mul00830114(.x(x_114), .z(tmp00_114_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830115(.x(x_115), .z(tmp00_115_83));
	booth__008 #(.WIDTH(WIDTH)) mul00830116(.x(x_116), .z(tmp00_116_83));
	booth_0004 #(.WIDTH(WIDTH)) mul00830117(.x(x_117), .z(tmp00_117_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830118(.x(x_118), .z(tmp00_118_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830119(.x(x_119), .z(tmp00_119_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830120(.x(x_120), .z(tmp00_120_83));
	booth_0018 #(.WIDTH(WIDTH)) mul00830121(.x(x_121), .z(tmp00_121_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830122(.x(x_122), .z(tmp00_122_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830123(.x(x_123), .z(tmp00_123_83));
	booth_0000 #(.WIDTH(WIDTH)) mul00830124(.x(x_124), .z(tmp00_124_83));
	booth__004 #(.WIDTH(WIDTH)) mul00830125(.x(x_125), .z(tmp00_125_83));
	booth_0008 #(.WIDTH(WIDTH)) mul00830126(.x(x_126), .z(tmp00_126_83));
	booth__006 #(.WIDTH(WIDTH)) mul00830127(.x(x_127), .z(tmp00_127_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000000(.in0(tmp00_0_0), .in1(tmp00_1_0), .out(tmp01_0_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000001(.in0(tmp00_2_0), .in1(tmp00_3_0), .out(tmp01_1_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000002(.in0(tmp00_4_0), .in1(tmp00_5_0), .out(tmp01_2_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000003(.in0(tmp00_6_0), .in1(tmp00_7_0), .out(tmp01_3_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000004(.in0(tmp00_8_0), .in1(tmp00_9_0), .out(tmp01_4_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000005(.in0(tmp00_10_0), .in1(tmp00_11_0), .out(tmp01_5_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000006(.in0(tmp00_12_0), .in1(tmp00_13_0), .out(tmp01_6_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000007(.in0(tmp00_14_0), .in1(tmp00_15_0), .out(tmp01_7_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000008(.in0(tmp00_16_0), .in1(tmp00_17_0), .out(tmp01_8_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000009(.in0(tmp00_18_0), .in1(tmp00_19_0), .out(tmp01_9_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000010(.in0(tmp00_20_0), .in1(tmp00_21_0), .out(tmp01_10_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000011(.in0(tmp00_22_0), .in1(tmp00_23_0), .out(tmp01_11_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000012(.in0(tmp00_24_0), .in1(tmp00_25_0), .out(tmp01_12_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000013(.in0(tmp00_26_0), .in1(tmp00_27_0), .out(tmp01_13_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000014(.in0(tmp00_28_0), .in1(tmp00_29_0), .out(tmp01_14_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000015(.in0(tmp00_30_0), .in1(tmp00_31_0), .out(tmp01_15_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000016(.in0(tmp00_32_0), .in1(tmp00_33_0), .out(tmp01_16_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000017(.in0(tmp00_34_0), .in1(tmp00_35_0), .out(tmp01_17_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000018(.in0(tmp00_36_0), .in1(tmp00_37_0), .out(tmp01_18_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000019(.in0(tmp00_38_0), .in1(tmp00_39_0), .out(tmp01_19_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000020(.in0(tmp00_40_0), .in1(tmp00_41_0), .out(tmp01_20_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000021(.in0(tmp00_42_0), .in1(tmp00_43_0), .out(tmp01_21_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000022(.in0(tmp00_44_0), .in1(tmp00_45_0), .out(tmp01_22_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000023(.in0(tmp00_46_0), .in1(tmp00_47_0), .out(tmp01_23_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000024(.in0(tmp00_48_0), .in1(tmp00_49_0), .out(tmp01_24_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000025(.in0(tmp00_50_0), .in1(tmp00_51_0), .out(tmp01_25_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000026(.in0(tmp00_52_0), .in1(tmp00_53_0), .out(tmp01_26_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000027(.in0(tmp00_54_0), .in1(tmp00_55_0), .out(tmp01_27_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000028(.in0(tmp00_56_0), .in1(tmp00_57_0), .out(tmp01_28_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000029(.in0(tmp00_58_0), .in1(tmp00_59_0), .out(tmp01_29_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000030(.in0(tmp00_60_0), .in1(tmp00_61_0), .out(tmp01_30_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000031(.in0(tmp00_62_0), .in1(tmp00_63_0), .out(tmp01_31_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000032(.in0(tmp00_64_0), .in1(tmp00_65_0), .out(tmp01_32_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000033(.in0(tmp00_66_0), .in1(tmp00_67_0), .out(tmp01_33_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000034(.in0(tmp00_68_0), .in1(tmp00_69_0), .out(tmp01_34_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000035(.in0(tmp00_70_0), .in1(tmp00_71_0), .out(tmp01_35_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000036(.in0(tmp00_72_0), .in1(tmp00_73_0), .out(tmp01_36_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000037(.in0(tmp00_74_0), .in1(tmp00_75_0), .out(tmp01_37_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000038(.in0(tmp00_76_0), .in1(tmp00_77_0), .out(tmp01_38_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000039(.in0(tmp00_78_0), .in1(tmp00_79_0), .out(tmp01_39_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000040(.in0(tmp00_80_0), .in1(tmp00_81_0), .out(tmp01_40_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000041(.in0(tmp00_82_0), .in1(tmp00_83_0), .out(tmp01_41_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000042(.in0(tmp00_84_0), .in1(tmp00_85_0), .out(tmp01_42_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000043(.in0(tmp00_86_0), .in1(tmp00_87_0), .out(tmp01_43_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000044(.in0(tmp00_88_0), .in1(tmp00_89_0), .out(tmp01_44_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000045(.in0(tmp00_90_0), .in1(tmp00_91_0), .out(tmp01_45_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000046(.in0(tmp00_92_0), .in1(tmp00_93_0), .out(tmp01_46_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000047(.in0(tmp00_94_0), .in1(tmp00_95_0), .out(tmp01_47_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000048(.in0(tmp00_96_0), .in1(tmp00_97_0), .out(tmp01_48_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000049(.in0(tmp00_98_0), .in1(tmp00_99_0), .out(tmp01_49_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000050(.in0(tmp00_100_0), .in1(tmp00_101_0), .out(tmp01_50_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000051(.in0(tmp00_102_0), .in1(tmp00_103_0), .out(tmp01_51_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000052(.in0(tmp00_104_0), .in1(tmp00_105_0), .out(tmp01_52_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000053(.in0(tmp00_106_0), .in1(tmp00_107_0), .out(tmp01_53_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000054(.in0(tmp00_108_0), .in1(tmp00_109_0), .out(tmp01_54_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000055(.in0(tmp00_110_0), .in1(tmp00_111_0), .out(tmp01_55_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000056(.in0(tmp00_112_0), .in1(tmp00_113_0), .out(tmp01_56_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000057(.in0(tmp00_114_0), .in1(tmp00_115_0), .out(tmp01_57_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000058(.in0(tmp00_116_0), .in1(tmp00_117_0), .out(tmp01_58_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000059(.in0(tmp00_118_0), .in1(tmp00_119_0), .out(tmp01_59_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000060(.in0(tmp00_120_0), .in1(tmp00_121_0), .out(tmp01_60_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000061(.in0(tmp00_122_0), .in1(tmp00_123_0), .out(tmp01_61_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000062(.in0(tmp00_124_0), .in1(tmp00_125_0), .out(tmp01_62_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000063(.in0(tmp00_126_0), .in1(tmp00_127_0), .out(tmp01_63_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000064(.in0(tmp01_0_0), .in1(tmp01_1_0), .out(tmp02_0_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000065(.in0(tmp01_2_0), .in1(tmp01_3_0), .out(tmp02_1_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000066(.in0(tmp01_4_0), .in1(tmp01_5_0), .out(tmp02_2_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000067(.in0(tmp01_6_0), .in1(tmp01_7_0), .out(tmp02_3_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000068(.in0(tmp01_8_0), .in1(tmp01_9_0), .out(tmp02_4_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000069(.in0(tmp01_10_0), .in1(tmp01_11_0), .out(tmp02_5_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000070(.in0(tmp01_12_0), .in1(tmp01_13_0), .out(tmp02_6_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000071(.in0(tmp01_14_0), .in1(tmp01_15_0), .out(tmp02_7_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000072(.in0(tmp01_16_0), .in1(tmp01_17_0), .out(tmp02_8_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000073(.in0(tmp01_18_0), .in1(tmp01_19_0), .out(tmp02_9_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000074(.in0(tmp01_20_0), .in1(tmp01_21_0), .out(tmp02_10_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000075(.in0(tmp01_22_0), .in1(tmp01_23_0), .out(tmp02_11_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000076(.in0(tmp01_24_0), .in1(tmp01_25_0), .out(tmp02_12_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000077(.in0(tmp01_26_0), .in1(tmp01_27_0), .out(tmp02_13_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000078(.in0(tmp01_28_0), .in1(tmp01_29_0), .out(tmp02_14_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000079(.in0(tmp01_30_0), .in1(tmp01_31_0), .out(tmp02_15_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000080(.in0(tmp01_32_0), .in1(tmp01_33_0), .out(tmp02_16_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000081(.in0(tmp01_34_0), .in1(tmp01_35_0), .out(tmp02_17_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000082(.in0(tmp01_36_0), .in1(tmp01_37_0), .out(tmp02_18_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000083(.in0(tmp01_38_0), .in1(tmp01_39_0), .out(tmp02_19_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000084(.in0(tmp01_40_0), .in1(tmp01_41_0), .out(tmp02_20_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000085(.in0(tmp01_42_0), .in1(tmp01_43_0), .out(tmp02_21_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000086(.in0(tmp01_44_0), .in1(tmp01_45_0), .out(tmp02_22_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000087(.in0(tmp01_46_0), .in1(tmp01_47_0), .out(tmp02_23_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000088(.in0(tmp01_48_0), .in1(tmp01_49_0), .out(tmp02_24_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000089(.in0(tmp01_50_0), .in1(tmp01_51_0), .out(tmp02_25_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000090(.in0(tmp01_52_0), .in1(tmp01_53_0), .out(tmp02_26_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000091(.in0(tmp01_54_0), .in1(tmp01_55_0), .out(tmp02_27_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000092(.in0(tmp01_56_0), .in1(tmp01_57_0), .out(tmp02_28_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000093(.in0(tmp01_58_0), .in1(tmp01_59_0), .out(tmp02_29_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000094(.in0(tmp01_60_0), .in1(tmp01_61_0), .out(tmp02_30_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000095(.in0(tmp01_62_0), .in1(tmp01_63_0), .out(tmp02_31_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000096(.in0(tmp02_0_0), .in1(tmp02_1_0), .out(tmp03_0_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000097(.in0(tmp02_2_0), .in1(tmp02_3_0), .out(tmp03_1_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000098(.in0(tmp02_4_0), .in1(tmp02_5_0), .out(tmp03_2_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000099(.in0(tmp02_6_0), .in1(tmp02_7_0), .out(tmp03_3_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000100(.in0(tmp02_8_0), .in1(tmp02_9_0), .out(tmp03_4_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000101(.in0(tmp02_10_0), .in1(tmp02_11_0), .out(tmp03_5_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000102(.in0(tmp02_12_0), .in1(tmp02_13_0), .out(tmp03_6_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000103(.in0(tmp02_14_0), .in1(tmp02_15_0), .out(tmp03_7_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000104(.in0(tmp02_16_0), .in1(tmp02_17_0), .out(tmp03_8_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000105(.in0(tmp02_18_0), .in1(tmp02_19_0), .out(tmp03_9_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000106(.in0(tmp02_20_0), .in1(tmp02_21_0), .out(tmp03_10_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000107(.in0(tmp02_22_0), .in1(tmp02_23_0), .out(tmp03_11_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000108(.in0(tmp02_24_0), .in1(tmp02_25_0), .out(tmp03_12_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000109(.in0(tmp02_26_0), .in1(tmp02_27_0), .out(tmp03_13_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000110(.in0(tmp02_28_0), .in1(tmp02_29_0), .out(tmp03_14_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000111(.in0(tmp02_30_0), .in1(tmp02_31_0), .out(tmp03_15_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000112(.in0(tmp03_0_0), .in1(tmp03_1_0), .out(tmp04_0_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000113(.in0(tmp03_2_0), .in1(tmp03_3_0), .out(tmp04_1_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000114(.in0(tmp03_4_0), .in1(tmp03_5_0), .out(tmp04_2_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000115(.in0(tmp03_6_0), .in1(tmp03_7_0), .out(tmp04_3_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000116(.in0(tmp03_8_0), .in1(tmp03_9_0), .out(tmp04_4_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000117(.in0(tmp03_10_0), .in1(tmp03_11_0), .out(tmp04_5_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000118(.in0(tmp03_12_0), .in1(tmp03_13_0), .out(tmp04_6_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000119(.in0(tmp03_14_0), .in1(tmp03_15_0), .out(tmp04_7_0));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000120(.in0(tmp04_0_0), .in1(tmp04_1_0), .out(tmp05_0_0));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000121(.in0(tmp04_2_0), .in1(tmp04_3_0), .out(tmp05_1_0));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000122(.in0(tmp04_4_0), .in1(tmp04_5_0), .out(tmp05_2_0));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000123(.in0(tmp04_6_0), .in1(tmp04_7_0), .out(tmp05_3_0));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000124(.in0(tmp05_0_0), .in1(tmp05_1_0), .out(tmp06_0_0));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000125(.in0(tmp05_2_0), .in1(tmp05_3_0), .out(tmp06_1_0));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000126(.in0(tmp06_0_0), .in1(tmp06_1_0), .out(tmp07_0_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000127(.in0(tmp00_0_1), .in1(tmp00_1_1), .out(tmp01_0_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000128(.in0(tmp00_2_1), .in1(tmp00_3_1), .out(tmp01_1_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000129(.in0(tmp00_4_1), .in1(tmp00_5_1), .out(tmp01_2_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000130(.in0(tmp00_6_1), .in1(tmp00_7_1), .out(tmp01_3_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000131(.in0(tmp00_8_1), .in1(tmp00_9_1), .out(tmp01_4_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000132(.in0(tmp00_10_1), .in1(tmp00_11_1), .out(tmp01_5_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000133(.in0(tmp00_12_1), .in1(tmp00_13_1), .out(tmp01_6_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000134(.in0(tmp00_14_1), .in1(tmp00_15_1), .out(tmp01_7_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000135(.in0(tmp00_16_1), .in1(tmp00_17_1), .out(tmp01_8_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000136(.in0(tmp00_18_1), .in1(tmp00_19_1), .out(tmp01_9_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000137(.in0(tmp00_20_1), .in1(tmp00_21_1), .out(tmp01_10_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000138(.in0(tmp00_22_1), .in1(tmp00_23_1), .out(tmp01_11_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000139(.in0(tmp00_24_1), .in1(tmp00_25_1), .out(tmp01_12_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000140(.in0(tmp00_26_1), .in1(tmp00_27_1), .out(tmp01_13_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000141(.in0(tmp00_28_1), .in1(tmp00_29_1), .out(tmp01_14_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000142(.in0(tmp00_30_1), .in1(tmp00_31_1), .out(tmp01_15_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000143(.in0(tmp00_32_1), .in1(tmp00_33_1), .out(tmp01_16_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000144(.in0(tmp00_34_1), .in1(tmp00_35_1), .out(tmp01_17_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000145(.in0(tmp00_36_1), .in1(tmp00_37_1), .out(tmp01_18_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000146(.in0(tmp00_38_1), .in1(tmp00_39_1), .out(tmp01_19_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000147(.in0(tmp00_40_1), .in1(tmp00_41_1), .out(tmp01_20_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000148(.in0(tmp00_42_1), .in1(tmp00_43_1), .out(tmp01_21_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000149(.in0(tmp00_44_1), .in1(tmp00_45_1), .out(tmp01_22_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000150(.in0(tmp00_46_1), .in1(tmp00_47_1), .out(tmp01_23_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000151(.in0(tmp00_48_1), .in1(tmp00_49_1), .out(tmp01_24_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000152(.in0(tmp00_50_1), .in1(tmp00_51_1), .out(tmp01_25_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000153(.in0(tmp00_52_1), .in1(tmp00_53_1), .out(tmp01_26_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000154(.in0(tmp00_54_1), .in1(tmp00_55_1), .out(tmp01_27_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000155(.in0(tmp00_56_1), .in1(tmp00_57_1), .out(tmp01_28_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000156(.in0(tmp00_58_1), .in1(tmp00_59_1), .out(tmp01_29_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000157(.in0(tmp00_60_1), .in1(tmp00_61_1), .out(tmp01_30_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000158(.in0(tmp00_62_1), .in1(tmp00_63_1), .out(tmp01_31_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000159(.in0(tmp00_64_1), .in1(tmp00_65_1), .out(tmp01_32_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000160(.in0(tmp00_66_1), .in1(tmp00_67_1), .out(tmp01_33_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000161(.in0(tmp00_68_1), .in1(tmp00_69_1), .out(tmp01_34_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000162(.in0(tmp00_70_1), .in1(tmp00_71_1), .out(tmp01_35_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000163(.in0(tmp00_72_1), .in1(tmp00_73_1), .out(tmp01_36_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000164(.in0(tmp00_74_1), .in1(tmp00_75_1), .out(tmp01_37_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000165(.in0(tmp00_76_1), .in1(tmp00_77_1), .out(tmp01_38_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000166(.in0(tmp00_78_1), .in1(tmp00_79_1), .out(tmp01_39_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000167(.in0(tmp00_80_1), .in1(tmp00_81_1), .out(tmp01_40_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000168(.in0(tmp00_82_1), .in1(tmp00_83_1), .out(tmp01_41_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000169(.in0(tmp00_84_1), .in1(tmp00_85_1), .out(tmp01_42_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000170(.in0(tmp00_86_1), .in1(tmp00_87_1), .out(tmp01_43_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000171(.in0(tmp00_88_1), .in1(tmp00_89_1), .out(tmp01_44_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000172(.in0(tmp00_90_1), .in1(tmp00_91_1), .out(tmp01_45_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000173(.in0(tmp00_92_1), .in1(tmp00_93_1), .out(tmp01_46_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000174(.in0(tmp00_94_1), .in1(tmp00_95_1), .out(tmp01_47_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000175(.in0(tmp00_96_1), .in1(tmp00_97_1), .out(tmp01_48_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000176(.in0(tmp00_98_1), .in1(tmp00_99_1), .out(tmp01_49_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000177(.in0(tmp00_100_1), .in1(tmp00_101_1), .out(tmp01_50_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000178(.in0(tmp00_102_1), .in1(tmp00_103_1), .out(tmp01_51_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000179(.in0(tmp00_104_1), .in1(tmp00_105_1), .out(tmp01_52_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000180(.in0(tmp00_106_1), .in1(tmp00_107_1), .out(tmp01_53_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000181(.in0(tmp00_108_1), .in1(tmp00_109_1), .out(tmp01_54_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000182(.in0(tmp00_110_1), .in1(tmp00_111_1), .out(tmp01_55_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000183(.in0(tmp00_112_1), .in1(tmp00_113_1), .out(tmp01_56_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000184(.in0(tmp00_114_1), .in1(tmp00_115_1), .out(tmp01_57_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000185(.in0(tmp00_116_1), .in1(tmp00_117_1), .out(tmp01_58_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000186(.in0(tmp00_118_1), .in1(tmp00_119_1), .out(tmp01_59_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000187(.in0(tmp00_120_1), .in1(tmp00_121_1), .out(tmp01_60_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000188(.in0(tmp00_122_1), .in1(tmp00_123_1), .out(tmp01_61_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000189(.in0(tmp00_124_1), .in1(tmp00_125_1), .out(tmp01_62_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000190(.in0(tmp00_126_1), .in1(tmp00_127_1), .out(tmp01_63_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000191(.in0(tmp01_0_1), .in1(tmp01_1_1), .out(tmp02_0_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000192(.in0(tmp01_2_1), .in1(tmp01_3_1), .out(tmp02_1_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000193(.in0(tmp01_4_1), .in1(tmp01_5_1), .out(tmp02_2_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000194(.in0(tmp01_6_1), .in1(tmp01_7_1), .out(tmp02_3_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000195(.in0(tmp01_8_1), .in1(tmp01_9_1), .out(tmp02_4_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000196(.in0(tmp01_10_1), .in1(tmp01_11_1), .out(tmp02_5_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000197(.in0(tmp01_12_1), .in1(tmp01_13_1), .out(tmp02_6_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000198(.in0(tmp01_14_1), .in1(tmp01_15_1), .out(tmp02_7_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000199(.in0(tmp01_16_1), .in1(tmp01_17_1), .out(tmp02_8_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000200(.in0(tmp01_18_1), .in1(tmp01_19_1), .out(tmp02_9_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000201(.in0(tmp01_20_1), .in1(tmp01_21_1), .out(tmp02_10_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000202(.in0(tmp01_22_1), .in1(tmp01_23_1), .out(tmp02_11_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000203(.in0(tmp01_24_1), .in1(tmp01_25_1), .out(tmp02_12_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000204(.in0(tmp01_26_1), .in1(tmp01_27_1), .out(tmp02_13_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000205(.in0(tmp01_28_1), .in1(tmp01_29_1), .out(tmp02_14_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000206(.in0(tmp01_30_1), .in1(tmp01_31_1), .out(tmp02_15_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000207(.in0(tmp01_32_1), .in1(tmp01_33_1), .out(tmp02_16_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000208(.in0(tmp01_34_1), .in1(tmp01_35_1), .out(tmp02_17_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000209(.in0(tmp01_36_1), .in1(tmp01_37_1), .out(tmp02_18_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000210(.in0(tmp01_38_1), .in1(tmp01_39_1), .out(tmp02_19_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000211(.in0(tmp01_40_1), .in1(tmp01_41_1), .out(tmp02_20_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000212(.in0(tmp01_42_1), .in1(tmp01_43_1), .out(tmp02_21_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000213(.in0(tmp01_44_1), .in1(tmp01_45_1), .out(tmp02_22_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000214(.in0(tmp01_46_1), .in1(tmp01_47_1), .out(tmp02_23_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000215(.in0(tmp01_48_1), .in1(tmp01_49_1), .out(tmp02_24_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000216(.in0(tmp01_50_1), .in1(tmp01_51_1), .out(tmp02_25_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000217(.in0(tmp01_52_1), .in1(tmp01_53_1), .out(tmp02_26_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000218(.in0(tmp01_54_1), .in1(tmp01_55_1), .out(tmp02_27_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000219(.in0(tmp01_56_1), .in1(tmp01_57_1), .out(tmp02_28_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000220(.in0(tmp01_58_1), .in1(tmp01_59_1), .out(tmp02_29_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000221(.in0(tmp01_60_1), .in1(tmp01_61_1), .out(tmp02_30_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000222(.in0(tmp01_62_1), .in1(tmp01_63_1), .out(tmp02_31_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000223(.in0(tmp02_0_1), .in1(tmp02_1_1), .out(tmp03_0_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000224(.in0(tmp02_2_1), .in1(tmp02_3_1), .out(tmp03_1_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000225(.in0(tmp02_4_1), .in1(tmp02_5_1), .out(tmp03_2_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000226(.in0(tmp02_6_1), .in1(tmp02_7_1), .out(tmp03_3_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000227(.in0(tmp02_8_1), .in1(tmp02_9_1), .out(tmp03_4_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000228(.in0(tmp02_10_1), .in1(tmp02_11_1), .out(tmp03_5_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000229(.in0(tmp02_12_1), .in1(tmp02_13_1), .out(tmp03_6_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000230(.in0(tmp02_14_1), .in1(tmp02_15_1), .out(tmp03_7_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000231(.in0(tmp02_16_1), .in1(tmp02_17_1), .out(tmp03_8_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000232(.in0(tmp02_18_1), .in1(tmp02_19_1), .out(tmp03_9_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000233(.in0(tmp02_20_1), .in1(tmp02_21_1), .out(tmp03_10_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000234(.in0(tmp02_22_1), .in1(tmp02_23_1), .out(tmp03_11_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000235(.in0(tmp02_24_1), .in1(tmp02_25_1), .out(tmp03_12_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000236(.in0(tmp02_26_1), .in1(tmp02_27_1), .out(tmp03_13_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000237(.in0(tmp02_28_1), .in1(tmp02_29_1), .out(tmp03_14_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000238(.in0(tmp02_30_1), .in1(tmp02_31_1), .out(tmp03_15_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000239(.in0(tmp03_0_1), .in1(tmp03_1_1), .out(tmp04_0_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000240(.in0(tmp03_2_1), .in1(tmp03_3_1), .out(tmp04_1_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000241(.in0(tmp03_4_1), .in1(tmp03_5_1), .out(tmp04_2_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000242(.in0(tmp03_6_1), .in1(tmp03_7_1), .out(tmp04_3_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000243(.in0(tmp03_8_1), .in1(tmp03_9_1), .out(tmp04_4_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000244(.in0(tmp03_10_1), .in1(tmp03_11_1), .out(tmp04_5_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000245(.in0(tmp03_12_1), .in1(tmp03_13_1), .out(tmp04_6_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000246(.in0(tmp03_14_1), .in1(tmp03_15_1), .out(tmp04_7_1));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000247(.in0(tmp04_0_1), .in1(tmp04_1_1), .out(tmp05_0_1));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000248(.in0(tmp04_2_1), .in1(tmp04_3_1), .out(tmp05_1_1));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000249(.in0(tmp04_4_1), .in1(tmp04_5_1), .out(tmp05_2_1));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000250(.in0(tmp04_6_1), .in1(tmp04_7_1), .out(tmp05_3_1));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000251(.in0(tmp05_0_1), .in1(tmp05_1_1), .out(tmp06_0_1));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000252(.in0(tmp05_2_1), .in1(tmp05_3_1), .out(tmp06_1_1));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000253(.in0(tmp06_0_1), .in1(tmp06_1_1), .out(tmp07_0_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000254(.in0(tmp00_0_2), .in1(tmp00_1_2), .out(tmp01_0_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000255(.in0(tmp00_2_2), .in1(tmp00_3_2), .out(tmp01_1_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000256(.in0(tmp00_4_2), .in1(tmp00_5_2), .out(tmp01_2_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000257(.in0(tmp00_6_2), .in1(tmp00_7_2), .out(tmp01_3_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000258(.in0(tmp00_8_2), .in1(tmp00_9_2), .out(tmp01_4_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000259(.in0(tmp00_10_2), .in1(tmp00_11_2), .out(tmp01_5_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000260(.in0(tmp00_12_2), .in1(tmp00_13_2), .out(tmp01_6_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000261(.in0(tmp00_14_2), .in1(tmp00_15_2), .out(tmp01_7_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000262(.in0(tmp00_16_2), .in1(tmp00_17_2), .out(tmp01_8_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000263(.in0(tmp00_18_2), .in1(tmp00_19_2), .out(tmp01_9_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000264(.in0(tmp00_20_2), .in1(tmp00_21_2), .out(tmp01_10_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000265(.in0(tmp00_22_2), .in1(tmp00_23_2), .out(tmp01_11_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000266(.in0(tmp00_24_2), .in1(tmp00_25_2), .out(tmp01_12_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000267(.in0(tmp00_26_2), .in1(tmp00_27_2), .out(tmp01_13_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000268(.in0(tmp00_28_2), .in1(tmp00_29_2), .out(tmp01_14_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000269(.in0(tmp00_30_2), .in1(tmp00_31_2), .out(tmp01_15_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000270(.in0(tmp00_32_2), .in1(tmp00_33_2), .out(tmp01_16_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000271(.in0(tmp00_34_2), .in1(tmp00_35_2), .out(tmp01_17_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000272(.in0(tmp00_36_2), .in1(tmp00_37_2), .out(tmp01_18_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000273(.in0(tmp00_38_2), .in1(tmp00_39_2), .out(tmp01_19_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000274(.in0(tmp00_40_2), .in1(tmp00_41_2), .out(tmp01_20_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000275(.in0(tmp00_42_2), .in1(tmp00_43_2), .out(tmp01_21_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000276(.in0(tmp00_44_2), .in1(tmp00_45_2), .out(tmp01_22_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000277(.in0(tmp00_46_2), .in1(tmp00_47_2), .out(tmp01_23_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000278(.in0(tmp00_48_2), .in1(tmp00_49_2), .out(tmp01_24_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000279(.in0(tmp00_50_2), .in1(tmp00_51_2), .out(tmp01_25_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000280(.in0(tmp00_52_2), .in1(tmp00_53_2), .out(tmp01_26_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000281(.in0(tmp00_54_2), .in1(tmp00_55_2), .out(tmp01_27_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000282(.in0(tmp00_56_2), .in1(tmp00_57_2), .out(tmp01_28_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000283(.in0(tmp00_58_2), .in1(tmp00_59_2), .out(tmp01_29_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000284(.in0(tmp00_60_2), .in1(tmp00_61_2), .out(tmp01_30_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000285(.in0(tmp00_62_2), .in1(tmp00_63_2), .out(tmp01_31_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000286(.in0(tmp00_64_2), .in1(tmp00_65_2), .out(tmp01_32_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000287(.in0(tmp00_66_2), .in1(tmp00_67_2), .out(tmp01_33_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000288(.in0(tmp00_68_2), .in1(tmp00_69_2), .out(tmp01_34_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000289(.in0(tmp00_70_2), .in1(tmp00_71_2), .out(tmp01_35_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000290(.in0(tmp00_72_2), .in1(tmp00_73_2), .out(tmp01_36_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000291(.in0(tmp00_74_2), .in1(tmp00_75_2), .out(tmp01_37_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000292(.in0(tmp00_76_2), .in1(tmp00_77_2), .out(tmp01_38_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000293(.in0(tmp00_78_2), .in1(tmp00_79_2), .out(tmp01_39_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000294(.in0(tmp00_80_2), .in1(tmp00_81_2), .out(tmp01_40_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000295(.in0(tmp00_82_2), .in1(tmp00_83_2), .out(tmp01_41_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000296(.in0(tmp00_84_2), .in1(tmp00_85_2), .out(tmp01_42_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000297(.in0(tmp00_86_2), .in1(tmp00_87_2), .out(tmp01_43_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000298(.in0(tmp00_88_2), .in1(tmp00_89_2), .out(tmp01_44_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000299(.in0(tmp00_90_2), .in1(tmp00_91_2), .out(tmp01_45_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000300(.in0(tmp00_92_2), .in1(tmp00_93_2), .out(tmp01_46_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000301(.in0(tmp00_94_2), .in1(tmp00_95_2), .out(tmp01_47_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000302(.in0(tmp00_96_2), .in1(tmp00_97_2), .out(tmp01_48_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000303(.in0(tmp00_98_2), .in1(tmp00_99_2), .out(tmp01_49_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000304(.in0(tmp00_100_2), .in1(tmp00_101_2), .out(tmp01_50_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000305(.in0(tmp00_102_2), .in1(tmp00_103_2), .out(tmp01_51_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000306(.in0(tmp00_104_2), .in1(tmp00_105_2), .out(tmp01_52_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000307(.in0(tmp00_106_2), .in1(tmp00_107_2), .out(tmp01_53_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000308(.in0(tmp00_108_2), .in1(tmp00_109_2), .out(tmp01_54_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000309(.in0(tmp00_110_2), .in1(tmp00_111_2), .out(tmp01_55_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000310(.in0(tmp00_112_2), .in1(tmp00_113_2), .out(tmp01_56_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000311(.in0(tmp00_114_2), .in1(tmp00_115_2), .out(tmp01_57_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000312(.in0(tmp00_116_2), .in1(tmp00_117_2), .out(tmp01_58_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000313(.in0(tmp00_118_2), .in1(tmp00_119_2), .out(tmp01_59_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000314(.in0(tmp00_120_2), .in1(tmp00_121_2), .out(tmp01_60_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000315(.in0(tmp00_122_2), .in1(tmp00_123_2), .out(tmp01_61_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000316(.in0(tmp00_124_2), .in1(tmp00_125_2), .out(tmp01_62_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000317(.in0(tmp00_126_2), .in1(tmp00_127_2), .out(tmp01_63_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000318(.in0(tmp01_0_2), .in1(tmp01_1_2), .out(tmp02_0_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000319(.in0(tmp01_2_2), .in1(tmp01_3_2), .out(tmp02_1_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000320(.in0(tmp01_4_2), .in1(tmp01_5_2), .out(tmp02_2_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000321(.in0(tmp01_6_2), .in1(tmp01_7_2), .out(tmp02_3_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000322(.in0(tmp01_8_2), .in1(tmp01_9_2), .out(tmp02_4_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000323(.in0(tmp01_10_2), .in1(tmp01_11_2), .out(tmp02_5_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000324(.in0(tmp01_12_2), .in1(tmp01_13_2), .out(tmp02_6_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000325(.in0(tmp01_14_2), .in1(tmp01_15_2), .out(tmp02_7_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000326(.in0(tmp01_16_2), .in1(tmp01_17_2), .out(tmp02_8_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000327(.in0(tmp01_18_2), .in1(tmp01_19_2), .out(tmp02_9_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000328(.in0(tmp01_20_2), .in1(tmp01_21_2), .out(tmp02_10_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000329(.in0(tmp01_22_2), .in1(tmp01_23_2), .out(tmp02_11_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000330(.in0(tmp01_24_2), .in1(tmp01_25_2), .out(tmp02_12_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000331(.in0(tmp01_26_2), .in1(tmp01_27_2), .out(tmp02_13_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000332(.in0(tmp01_28_2), .in1(tmp01_29_2), .out(tmp02_14_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000333(.in0(tmp01_30_2), .in1(tmp01_31_2), .out(tmp02_15_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000334(.in0(tmp01_32_2), .in1(tmp01_33_2), .out(tmp02_16_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000335(.in0(tmp01_34_2), .in1(tmp01_35_2), .out(tmp02_17_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000336(.in0(tmp01_36_2), .in1(tmp01_37_2), .out(tmp02_18_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000337(.in0(tmp01_38_2), .in1(tmp01_39_2), .out(tmp02_19_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000338(.in0(tmp01_40_2), .in1(tmp01_41_2), .out(tmp02_20_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000339(.in0(tmp01_42_2), .in1(tmp01_43_2), .out(tmp02_21_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000340(.in0(tmp01_44_2), .in1(tmp01_45_2), .out(tmp02_22_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000341(.in0(tmp01_46_2), .in1(tmp01_47_2), .out(tmp02_23_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000342(.in0(tmp01_48_2), .in1(tmp01_49_2), .out(tmp02_24_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000343(.in0(tmp01_50_2), .in1(tmp01_51_2), .out(tmp02_25_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000344(.in0(tmp01_52_2), .in1(tmp01_53_2), .out(tmp02_26_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000345(.in0(tmp01_54_2), .in1(tmp01_55_2), .out(tmp02_27_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000346(.in0(tmp01_56_2), .in1(tmp01_57_2), .out(tmp02_28_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000347(.in0(tmp01_58_2), .in1(tmp01_59_2), .out(tmp02_29_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000348(.in0(tmp01_60_2), .in1(tmp01_61_2), .out(tmp02_30_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000349(.in0(tmp01_62_2), .in1(tmp01_63_2), .out(tmp02_31_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000350(.in0(tmp02_0_2), .in1(tmp02_1_2), .out(tmp03_0_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000351(.in0(tmp02_2_2), .in1(tmp02_3_2), .out(tmp03_1_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000352(.in0(tmp02_4_2), .in1(tmp02_5_2), .out(tmp03_2_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000353(.in0(tmp02_6_2), .in1(tmp02_7_2), .out(tmp03_3_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000354(.in0(tmp02_8_2), .in1(tmp02_9_2), .out(tmp03_4_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000355(.in0(tmp02_10_2), .in1(tmp02_11_2), .out(tmp03_5_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000356(.in0(tmp02_12_2), .in1(tmp02_13_2), .out(tmp03_6_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000357(.in0(tmp02_14_2), .in1(tmp02_15_2), .out(tmp03_7_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000358(.in0(tmp02_16_2), .in1(tmp02_17_2), .out(tmp03_8_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000359(.in0(tmp02_18_2), .in1(tmp02_19_2), .out(tmp03_9_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000360(.in0(tmp02_20_2), .in1(tmp02_21_2), .out(tmp03_10_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000361(.in0(tmp02_22_2), .in1(tmp02_23_2), .out(tmp03_11_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000362(.in0(tmp02_24_2), .in1(tmp02_25_2), .out(tmp03_12_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000363(.in0(tmp02_26_2), .in1(tmp02_27_2), .out(tmp03_13_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000364(.in0(tmp02_28_2), .in1(tmp02_29_2), .out(tmp03_14_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000365(.in0(tmp02_30_2), .in1(tmp02_31_2), .out(tmp03_15_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000366(.in0(tmp03_0_2), .in1(tmp03_1_2), .out(tmp04_0_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000367(.in0(tmp03_2_2), .in1(tmp03_3_2), .out(tmp04_1_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000368(.in0(tmp03_4_2), .in1(tmp03_5_2), .out(tmp04_2_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000369(.in0(tmp03_6_2), .in1(tmp03_7_2), .out(tmp04_3_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000370(.in0(tmp03_8_2), .in1(tmp03_9_2), .out(tmp04_4_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000371(.in0(tmp03_10_2), .in1(tmp03_11_2), .out(tmp04_5_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000372(.in0(tmp03_12_2), .in1(tmp03_13_2), .out(tmp04_6_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000373(.in0(tmp03_14_2), .in1(tmp03_15_2), .out(tmp04_7_2));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000374(.in0(tmp04_0_2), .in1(tmp04_1_2), .out(tmp05_0_2));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000375(.in0(tmp04_2_2), .in1(tmp04_3_2), .out(tmp05_1_2));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000376(.in0(tmp04_4_2), .in1(tmp04_5_2), .out(tmp05_2_2));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000377(.in0(tmp04_6_2), .in1(tmp04_7_2), .out(tmp05_3_2));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000378(.in0(tmp05_0_2), .in1(tmp05_1_2), .out(tmp06_0_2));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000379(.in0(tmp05_2_2), .in1(tmp05_3_2), .out(tmp06_1_2));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000380(.in0(tmp06_0_2), .in1(tmp06_1_2), .out(tmp07_0_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000381(.in0(tmp00_0_3), .in1(tmp00_1_3), .out(tmp01_0_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000382(.in0(tmp00_2_3), .in1(tmp00_3_3), .out(tmp01_1_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000383(.in0(tmp00_4_3), .in1(tmp00_5_3), .out(tmp01_2_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000384(.in0(tmp00_6_3), .in1(tmp00_7_3), .out(tmp01_3_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000385(.in0(tmp00_8_3), .in1(tmp00_9_3), .out(tmp01_4_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000386(.in0(tmp00_10_3), .in1(tmp00_11_3), .out(tmp01_5_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000387(.in0(tmp00_12_3), .in1(tmp00_13_3), .out(tmp01_6_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000388(.in0(tmp00_14_3), .in1(tmp00_15_3), .out(tmp01_7_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000389(.in0(tmp00_16_3), .in1(tmp00_17_3), .out(tmp01_8_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000390(.in0(tmp00_18_3), .in1(tmp00_19_3), .out(tmp01_9_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000391(.in0(tmp00_20_3), .in1(tmp00_21_3), .out(tmp01_10_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000392(.in0(tmp00_22_3), .in1(tmp00_23_3), .out(tmp01_11_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000393(.in0(tmp00_24_3), .in1(tmp00_25_3), .out(tmp01_12_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000394(.in0(tmp00_26_3), .in1(tmp00_27_3), .out(tmp01_13_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000395(.in0(tmp00_28_3), .in1(tmp00_29_3), .out(tmp01_14_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000396(.in0(tmp00_30_3), .in1(tmp00_31_3), .out(tmp01_15_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000397(.in0(tmp00_32_3), .in1(tmp00_33_3), .out(tmp01_16_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000398(.in0(tmp00_34_3), .in1(tmp00_35_3), .out(tmp01_17_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000399(.in0(tmp00_36_3), .in1(tmp00_37_3), .out(tmp01_18_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000400(.in0(tmp00_38_3), .in1(tmp00_39_3), .out(tmp01_19_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000401(.in0(tmp00_40_3), .in1(tmp00_41_3), .out(tmp01_20_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000402(.in0(tmp00_42_3), .in1(tmp00_43_3), .out(tmp01_21_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000403(.in0(tmp00_44_3), .in1(tmp00_45_3), .out(tmp01_22_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000404(.in0(tmp00_46_3), .in1(tmp00_47_3), .out(tmp01_23_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000405(.in0(tmp00_48_3), .in1(tmp00_49_3), .out(tmp01_24_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000406(.in0(tmp00_50_3), .in1(tmp00_51_3), .out(tmp01_25_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000407(.in0(tmp00_52_3), .in1(tmp00_53_3), .out(tmp01_26_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000408(.in0(tmp00_54_3), .in1(tmp00_55_3), .out(tmp01_27_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000409(.in0(tmp00_56_3), .in1(tmp00_57_3), .out(tmp01_28_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000410(.in0(tmp00_58_3), .in1(tmp00_59_3), .out(tmp01_29_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000411(.in0(tmp00_60_3), .in1(tmp00_61_3), .out(tmp01_30_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000412(.in0(tmp00_62_3), .in1(tmp00_63_3), .out(tmp01_31_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000413(.in0(tmp00_64_3), .in1(tmp00_65_3), .out(tmp01_32_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000414(.in0(tmp00_66_3), .in1(tmp00_67_3), .out(tmp01_33_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000415(.in0(tmp00_68_3), .in1(tmp00_69_3), .out(tmp01_34_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000416(.in0(tmp00_70_3), .in1(tmp00_71_3), .out(tmp01_35_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000417(.in0(tmp00_72_3), .in1(tmp00_73_3), .out(tmp01_36_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000418(.in0(tmp00_74_3), .in1(tmp00_75_3), .out(tmp01_37_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000419(.in0(tmp00_76_3), .in1(tmp00_77_3), .out(tmp01_38_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000420(.in0(tmp00_78_3), .in1(tmp00_79_3), .out(tmp01_39_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000421(.in0(tmp00_80_3), .in1(tmp00_81_3), .out(tmp01_40_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000422(.in0(tmp00_82_3), .in1(tmp00_83_3), .out(tmp01_41_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000423(.in0(tmp00_84_3), .in1(tmp00_85_3), .out(tmp01_42_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000424(.in0(tmp00_86_3), .in1(tmp00_87_3), .out(tmp01_43_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000425(.in0(tmp00_88_3), .in1(tmp00_89_3), .out(tmp01_44_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000426(.in0(tmp00_90_3), .in1(tmp00_91_3), .out(tmp01_45_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000427(.in0(tmp00_92_3), .in1(tmp00_93_3), .out(tmp01_46_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000428(.in0(tmp00_94_3), .in1(tmp00_95_3), .out(tmp01_47_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000429(.in0(tmp00_96_3), .in1(tmp00_97_3), .out(tmp01_48_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000430(.in0(tmp00_98_3), .in1(tmp00_99_3), .out(tmp01_49_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000431(.in0(tmp00_100_3), .in1(tmp00_101_3), .out(tmp01_50_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000432(.in0(tmp00_102_3), .in1(tmp00_103_3), .out(tmp01_51_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000433(.in0(tmp00_104_3), .in1(tmp00_105_3), .out(tmp01_52_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000434(.in0(tmp00_106_3), .in1(tmp00_107_3), .out(tmp01_53_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000435(.in0(tmp00_108_3), .in1(tmp00_109_3), .out(tmp01_54_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000436(.in0(tmp00_110_3), .in1(tmp00_111_3), .out(tmp01_55_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000437(.in0(tmp00_112_3), .in1(tmp00_113_3), .out(tmp01_56_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000438(.in0(tmp00_114_3), .in1(tmp00_115_3), .out(tmp01_57_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000439(.in0(tmp00_116_3), .in1(tmp00_117_3), .out(tmp01_58_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000440(.in0(tmp00_118_3), .in1(tmp00_119_3), .out(tmp01_59_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000441(.in0(tmp00_120_3), .in1(tmp00_121_3), .out(tmp01_60_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000442(.in0(tmp00_122_3), .in1(tmp00_123_3), .out(tmp01_61_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000443(.in0(tmp00_124_3), .in1(tmp00_125_3), .out(tmp01_62_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000444(.in0(tmp00_126_3), .in1(tmp00_127_3), .out(tmp01_63_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000445(.in0(tmp01_0_3), .in1(tmp01_1_3), .out(tmp02_0_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000446(.in0(tmp01_2_3), .in1(tmp01_3_3), .out(tmp02_1_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000447(.in0(tmp01_4_3), .in1(tmp01_5_3), .out(tmp02_2_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000448(.in0(tmp01_6_3), .in1(tmp01_7_3), .out(tmp02_3_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000449(.in0(tmp01_8_3), .in1(tmp01_9_3), .out(tmp02_4_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000450(.in0(tmp01_10_3), .in1(tmp01_11_3), .out(tmp02_5_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000451(.in0(tmp01_12_3), .in1(tmp01_13_3), .out(tmp02_6_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000452(.in0(tmp01_14_3), .in1(tmp01_15_3), .out(tmp02_7_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000453(.in0(tmp01_16_3), .in1(tmp01_17_3), .out(tmp02_8_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000454(.in0(tmp01_18_3), .in1(tmp01_19_3), .out(tmp02_9_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000455(.in0(tmp01_20_3), .in1(tmp01_21_3), .out(tmp02_10_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000456(.in0(tmp01_22_3), .in1(tmp01_23_3), .out(tmp02_11_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000457(.in0(tmp01_24_3), .in1(tmp01_25_3), .out(tmp02_12_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000458(.in0(tmp01_26_3), .in1(tmp01_27_3), .out(tmp02_13_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000459(.in0(tmp01_28_3), .in1(tmp01_29_3), .out(tmp02_14_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000460(.in0(tmp01_30_3), .in1(tmp01_31_3), .out(tmp02_15_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000461(.in0(tmp01_32_3), .in1(tmp01_33_3), .out(tmp02_16_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000462(.in0(tmp01_34_3), .in1(tmp01_35_3), .out(tmp02_17_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000463(.in0(tmp01_36_3), .in1(tmp01_37_3), .out(tmp02_18_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000464(.in0(tmp01_38_3), .in1(tmp01_39_3), .out(tmp02_19_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000465(.in0(tmp01_40_3), .in1(tmp01_41_3), .out(tmp02_20_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000466(.in0(tmp01_42_3), .in1(tmp01_43_3), .out(tmp02_21_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000467(.in0(tmp01_44_3), .in1(tmp01_45_3), .out(tmp02_22_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000468(.in0(tmp01_46_3), .in1(tmp01_47_3), .out(tmp02_23_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000469(.in0(tmp01_48_3), .in1(tmp01_49_3), .out(tmp02_24_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000470(.in0(tmp01_50_3), .in1(tmp01_51_3), .out(tmp02_25_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000471(.in0(tmp01_52_3), .in1(tmp01_53_3), .out(tmp02_26_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000472(.in0(tmp01_54_3), .in1(tmp01_55_3), .out(tmp02_27_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000473(.in0(tmp01_56_3), .in1(tmp01_57_3), .out(tmp02_28_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000474(.in0(tmp01_58_3), .in1(tmp01_59_3), .out(tmp02_29_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000475(.in0(tmp01_60_3), .in1(tmp01_61_3), .out(tmp02_30_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000476(.in0(tmp01_62_3), .in1(tmp01_63_3), .out(tmp02_31_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000477(.in0(tmp02_0_3), .in1(tmp02_1_3), .out(tmp03_0_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000478(.in0(tmp02_2_3), .in1(tmp02_3_3), .out(tmp03_1_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000479(.in0(tmp02_4_3), .in1(tmp02_5_3), .out(tmp03_2_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000480(.in0(tmp02_6_3), .in1(tmp02_7_3), .out(tmp03_3_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000481(.in0(tmp02_8_3), .in1(tmp02_9_3), .out(tmp03_4_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000482(.in0(tmp02_10_3), .in1(tmp02_11_3), .out(tmp03_5_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000483(.in0(tmp02_12_3), .in1(tmp02_13_3), .out(tmp03_6_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000484(.in0(tmp02_14_3), .in1(tmp02_15_3), .out(tmp03_7_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000485(.in0(tmp02_16_3), .in1(tmp02_17_3), .out(tmp03_8_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000486(.in0(tmp02_18_3), .in1(tmp02_19_3), .out(tmp03_9_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000487(.in0(tmp02_20_3), .in1(tmp02_21_3), .out(tmp03_10_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000488(.in0(tmp02_22_3), .in1(tmp02_23_3), .out(tmp03_11_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000489(.in0(tmp02_24_3), .in1(tmp02_25_3), .out(tmp03_12_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000490(.in0(tmp02_26_3), .in1(tmp02_27_3), .out(tmp03_13_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000491(.in0(tmp02_28_3), .in1(tmp02_29_3), .out(tmp03_14_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000492(.in0(tmp02_30_3), .in1(tmp02_31_3), .out(tmp03_15_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000493(.in0(tmp03_0_3), .in1(tmp03_1_3), .out(tmp04_0_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000494(.in0(tmp03_2_3), .in1(tmp03_3_3), .out(tmp04_1_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000495(.in0(tmp03_4_3), .in1(tmp03_5_3), .out(tmp04_2_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000496(.in0(tmp03_6_3), .in1(tmp03_7_3), .out(tmp04_3_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000497(.in0(tmp03_8_3), .in1(tmp03_9_3), .out(tmp04_4_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000498(.in0(tmp03_10_3), .in1(tmp03_11_3), .out(tmp04_5_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000499(.in0(tmp03_12_3), .in1(tmp03_13_3), .out(tmp04_6_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000500(.in0(tmp03_14_3), .in1(tmp03_15_3), .out(tmp04_7_3));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000501(.in0(tmp04_0_3), .in1(tmp04_1_3), .out(tmp05_0_3));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000502(.in0(tmp04_2_3), .in1(tmp04_3_3), .out(tmp05_1_3));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000503(.in0(tmp04_4_3), .in1(tmp04_5_3), .out(tmp05_2_3));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000504(.in0(tmp04_6_3), .in1(tmp04_7_3), .out(tmp05_3_3));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000505(.in0(tmp05_0_3), .in1(tmp05_1_3), .out(tmp06_0_3));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000506(.in0(tmp05_2_3), .in1(tmp05_3_3), .out(tmp06_1_3));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000507(.in0(tmp06_0_3), .in1(tmp06_1_3), .out(tmp07_0_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000508(.in0(tmp00_0_4), .in1(tmp00_1_4), .out(tmp01_0_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000509(.in0(tmp00_2_4), .in1(tmp00_3_4), .out(tmp01_1_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000510(.in0(tmp00_4_4), .in1(tmp00_5_4), .out(tmp01_2_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000511(.in0(tmp00_6_4), .in1(tmp00_7_4), .out(tmp01_3_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000512(.in0(tmp00_8_4), .in1(tmp00_9_4), .out(tmp01_4_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000513(.in0(tmp00_10_4), .in1(tmp00_11_4), .out(tmp01_5_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000514(.in0(tmp00_12_4), .in1(tmp00_13_4), .out(tmp01_6_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000515(.in0(tmp00_14_4), .in1(tmp00_15_4), .out(tmp01_7_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000516(.in0(tmp00_16_4), .in1(tmp00_17_4), .out(tmp01_8_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000517(.in0(tmp00_18_4), .in1(tmp00_19_4), .out(tmp01_9_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000518(.in0(tmp00_20_4), .in1(tmp00_21_4), .out(tmp01_10_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000519(.in0(tmp00_22_4), .in1(tmp00_23_4), .out(tmp01_11_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000520(.in0(tmp00_24_4), .in1(tmp00_25_4), .out(tmp01_12_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000521(.in0(tmp00_26_4), .in1(tmp00_27_4), .out(tmp01_13_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000522(.in0(tmp00_28_4), .in1(tmp00_29_4), .out(tmp01_14_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000523(.in0(tmp00_30_4), .in1(tmp00_31_4), .out(tmp01_15_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000524(.in0(tmp00_32_4), .in1(tmp00_33_4), .out(tmp01_16_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000525(.in0(tmp00_34_4), .in1(tmp00_35_4), .out(tmp01_17_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000526(.in0(tmp00_36_4), .in1(tmp00_37_4), .out(tmp01_18_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000527(.in0(tmp00_38_4), .in1(tmp00_39_4), .out(tmp01_19_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000528(.in0(tmp00_40_4), .in1(tmp00_41_4), .out(tmp01_20_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000529(.in0(tmp00_42_4), .in1(tmp00_43_4), .out(tmp01_21_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000530(.in0(tmp00_44_4), .in1(tmp00_45_4), .out(tmp01_22_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000531(.in0(tmp00_46_4), .in1(tmp00_47_4), .out(tmp01_23_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000532(.in0(tmp00_48_4), .in1(tmp00_49_4), .out(tmp01_24_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000533(.in0(tmp00_50_4), .in1(tmp00_51_4), .out(tmp01_25_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000534(.in0(tmp00_52_4), .in1(tmp00_53_4), .out(tmp01_26_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000535(.in0(tmp00_54_4), .in1(tmp00_55_4), .out(tmp01_27_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000536(.in0(tmp00_56_4), .in1(tmp00_57_4), .out(tmp01_28_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000537(.in0(tmp00_58_4), .in1(tmp00_59_4), .out(tmp01_29_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000538(.in0(tmp00_60_4), .in1(tmp00_61_4), .out(tmp01_30_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000539(.in0(tmp00_62_4), .in1(tmp00_63_4), .out(tmp01_31_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000540(.in0(tmp00_64_4), .in1(tmp00_65_4), .out(tmp01_32_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000541(.in0(tmp00_66_4), .in1(tmp00_67_4), .out(tmp01_33_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000542(.in0(tmp00_68_4), .in1(tmp00_69_4), .out(tmp01_34_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000543(.in0(tmp00_70_4), .in1(tmp00_71_4), .out(tmp01_35_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000544(.in0(tmp00_72_4), .in1(tmp00_73_4), .out(tmp01_36_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000545(.in0(tmp00_74_4), .in1(tmp00_75_4), .out(tmp01_37_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000546(.in0(tmp00_76_4), .in1(tmp00_77_4), .out(tmp01_38_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000547(.in0(tmp00_78_4), .in1(tmp00_79_4), .out(tmp01_39_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000548(.in0(tmp00_80_4), .in1(tmp00_81_4), .out(tmp01_40_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000549(.in0(tmp00_82_4), .in1(tmp00_83_4), .out(tmp01_41_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000550(.in0(tmp00_84_4), .in1(tmp00_85_4), .out(tmp01_42_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000551(.in0(tmp00_86_4), .in1(tmp00_87_4), .out(tmp01_43_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000552(.in0(tmp00_88_4), .in1(tmp00_89_4), .out(tmp01_44_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000553(.in0(tmp00_90_4), .in1(tmp00_91_4), .out(tmp01_45_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000554(.in0(tmp00_92_4), .in1(tmp00_93_4), .out(tmp01_46_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000555(.in0(tmp00_94_4), .in1(tmp00_95_4), .out(tmp01_47_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000556(.in0(tmp00_96_4), .in1(tmp00_97_4), .out(tmp01_48_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000557(.in0(tmp00_98_4), .in1(tmp00_99_4), .out(tmp01_49_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000558(.in0(tmp00_100_4), .in1(tmp00_101_4), .out(tmp01_50_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000559(.in0(tmp00_102_4), .in1(tmp00_103_4), .out(tmp01_51_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000560(.in0(tmp00_104_4), .in1(tmp00_105_4), .out(tmp01_52_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000561(.in0(tmp00_106_4), .in1(tmp00_107_4), .out(tmp01_53_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000562(.in0(tmp00_108_4), .in1(tmp00_109_4), .out(tmp01_54_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000563(.in0(tmp00_110_4), .in1(tmp00_111_4), .out(tmp01_55_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000564(.in0(tmp00_112_4), .in1(tmp00_113_4), .out(tmp01_56_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000565(.in0(tmp00_114_4), .in1(tmp00_115_4), .out(tmp01_57_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000566(.in0(tmp00_116_4), .in1(tmp00_117_4), .out(tmp01_58_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000567(.in0(tmp00_118_4), .in1(tmp00_119_4), .out(tmp01_59_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000568(.in0(tmp00_120_4), .in1(tmp00_121_4), .out(tmp01_60_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000569(.in0(tmp00_122_4), .in1(tmp00_123_4), .out(tmp01_61_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000570(.in0(tmp00_124_4), .in1(tmp00_125_4), .out(tmp01_62_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000571(.in0(tmp00_126_4), .in1(tmp00_127_4), .out(tmp01_63_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000572(.in0(tmp01_0_4), .in1(tmp01_1_4), .out(tmp02_0_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000573(.in0(tmp01_2_4), .in1(tmp01_3_4), .out(tmp02_1_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000574(.in0(tmp01_4_4), .in1(tmp01_5_4), .out(tmp02_2_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000575(.in0(tmp01_6_4), .in1(tmp01_7_4), .out(tmp02_3_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000576(.in0(tmp01_8_4), .in1(tmp01_9_4), .out(tmp02_4_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000577(.in0(tmp01_10_4), .in1(tmp01_11_4), .out(tmp02_5_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000578(.in0(tmp01_12_4), .in1(tmp01_13_4), .out(tmp02_6_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000579(.in0(tmp01_14_4), .in1(tmp01_15_4), .out(tmp02_7_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000580(.in0(tmp01_16_4), .in1(tmp01_17_4), .out(tmp02_8_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000581(.in0(tmp01_18_4), .in1(tmp01_19_4), .out(tmp02_9_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000582(.in0(tmp01_20_4), .in1(tmp01_21_4), .out(tmp02_10_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000583(.in0(tmp01_22_4), .in1(tmp01_23_4), .out(tmp02_11_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000584(.in0(tmp01_24_4), .in1(tmp01_25_4), .out(tmp02_12_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000585(.in0(tmp01_26_4), .in1(tmp01_27_4), .out(tmp02_13_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000586(.in0(tmp01_28_4), .in1(tmp01_29_4), .out(tmp02_14_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000587(.in0(tmp01_30_4), .in1(tmp01_31_4), .out(tmp02_15_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000588(.in0(tmp01_32_4), .in1(tmp01_33_4), .out(tmp02_16_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000589(.in0(tmp01_34_4), .in1(tmp01_35_4), .out(tmp02_17_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000590(.in0(tmp01_36_4), .in1(tmp01_37_4), .out(tmp02_18_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000591(.in0(tmp01_38_4), .in1(tmp01_39_4), .out(tmp02_19_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000592(.in0(tmp01_40_4), .in1(tmp01_41_4), .out(tmp02_20_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000593(.in0(tmp01_42_4), .in1(tmp01_43_4), .out(tmp02_21_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000594(.in0(tmp01_44_4), .in1(tmp01_45_4), .out(tmp02_22_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000595(.in0(tmp01_46_4), .in1(tmp01_47_4), .out(tmp02_23_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000596(.in0(tmp01_48_4), .in1(tmp01_49_4), .out(tmp02_24_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000597(.in0(tmp01_50_4), .in1(tmp01_51_4), .out(tmp02_25_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000598(.in0(tmp01_52_4), .in1(tmp01_53_4), .out(tmp02_26_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000599(.in0(tmp01_54_4), .in1(tmp01_55_4), .out(tmp02_27_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000600(.in0(tmp01_56_4), .in1(tmp01_57_4), .out(tmp02_28_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000601(.in0(tmp01_58_4), .in1(tmp01_59_4), .out(tmp02_29_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000602(.in0(tmp01_60_4), .in1(tmp01_61_4), .out(tmp02_30_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000603(.in0(tmp01_62_4), .in1(tmp01_63_4), .out(tmp02_31_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000604(.in0(tmp02_0_4), .in1(tmp02_1_4), .out(tmp03_0_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000605(.in0(tmp02_2_4), .in1(tmp02_3_4), .out(tmp03_1_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000606(.in0(tmp02_4_4), .in1(tmp02_5_4), .out(tmp03_2_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000607(.in0(tmp02_6_4), .in1(tmp02_7_4), .out(tmp03_3_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000608(.in0(tmp02_8_4), .in1(tmp02_9_4), .out(tmp03_4_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000609(.in0(tmp02_10_4), .in1(tmp02_11_4), .out(tmp03_5_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000610(.in0(tmp02_12_4), .in1(tmp02_13_4), .out(tmp03_6_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000611(.in0(tmp02_14_4), .in1(tmp02_15_4), .out(tmp03_7_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000612(.in0(tmp02_16_4), .in1(tmp02_17_4), .out(tmp03_8_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000613(.in0(tmp02_18_4), .in1(tmp02_19_4), .out(tmp03_9_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000614(.in0(tmp02_20_4), .in1(tmp02_21_4), .out(tmp03_10_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000615(.in0(tmp02_22_4), .in1(tmp02_23_4), .out(tmp03_11_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000616(.in0(tmp02_24_4), .in1(tmp02_25_4), .out(tmp03_12_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000617(.in0(tmp02_26_4), .in1(tmp02_27_4), .out(tmp03_13_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000618(.in0(tmp02_28_4), .in1(tmp02_29_4), .out(tmp03_14_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000619(.in0(tmp02_30_4), .in1(tmp02_31_4), .out(tmp03_15_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000620(.in0(tmp03_0_4), .in1(tmp03_1_4), .out(tmp04_0_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000621(.in0(tmp03_2_4), .in1(tmp03_3_4), .out(tmp04_1_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000622(.in0(tmp03_4_4), .in1(tmp03_5_4), .out(tmp04_2_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000623(.in0(tmp03_6_4), .in1(tmp03_7_4), .out(tmp04_3_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000624(.in0(tmp03_8_4), .in1(tmp03_9_4), .out(tmp04_4_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000625(.in0(tmp03_10_4), .in1(tmp03_11_4), .out(tmp04_5_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000626(.in0(tmp03_12_4), .in1(tmp03_13_4), .out(tmp04_6_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000627(.in0(tmp03_14_4), .in1(tmp03_15_4), .out(tmp04_7_4));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000628(.in0(tmp04_0_4), .in1(tmp04_1_4), .out(tmp05_0_4));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000629(.in0(tmp04_2_4), .in1(tmp04_3_4), .out(tmp05_1_4));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000630(.in0(tmp04_4_4), .in1(tmp04_5_4), .out(tmp05_2_4));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000631(.in0(tmp04_6_4), .in1(tmp04_7_4), .out(tmp05_3_4));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000632(.in0(tmp05_0_4), .in1(tmp05_1_4), .out(tmp06_0_4));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000633(.in0(tmp05_2_4), .in1(tmp05_3_4), .out(tmp06_1_4));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000634(.in0(tmp06_0_4), .in1(tmp06_1_4), .out(tmp07_0_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000635(.in0(tmp00_0_5), .in1(tmp00_1_5), .out(tmp01_0_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000636(.in0(tmp00_2_5), .in1(tmp00_3_5), .out(tmp01_1_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000637(.in0(tmp00_4_5), .in1(tmp00_5_5), .out(tmp01_2_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000638(.in0(tmp00_6_5), .in1(tmp00_7_5), .out(tmp01_3_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000639(.in0(tmp00_8_5), .in1(tmp00_9_5), .out(tmp01_4_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000640(.in0(tmp00_10_5), .in1(tmp00_11_5), .out(tmp01_5_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000641(.in0(tmp00_12_5), .in1(tmp00_13_5), .out(tmp01_6_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000642(.in0(tmp00_14_5), .in1(tmp00_15_5), .out(tmp01_7_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000643(.in0(tmp00_16_5), .in1(tmp00_17_5), .out(tmp01_8_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000644(.in0(tmp00_18_5), .in1(tmp00_19_5), .out(tmp01_9_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000645(.in0(tmp00_20_5), .in1(tmp00_21_5), .out(tmp01_10_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000646(.in0(tmp00_22_5), .in1(tmp00_23_5), .out(tmp01_11_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000647(.in0(tmp00_24_5), .in1(tmp00_25_5), .out(tmp01_12_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000648(.in0(tmp00_26_5), .in1(tmp00_27_5), .out(tmp01_13_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000649(.in0(tmp00_28_5), .in1(tmp00_29_5), .out(tmp01_14_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000650(.in0(tmp00_30_5), .in1(tmp00_31_5), .out(tmp01_15_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000651(.in0(tmp00_32_5), .in1(tmp00_33_5), .out(tmp01_16_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000652(.in0(tmp00_34_5), .in1(tmp00_35_5), .out(tmp01_17_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000653(.in0(tmp00_36_5), .in1(tmp00_37_5), .out(tmp01_18_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000654(.in0(tmp00_38_5), .in1(tmp00_39_5), .out(tmp01_19_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000655(.in0(tmp00_40_5), .in1(tmp00_41_5), .out(tmp01_20_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000656(.in0(tmp00_42_5), .in1(tmp00_43_5), .out(tmp01_21_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000657(.in0(tmp00_44_5), .in1(tmp00_45_5), .out(tmp01_22_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000658(.in0(tmp00_46_5), .in1(tmp00_47_5), .out(tmp01_23_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000659(.in0(tmp00_48_5), .in1(tmp00_49_5), .out(tmp01_24_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000660(.in0(tmp00_50_5), .in1(tmp00_51_5), .out(tmp01_25_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000661(.in0(tmp00_52_5), .in1(tmp00_53_5), .out(tmp01_26_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000662(.in0(tmp00_54_5), .in1(tmp00_55_5), .out(tmp01_27_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000663(.in0(tmp00_56_5), .in1(tmp00_57_5), .out(tmp01_28_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000664(.in0(tmp00_58_5), .in1(tmp00_59_5), .out(tmp01_29_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000665(.in0(tmp00_60_5), .in1(tmp00_61_5), .out(tmp01_30_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000666(.in0(tmp00_62_5), .in1(tmp00_63_5), .out(tmp01_31_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000667(.in0(tmp00_64_5), .in1(tmp00_65_5), .out(tmp01_32_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000668(.in0(tmp00_66_5), .in1(tmp00_67_5), .out(tmp01_33_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000669(.in0(tmp00_68_5), .in1(tmp00_69_5), .out(tmp01_34_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000670(.in0(tmp00_70_5), .in1(tmp00_71_5), .out(tmp01_35_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000671(.in0(tmp00_72_5), .in1(tmp00_73_5), .out(tmp01_36_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000672(.in0(tmp00_74_5), .in1(tmp00_75_5), .out(tmp01_37_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000673(.in0(tmp00_76_5), .in1(tmp00_77_5), .out(tmp01_38_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000674(.in0(tmp00_78_5), .in1(tmp00_79_5), .out(tmp01_39_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000675(.in0(tmp00_80_5), .in1(tmp00_81_5), .out(tmp01_40_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000676(.in0(tmp00_82_5), .in1(tmp00_83_5), .out(tmp01_41_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000677(.in0(tmp00_84_5), .in1(tmp00_85_5), .out(tmp01_42_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000678(.in0(tmp00_86_5), .in1(tmp00_87_5), .out(tmp01_43_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000679(.in0(tmp00_88_5), .in1(tmp00_89_5), .out(tmp01_44_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000680(.in0(tmp00_90_5), .in1(tmp00_91_5), .out(tmp01_45_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000681(.in0(tmp00_92_5), .in1(tmp00_93_5), .out(tmp01_46_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000682(.in0(tmp00_94_5), .in1(tmp00_95_5), .out(tmp01_47_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000683(.in0(tmp00_96_5), .in1(tmp00_97_5), .out(tmp01_48_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000684(.in0(tmp00_98_5), .in1(tmp00_99_5), .out(tmp01_49_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000685(.in0(tmp00_100_5), .in1(tmp00_101_5), .out(tmp01_50_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000686(.in0(tmp00_102_5), .in1(tmp00_103_5), .out(tmp01_51_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000687(.in0(tmp00_104_5), .in1(tmp00_105_5), .out(tmp01_52_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000688(.in0(tmp00_106_5), .in1(tmp00_107_5), .out(tmp01_53_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000689(.in0(tmp00_108_5), .in1(tmp00_109_5), .out(tmp01_54_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000690(.in0(tmp00_110_5), .in1(tmp00_111_5), .out(tmp01_55_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000691(.in0(tmp00_112_5), .in1(tmp00_113_5), .out(tmp01_56_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000692(.in0(tmp00_114_5), .in1(tmp00_115_5), .out(tmp01_57_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000693(.in0(tmp00_116_5), .in1(tmp00_117_5), .out(tmp01_58_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000694(.in0(tmp00_118_5), .in1(tmp00_119_5), .out(tmp01_59_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000695(.in0(tmp00_120_5), .in1(tmp00_121_5), .out(tmp01_60_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000696(.in0(tmp00_122_5), .in1(tmp00_123_5), .out(tmp01_61_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000697(.in0(tmp00_124_5), .in1(tmp00_125_5), .out(tmp01_62_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000698(.in0(tmp00_126_5), .in1(tmp00_127_5), .out(tmp01_63_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000699(.in0(tmp01_0_5), .in1(tmp01_1_5), .out(tmp02_0_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000700(.in0(tmp01_2_5), .in1(tmp01_3_5), .out(tmp02_1_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000701(.in0(tmp01_4_5), .in1(tmp01_5_5), .out(tmp02_2_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000702(.in0(tmp01_6_5), .in1(tmp01_7_5), .out(tmp02_3_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000703(.in0(tmp01_8_5), .in1(tmp01_9_5), .out(tmp02_4_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000704(.in0(tmp01_10_5), .in1(tmp01_11_5), .out(tmp02_5_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000705(.in0(tmp01_12_5), .in1(tmp01_13_5), .out(tmp02_6_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000706(.in0(tmp01_14_5), .in1(tmp01_15_5), .out(tmp02_7_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000707(.in0(tmp01_16_5), .in1(tmp01_17_5), .out(tmp02_8_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000708(.in0(tmp01_18_5), .in1(tmp01_19_5), .out(tmp02_9_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000709(.in0(tmp01_20_5), .in1(tmp01_21_5), .out(tmp02_10_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000710(.in0(tmp01_22_5), .in1(tmp01_23_5), .out(tmp02_11_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000711(.in0(tmp01_24_5), .in1(tmp01_25_5), .out(tmp02_12_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000712(.in0(tmp01_26_5), .in1(tmp01_27_5), .out(tmp02_13_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000713(.in0(tmp01_28_5), .in1(tmp01_29_5), .out(tmp02_14_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000714(.in0(tmp01_30_5), .in1(tmp01_31_5), .out(tmp02_15_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000715(.in0(tmp01_32_5), .in1(tmp01_33_5), .out(tmp02_16_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000716(.in0(tmp01_34_5), .in1(tmp01_35_5), .out(tmp02_17_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000717(.in0(tmp01_36_5), .in1(tmp01_37_5), .out(tmp02_18_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000718(.in0(tmp01_38_5), .in1(tmp01_39_5), .out(tmp02_19_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000719(.in0(tmp01_40_5), .in1(tmp01_41_5), .out(tmp02_20_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000720(.in0(tmp01_42_5), .in1(tmp01_43_5), .out(tmp02_21_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000721(.in0(tmp01_44_5), .in1(tmp01_45_5), .out(tmp02_22_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000722(.in0(tmp01_46_5), .in1(tmp01_47_5), .out(tmp02_23_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000723(.in0(tmp01_48_5), .in1(tmp01_49_5), .out(tmp02_24_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000724(.in0(tmp01_50_5), .in1(tmp01_51_5), .out(tmp02_25_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000725(.in0(tmp01_52_5), .in1(tmp01_53_5), .out(tmp02_26_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000726(.in0(tmp01_54_5), .in1(tmp01_55_5), .out(tmp02_27_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000727(.in0(tmp01_56_5), .in1(tmp01_57_5), .out(tmp02_28_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000728(.in0(tmp01_58_5), .in1(tmp01_59_5), .out(tmp02_29_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000729(.in0(tmp01_60_5), .in1(tmp01_61_5), .out(tmp02_30_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000730(.in0(tmp01_62_5), .in1(tmp01_63_5), .out(tmp02_31_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000731(.in0(tmp02_0_5), .in1(tmp02_1_5), .out(tmp03_0_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000732(.in0(tmp02_2_5), .in1(tmp02_3_5), .out(tmp03_1_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000733(.in0(tmp02_4_5), .in1(tmp02_5_5), .out(tmp03_2_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000734(.in0(tmp02_6_5), .in1(tmp02_7_5), .out(tmp03_3_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000735(.in0(tmp02_8_5), .in1(tmp02_9_5), .out(tmp03_4_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000736(.in0(tmp02_10_5), .in1(tmp02_11_5), .out(tmp03_5_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000737(.in0(tmp02_12_5), .in1(tmp02_13_5), .out(tmp03_6_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000738(.in0(tmp02_14_5), .in1(tmp02_15_5), .out(tmp03_7_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000739(.in0(tmp02_16_5), .in1(tmp02_17_5), .out(tmp03_8_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000740(.in0(tmp02_18_5), .in1(tmp02_19_5), .out(tmp03_9_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000741(.in0(tmp02_20_5), .in1(tmp02_21_5), .out(tmp03_10_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000742(.in0(tmp02_22_5), .in1(tmp02_23_5), .out(tmp03_11_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000743(.in0(tmp02_24_5), .in1(tmp02_25_5), .out(tmp03_12_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000744(.in0(tmp02_26_5), .in1(tmp02_27_5), .out(tmp03_13_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000745(.in0(tmp02_28_5), .in1(tmp02_29_5), .out(tmp03_14_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000746(.in0(tmp02_30_5), .in1(tmp02_31_5), .out(tmp03_15_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000747(.in0(tmp03_0_5), .in1(tmp03_1_5), .out(tmp04_0_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000748(.in0(tmp03_2_5), .in1(tmp03_3_5), .out(tmp04_1_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000749(.in0(tmp03_4_5), .in1(tmp03_5_5), .out(tmp04_2_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000750(.in0(tmp03_6_5), .in1(tmp03_7_5), .out(tmp04_3_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000751(.in0(tmp03_8_5), .in1(tmp03_9_5), .out(tmp04_4_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000752(.in0(tmp03_10_5), .in1(tmp03_11_5), .out(tmp04_5_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000753(.in0(tmp03_12_5), .in1(tmp03_13_5), .out(tmp04_6_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000754(.in0(tmp03_14_5), .in1(tmp03_15_5), .out(tmp04_7_5));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000755(.in0(tmp04_0_5), .in1(tmp04_1_5), .out(tmp05_0_5));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000756(.in0(tmp04_2_5), .in1(tmp04_3_5), .out(tmp05_1_5));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000757(.in0(tmp04_4_5), .in1(tmp04_5_5), .out(tmp05_2_5));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000758(.in0(tmp04_6_5), .in1(tmp04_7_5), .out(tmp05_3_5));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000759(.in0(tmp05_0_5), .in1(tmp05_1_5), .out(tmp06_0_5));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000760(.in0(tmp05_2_5), .in1(tmp05_3_5), .out(tmp06_1_5));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000761(.in0(tmp06_0_5), .in1(tmp06_1_5), .out(tmp07_0_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000762(.in0(tmp00_0_6), .in1(tmp00_1_6), .out(tmp01_0_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000763(.in0(tmp00_2_6), .in1(tmp00_3_6), .out(tmp01_1_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000764(.in0(tmp00_4_6), .in1(tmp00_5_6), .out(tmp01_2_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000765(.in0(tmp00_6_6), .in1(tmp00_7_6), .out(tmp01_3_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000766(.in0(tmp00_8_6), .in1(tmp00_9_6), .out(tmp01_4_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000767(.in0(tmp00_10_6), .in1(tmp00_11_6), .out(tmp01_5_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000768(.in0(tmp00_12_6), .in1(tmp00_13_6), .out(tmp01_6_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000769(.in0(tmp00_14_6), .in1(tmp00_15_6), .out(tmp01_7_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000770(.in0(tmp00_16_6), .in1(tmp00_17_6), .out(tmp01_8_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000771(.in0(tmp00_18_6), .in1(tmp00_19_6), .out(tmp01_9_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000772(.in0(tmp00_20_6), .in1(tmp00_21_6), .out(tmp01_10_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000773(.in0(tmp00_22_6), .in1(tmp00_23_6), .out(tmp01_11_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000774(.in0(tmp00_24_6), .in1(tmp00_25_6), .out(tmp01_12_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000775(.in0(tmp00_26_6), .in1(tmp00_27_6), .out(tmp01_13_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000776(.in0(tmp00_28_6), .in1(tmp00_29_6), .out(tmp01_14_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000777(.in0(tmp00_30_6), .in1(tmp00_31_6), .out(tmp01_15_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000778(.in0(tmp00_32_6), .in1(tmp00_33_6), .out(tmp01_16_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000779(.in0(tmp00_34_6), .in1(tmp00_35_6), .out(tmp01_17_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000780(.in0(tmp00_36_6), .in1(tmp00_37_6), .out(tmp01_18_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000781(.in0(tmp00_38_6), .in1(tmp00_39_6), .out(tmp01_19_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000782(.in0(tmp00_40_6), .in1(tmp00_41_6), .out(tmp01_20_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000783(.in0(tmp00_42_6), .in1(tmp00_43_6), .out(tmp01_21_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000784(.in0(tmp00_44_6), .in1(tmp00_45_6), .out(tmp01_22_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000785(.in0(tmp00_46_6), .in1(tmp00_47_6), .out(tmp01_23_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000786(.in0(tmp00_48_6), .in1(tmp00_49_6), .out(tmp01_24_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000787(.in0(tmp00_50_6), .in1(tmp00_51_6), .out(tmp01_25_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000788(.in0(tmp00_52_6), .in1(tmp00_53_6), .out(tmp01_26_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000789(.in0(tmp00_54_6), .in1(tmp00_55_6), .out(tmp01_27_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000790(.in0(tmp00_56_6), .in1(tmp00_57_6), .out(tmp01_28_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000791(.in0(tmp00_58_6), .in1(tmp00_59_6), .out(tmp01_29_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000792(.in0(tmp00_60_6), .in1(tmp00_61_6), .out(tmp01_30_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000793(.in0(tmp00_62_6), .in1(tmp00_63_6), .out(tmp01_31_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000794(.in0(tmp00_64_6), .in1(tmp00_65_6), .out(tmp01_32_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000795(.in0(tmp00_66_6), .in1(tmp00_67_6), .out(tmp01_33_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000796(.in0(tmp00_68_6), .in1(tmp00_69_6), .out(tmp01_34_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000797(.in0(tmp00_70_6), .in1(tmp00_71_6), .out(tmp01_35_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000798(.in0(tmp00_72_6), .in1(tmp00_73_6), .out(tmp01_36_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000799(.in0(tmp00_74_6), .in1(tmp00_75_6), .out(tmp01_37_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000800(.in0(tmp00_76_6), .in1(tmp00_77_6), .out(tmp01_38_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000801(.in0(tmp00_78_6), .in1(tmp00_79_6), .out(tmp01_39_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000802(.in0(tmp00_80_6), .in1(tmp00_81_6), .out(tmp01_40_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000803(.in0(tmp00_82_6), .in1(tmp00_83_6), .out(tmp01_41_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000804(.in0(tmp00_84_6), .in1(tmp00_85_6), .out(tmp01_42_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000805(.in0(tmp00_86_6), .in1(tmp00_87_6), .out(tmp01_43_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000806(.in0(tmp00_88_6), .in1(tmp00_89_6), .out(tmp01_44_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000807(.in0(tmp00_90_6), .in1(tmp00_91_6), .out(tmp01_45_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000808(.in0(tmp00_92_6), .in1(tmp00_93_6), .out(tmp01_46_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000809(.in0(tmp00_94_6), .in1(tmp00_95_6), .out(tmp01_47_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000810(.in0(tmp00_96_6), .in1(tmp00_97_6), .out(tmp01_48_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000811(.in0(tmp00_98_6), .in1(tmp00_99_6), .out(tmp01_49_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000812(.in0(tmp00_100_6), .in1(tmp00_101_6), .out(tmp01_50_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000813(.in0(tmp00_102_6), .in1(tmp00_103_6), .out(tmp01_51_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000814(.in0(tmp00_104_6), .in1(tmp00_105_6), .out(tmp01_52_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000815(.in0(tmp00_106_6), .in1(tmp00_107_6), .out(tmp01_53_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000816(.in0(tmp00_108_6), .in1(tmp00_109_6), .out(tmp01_54_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000817(.in0(tmp00_110_6), .in1(tmp00_111_6), .out(tmp01_55_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000818(.in0(tmp00_112_6), .in1(tmp00_113_6), .out(tmp01_56_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000819(.in0(tmp00_114_6), .in1(tmp00_115_6), .out(tmp01_57_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000820(.in0(tmp00_116_6), .in1(tmp00_117_6), .out(tmp01_58_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000821(.in0(tmp00_118_6), .in1(tmp00_119_6), .out(tmp01_59_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000822(.in0(tmp00_120_6), .in1(tmp00_121_6), .out(tmp01_60_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000823(.in0(tmp00_122_6), .in1(tmp00_123_6), .out(tmp01_61_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000824(.in0(tmp00_124_6), .in1(tmp00_125_6), .out(tmp01_62_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000825(.in0(tmp00_126_6), .in1(tmp00_127_6), .out(tmp01_63_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000826(.in0(tmp01_0_6), .in1(tmp01_1_6), .out(tmp02_0_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000827(.in0(tmp01_2_6), .in1(tmp01_3_6), .out(tmp02_1_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000828(.in0(tmp01_4_6), .in1(tmp01_5_6), .out(tmp02_2_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000829(.in0(tmp01_6_6), .in1(tmp01_7_6), .out(tmp02_3_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000830(.in0(tmp01_8_6), .in1(tmp01_9_6), .out(tmp02_4_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000831(.in0(tmp01_10_6), .in1(tmp01_11_6), .out(tmp02_5_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000832(.in0(tmp01_12_6), .in1(tmp01_13_6), .out(tmp02_6_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000833(.in0(tmp01_14_6), .in1(tmp01_15_6), .out(tmp02_7_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000834(.in0(tmp01_16_6), .in1(tmp01_17_6), .out(tmp02_8_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000835(.in0(tmp01_18_6), .in1(tmp01_19_6), .out(tmp02_9_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000836(.in0(tmp01_20_6), .in1(tmp01_21_6), .out(tmp02_10_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000837(.in0(tmp01_22_6), .in1(tmp01_23_6), .out(tmp02_11_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000838(.in0(tmp01_24_6), .in1(tmp01_25_6), .out(tmp02_12_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000839(.in0(tmp01_26_6), .in1(tmp01_27_6), .out(tmp02_13_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000840(.in0(tmp01_28_6), .in1(tmp01_29_6), .out(tmp02_14_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000841(.in0(tmp01_30_6), .in1(tmp01_31_6), .out(tmp02_15_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000842(.in0(tmp01_32_6), .in1(tmp01_33_6), .out(tmp02_16_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000843(.in0(tmp01_34_6), .in1(tmp01_35_6), .out(tmp02_17_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000844(.in0(tmp01_36_6), .in1(tmp01_37_6), .out(tmp02_18_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000845(.in0(tmp01_38_6), .in1(tmp01_39_6), .out(tmp02_19_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000846(.in0(tmp01_40_6), .in1(tmp01_41_6), .out(tmp02_20_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000847(.in0(tmp01_42_6), .in1(tmp01_43_6), .out(tmp02_21_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000848(.in0(tmp01_44_6), .in1(tmp01_45_6), .out(tmp02_22_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000849(.in0(tmp01_46_6), .in1(tmp01_47_6), .out(tmp02_23_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000850(.in0(tmp01_48_6), .in1(tmp01_49_6), .out(tmp02_24_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000851(.in0(tmp01_50_6), .in1(tmp01_51_6), .out(tmp02_25_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000852(.in0(tmp01_52_6), .in1(tmp01_53_6), .out(tmp02_26_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000853(.in0(tmp01_54_6), .in1(tmp01_55_6), .out(tmp02_27_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000854(.in0(tmp01_56_6), .in1(tmp01_57_6), .out(tmp02_28_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000855(.in0(tmp01_58_6), .in1(tmp01_59_6), .out(tmp02_29_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000856(.in0(tmp01_60_6), .in1(tmp01_61_6), .out(tmp02_30_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000857(.in0(tmp01_62_6), .in1(tmp01_63_6), .out(tmp02_31_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000858(.in0(tmp02_0_6), .in1(tmp02_1_6), .out(tmp03_0_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000859(.in0(tmp02_2_6), .in1(tmp02_3_6), .out(tmp03_1_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000860(.in0(tmp02_4_6), .in1(tmp02_5_6), .out(tmp03_2_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000861(.in0(tmp02_6_6), .in1(tmp02_7_6), .out(tmp03_3_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000862(.in0(tmp02_8_6), .in1(tmp02_9_6), .out(tmp03_4_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000863(.in0(tmp02_10_6), .in1(tmp02_11_6), .out(tmp03_5_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000864(.in0(tmp02_12_6), .in1(tmp02_13_6), .out(tmp03_6_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000865(.in0(tmp02_14_6), .in1(tmp02_15_6), .out(tmp03_7_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000866(.in0(tmp02_16_6), .in1(tmp02_17_6), .out(tmp03_8_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000867(.in0(tmp02_18_6), .in1(tmp02_19_6), .out(tmp03_9_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000868(.in0(tmp02_20_6), .in1(tmp02_21_6), .out(tmp03_10_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000869(.in0(tmp02_22_6), .in1(tmp02_23_6), .out(tmp03_11_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000870(.in0(tmp02_24_6), .in1(tmp02_25_6), .out(tmp03_12_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000871(.in0(tmp02_26_6), .in1(tmp02_27_6), .out(tmp03_13_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000872(.in0(tmp02_28_6), .in1(tmp02_29_6), .out(tmp03_14_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000873(.in0(tmp02_30_6), .in1(tmp02_31_6), .out(tmp03_15_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000874(.in0(tmp03_0_6), .in1(tmp03_1_6), .out(tmp04_0_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000875(.in0(tmp03_2_6), .in1(tmp03_3_6), .out(tmp04_1_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000876(.in0(tmp03_4_6), .in1(tmp03_5_6), .out(tmp04_2_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000877(.in0(tmp03_6_6), .in1(tmp03_7_6), .out(tmp04_3_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000878(.in0(tmp03_8_6), .in1(tmp03_9_6), .out(tmp04_4_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000879(.in0(tmp03_10_6), .in1(tmp03_11_6), .out(tmp04_5_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000880(.in0(tmp03_12_6), .in1(tmp03_13_6), .out(tmp04_6_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000881(.in0(tmp03_14_6), .in1(tmp03_15_6), .out(tmp04_7_6));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000882(.in0(tmp04_0_6), .in1(tmp04_1_6), .out(tmp05_0_6));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000883(.in0(tmp04_2_6), .in1(tmp04_3_6), .out(tmp05_1_6));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000884(.in0(tmp04_4_6), .in1(tmp04_5_6), .out(tmp05_2_6));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000885(.in0(tmp04_6_6), .in1(tmp04_7_6), .out(tmp05_3_6));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000886(.in0(tmp05_0_6), .in1(tmp05_1_6), .out(tmp06_0_6));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000887(.in0(tmp05_2_6), .in1(tmp05_3_6), .out(tmp06_1_6));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000888(.in0(tmp06_0_6), .in1(tmp06_1_6), .out(tmp07_0_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000889(.in0(tmp00_0_7), .in1(tmp00_1_7), .out(tmp01_0_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000890(.in0(tmp00_2_7), .in1(tmp00_3_7), .out(tmp01_1_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000891(.in0(tmp00_4_7), .in1(tmp00_5_7), .out(tmp01_2_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000892(.in0(tmp00_6_7), .in1(tmp00_7_7), .out(tmp01_3_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000893(.in0(tmp00_8_7), .in1(tmp00_9_7), .out(tmp01_4_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000894(.in0(tmp00_10_7), .in1(tmp00_11_7), .out(tmp01_5_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000895(.in0(tmp00_12_7), .in1(tmp00_13_7), .out(tmp01_6_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000896(.in0(tmp00_14_7), .in1(tmp00_15_7), .out(tmp01_7_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000897(.in0(tmp00_16_7), .in1(tmp00_17_7), .out(tmp01_8_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000898(.in0(tmp00_18_7), .in1(tmp00_19_7), .out(tmp01_9_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000899(.in0(tmp00_20_7), .in1(tmp00_21_7), .out(tmp01_10_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000900(.in0(tmp00_22_7), .in1(tmp00_23_7), .out(tmp01_11_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000901(.in0(tmp00_24_7), .in1(tmp00_25_7), .out(tmp01_12_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000902(.in0(tmp00_26_7), .in1(tmp00_27_7), .out(tmp01_13_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000903(.in0(tmp00_28_7), .in1(tmp00_29_7), .out(tmp01_14_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000904(.in0(tmp00_30_7), .in1(tmp00_31_7), .out(tmp01_15_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000905(.in0(tmp00_32_7), .in1(tmp00_33_7), .out(tmp01_16_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000906(.in0(tmp00_34_7), .in1(tmp00_35_7), .out(tmp01_17_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000907(.in0(tmp00_36_7), .in1(tmp00_37_7), .out(tmp01_18_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000908(.in0(tmp00_38_7), .in1(tmp00_39_7), .out(tmp01_19_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000909(.in0(tmp00_40_7), .in1(tmp00_41_7), .out(tmp01_20_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000910(.in0(tmp00_42_7), .in1(tmp00_43_7), .out(tmp01_21_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000911(.in0(tmp00_44_7), .in1(tmp00_45_7), .out(tmp01_22_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000912(.in0(tmp00_46_7), .in1(tmp00_47_7), .out(tmp01_23_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000913(.in0(tmp00_48_7), .in1(tmp00_49_7), .out(tmp01_24_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000914(.in0(tmp00_50_7), .in1(tmp00_51_7), .out(tmp01_25_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000915(.in0(tmp00_52_7), .in1(tmp00_53_7), .out(tmp01_26_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000916(.in0(tmp00_54_7), .in1(tmp00_55_7), .out(tmp01_27_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000917(.in0(tmp00_56_7), .in1(tmp00_57_7), .out(tmp01_28_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000918(.in0(tmp00_58_7), .in1(tmp00_59_7), .out(tmp01_29_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000919(.in0(tmp00_60_7), .in1(tmp00_61_7), .out(tmp01_30_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000920(.in0(tmp00_62_7), .in1(tmp00_63_7), .out(tmp01_31_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000921(.in0(tmp00_64_7), .in1(tmp00_65_7), .out(tmp01_32_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000922(.in0(tmp00_66_7), .in1(tmp00_67_7), .out(tmp01_33_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000923(.in0(tmp00_68_7), .in1(tmp00_69_7), .out(tmp01_34_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000924(.in0(tmp00_70_7), .in1(tmp00_71_7), .out(tmp01_35_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000925(.in0(tmp00_72_7), .in1(tmp00_73_7), .out(tmp01_36_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000926(.in0(tmp00_74_7), .in1(tmp00_75_7), .out(tmp01_37_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000927(.in0(tmp00_76_7), .in1(tmp00_77_7), .out(tmp01_38_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000928(.in0(tmp00_78_7), .in1(tmp00_79_7), .out(tmp01_39_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000929(.in0(tmp00_80_7), .in1(tmp00_81_7), .out(tmp01_40_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000930(.in0(tmp00_82_7), .in1(tmp00_83_7), .out(tmp01_41_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000931(.in0(tmp00_84_7), .in1(tmp00_85_7), .out(tmp01_42_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000932(.in0(tmp00_86_7), .in1(tmp00_87_7), .out(tmp01_43_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000933(.in0(tmp00_88_7), .in1(tmp00_89_7), .out(tmp01_44_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000934(.in0(tmp00_90_7), .in1(tmp00_91_7), .out(tmp01_45_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000935(.in0(tmp00_92_7), .in1(tmp00_93_7), .out(tmp01_46_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000936(.in0(tmp00_94_7), .in1(tmp00_95_7), .out(tmp01_47_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000937(.in0(tmp00_96_7), .in1(tmp00_97_7), .out(tmp01_48_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000938(.in0(tmp00_98_7), .in1(tmp00_99_7), .out(tmp01_49_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000939(.in0(tmp00_100_7), .in1(tmp00_101_7), .out(tmp01_50_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000940(.in0(tmp00_102_7), .in1(tmp00_103_7), .out(tmp01_51_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000941(.in0(tmp00_104_7), .in1(tmp00_105_7), .out(tmp01_52_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000942(.in0(tmp00_106_7), .in1(tmp00_107_7), .out(tmp01_53_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000943(.in0(tmp00_108_7), .in1(tmp00_109_7), .out(tmp01_54_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000944(.in0(tmp00_110_7), .in1(tmp00_111_7), .out(tmp01_55_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000945(.in0(tmp00_112_7), .in1(tmp00_113_7), .out(tmp01_56_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000946(.in0(tmp00_114_7), .in1(tmp00_115_7), .out(tmp01_57_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000947(.in0(tmp00_116_7), .in1(tmp00_117_7), .out(tmp01_58_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000948(.in0(tmp00_118_7), .in1(tmp00_119_7), .out(tmp01_59_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000949(.in0(tmp00_120_7), .in1(tmp00_121_7), .out(tmp01_60_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000950(.in0(tmp00_122_7), .in1(tmp00_123_7), .out(tmp01_61_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000951(.in0(tmp00_124_7), .in1(tmp00_125_7), .out(tmp01_62_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000952(.in0(tmp00_126_7), .in1(tmp00_127_7), .out(tmp01_63_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000953(.in0(tmp01_0_7), .in1(tmp01_1_7), .out(tmp02_0_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000954(.in0(tmp01_2_7), .in1(tmp01_3_7), .out(tmp02_1_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000955(.in0(tmp01_4_7), .in1(tmp01_5_7), .out(tmp02_2_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000956(.in0(tmp01_6_7), .in1(tmp01_7_7), .out(tmp02_3_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000957(.in0(tmp01_8_7), .in1(tmp01_9_7), .out(tmp02_4_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000958(.in0(tmp01_10_7), .in1(tmp01_11_7), .out(tmp02_5_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000959(.in0(tmp01_12_7), .in1(tmp01_13_7), .out(tmp02_6_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000960(.in0(tmp01_14_7), .in1(tmp01_15_7), .out(tmp02_7_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000961(.in0(tmp01_16_7), .in1(tmp01_17_7), .out(tmp02_8_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000962(.in0(tmp01_18_7), .in1(tmp01_19_7), .out(tmp02_9_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000963(.in0(tmp01_20_7), .in1(tmp01_21_7), .out(tmp02_10_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000964(.in0(tmp01_22_7), .in1(tmp01_23_7), .out(tmp02_11_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000965(.in0(tmp01_24_7), .in1(tmp01_25_7), .out(tmp02_12_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000966(.in0(tmp01_26_7), .in1(tmp01_27_7), .out(tmp02_13_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000967(.in0(tmp01_28_7), .in1(tmp01_29_7), .out(tmp02_14_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000968(.in0(tmp01_30_7), .in1(tmp01_31_7), .out(tmp02_15_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000969(.in0(tmp01_32_7), .in1(tmp01_33_7), .out(tmp02_16_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000970(.in0(tmp01_34_7), .in1(tmp01_35_7), .out(tmp02_17_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000971(.in0(tmp01_36_7), .in1(tmp01_37_7), .out(tmp02_18_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000972(.in0(tmp01_38_7), .in1(tmp01_39_7), .out(tmp02_19_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000973(.in0(tmp01_40_7), .in1(tmp01_41_7), .out(tmp02_20_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000974(.in0(tmp01_42_7), .in1(tmp01_43_7), .out(tmp02_21_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000975(.in0(tmp01_44_7), .in1(tmp01_45_7), .out(tmp02_22_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000976(.in0(tmp01_46_7), .in1(tmp01_47_7), .out(tmp02_23_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000977(.in0(tmp01_48_7), .in1(tmp01_49_7), .out(tmp02_24_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000978(.in0(tmp01_50_7), .in1(tmp01_51_7), .out(tmp02_25_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000979(.in0(tmp01_52_7), .in1(tmp01_53_7), .out(tmp02_26_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000980(.in0(tmp01_54_7), .in1(tmp01_55_7), .out(tmp02_27_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000981(.in0(tmp01_56_7), .in1(tmp01_57_7), .out(tmp02_28_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000982(.in0(tmp01_58_7), .in1(tmp01_59_7), .out(tmp02_29_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000983(.in0(tmp01_60_7), .in1(tmp01_61_7), .out(tmp02_30_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000984(.in0(tmp01_62_7), .in1(tmp01_63_7), .out(tmp02_31_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000985(.in0(tmp02_0_7), .in1(tmp02_1_7), .out(tmp03_0_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000986(.in0(tmp02_2_7), .in1(tmp02_3_7), .out(tmp03_1_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000987(.in0(tmp02_4_7), .in1(tmp02_5_7), .out(tmp03_2_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000988(.in0(tmp02_6_7), .in1(tmp02_7_7), .out(tmp03_3_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000989(.in0(tmp02_8_7), .in1(tmp02_9_7), .out(tmp03_4_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000990(.in0(tmp02_10_7), .in1(tmp02_11_7), .out(tmp03_5_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000991(.in0(tmp02_12_7), .in1(tmp02_13_7), .out(tmp03_6_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000992(.in0(tmp02_14_7), .in1(tmp02_15_7), .out(tmp03_7_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000993(.in0(tmp02_16_7), .in1(tmp02_17_7), .out(tmp03_8_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000994(.in0(tmp02_18_7), .in1(tmp02_19_7), .out(tmp03_9_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000995(.in0(tmp02_20_7), .in1(tmp02_21_7), .out(tmp03_10_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000996(.in0(tmp02_22_7), .in1(tmp02_23_7), .out(tmp03_11_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000997(.in0(tmp02_24_7), .in1(tmp02_25_7), .out(tmp03_12_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000998(.in0(tmp02_26_7), .in1(tmp02_27_7), .out(tmp03_13_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000999(.in0(tmp02_28_7), .in1(tmp02_29_7), .out(tmp03_14_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001000(.in0(tmp02_30_7), .in1(tmp02_31_7), .out(tmp03_15_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001001(.in0(tmp03_0_7), .in1(tmp03_1_7), .out(tmp04_0_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001002(.in0(tmp03_2_7), .in1(tmp03_3_7), .out(tmp04_1_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001003(.in0(tmp03_4_7), .in1(tmp03_5_7), .out(tmp04_2_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001004(.in0(tmp03_6_7), .in1(tmp03_7_7), .out(tmp04_3_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001005(.in0(tmp03_8_7), .in1(tmp03_9_7), .out(tmp04_4_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001006(.in0(tmp03_10_7), .in1(tmp03_11_7), .out(tmp04_5_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001007(.in0(tmp03_12_7), .in1(tmp03_13_7), .out(tmp04_6_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001008(.in0(tmp03_14_7), .in1(tmp03_15_7), .out(tmp04_7_7));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001009(.in0(tmp04_0_7), .in1(tmp04_1_7), .out(tmp05_0_7));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001010(.in0(tmp04_2_7), .in1(tmp04_3_7), .out(tmp05_1_7));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001011(.in0(tmp04_4_7), .in1(tmp04_5_7), .out(tmp05_2_7));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001012(.in0(tmp04_6_7), .in1(tmp04_7_7), .out(tmp05_3_7));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001013(.in0(tmp05_0_7), .in1(tmp05_1_7), .out(tmp06_0_7));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001014(.in0(tmp05_2_7), .in1(tmp05_3_7), .out(tmp06_1_7));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add001015(.in0(tmp06_0_7), .in1(tmp06_1_7), .out(tmp07_0_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001016(.in0(tmp00_0_8), .in1(tmp00_1_8), .out(tmp01_0_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001017(.in0(tmp00_2_8), .in1(tmp00_3_8), .out(tmp01_1_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001018(.in0(tmp00_4_8), .in1(tmp00_5_8), .out(tmp01_2_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001019(.in0(tmp00_6_8), .in1(tmp00_7_8), .out(tmp01_3_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001020(.in0(tmp00_8_8), .in1(tmp00_9_8), .out(tmp01_4_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001021(.in0(tmp00_10_8), .in1(tmp00_11_8), .out(tmp01_5_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001022(.in0(tmp00_12_8), .in1(tmp00_13_8), .out(tmp01_6_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001023(.in0(tmp00_14_8), .in1(tmp00_15_8), .out(tmp01_7_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001024(.in0(tmp00_16_8), .in1(tmp00_17_8), .out(tmp01_8_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001025(.in0(tmp00_18_8), .in1(tmp00_19_8), .out(tmp01_9_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001026(.in0(tmp00_20_8), .in1(tmp00_21_8), .out(tmp01_10_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001027(.in0(tmp00_22_8), .in1(tmp00_23_8), .out(tmp01_11_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001028(.in0(tmp00_24_8), .in1(tmp00_25_8), .out(tmp01_12_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001029(.in0(tmp00_26_8), .in1(tmp00_27_8), .out(tmp01_13_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001030(.in0(tmp00_28_8), .in1(tmp00_29_8), .out(tmp01_14_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001031(.in0(tmp00_30_8), .in1(tmp00_31_8), .out(tmp01_15_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001032(.in0(tmp00_32_8), .in1(tmp00_33_8), .out(tmp01_16_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001033(.in0(tmp00_34_8), .in1(tmp00_35_8), .out(tmp01_17_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001034(.in0(tmp00_36_8), .in1(tmp00_37_8), .out(tmp01_18_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001035(.in0(tmp00_38_8), .in1(tmp00_39_8), .out(tmp01_19_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001036(.in0(tmp00_40_8), .in1(tmp00_41_8), .out(tmp01_20_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001037(.in0(tmp00_42_8), .in1(tmp00_43_8), .out(tmp01_21_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001038(.in0(tmp00_44_8), .in1(tmp00_45_8), .out(tmp01_22_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001039(.in0(tmp00_46_8), .in1(tmp00_47_8), .out(tmp01_23_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001040(.in0(tmp00_48_8), .in1(tmp00_49_8), .out(tmp01_24_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001041(.in0(tmp00_50_8), .in1(tmp00_51_8), .out(tmp01_25_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001042(.in0(tmp00_52_8), .in1(tmp00_53_8), .out(tmp01_26_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001043(.in0(tmp00_54_8), .in1(tmp00_55_8), .out(tmp01_27_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001044(.in0(tmp00_56_8), .in1(tmp00_57_8), .out(tmp01_28_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001045(.in0(tmp00_58_8), .in1(tmp00_59_8), .out(tmp01_29_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001046(.in0(tmp00_60_8), .in1(tmp00_61_8), .out(tmp01_30_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001047(.in0(tmp00_62_8), .in1(tmp00_63_8), .out(tmp01_31_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001048(.in0(tmp00_64_8), .in1(tmp00_65_8), .out(tmp01_32_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001049(.in0(tmp00_66_8), .in1(tmp00_67_8), .out(tmp01_33_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001050(.in0(tmp00_68_8), .in1(tmp00_69_8), .out(tmp01_34_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001051(.in0(tmp00_70_8), .in1(tmp00_71_8), .out(tmp01_35_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001052(.in0(tmp00_72_8), .in1(tmp00_73_8), .out(tmp01_36_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001053(.in0(tmp00_74_8), .in1(tmp00_75_8), .out(tmp01_37_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001054(.in0(tmp00_76_8), .in1(tmp00_77_8), .out(tmp01_38_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001055(.in0(tmp00_78_8), .in1(tmp00_79_8), .out(tmp01_39_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001056(.in0(tmp00_80_8), .in1(tmp00_81_8), .out(tmp01_40_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001057(.in0(tmp00_82_8), .in1(tmp00_83_8), .out(tmp01_41_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001058(.in0(tmp00_84_8), .in1(tmp00_85_8), .out(tmp01_42_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001059(.in0(tmp00_86_8), .in1(tmp00_87_8), .out(tmp01_43_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001060(.in0(tmp00_88_8), .in1(tmp00_89_8), .out(tmp01_44_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001061(.in0(tmp00_90_8), .in1(tmp00_91_8), .out(tmp01_45_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001062(.in0(tmp00_92_8), .in1(tmp00_93_8), .out(tmp01_46_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001063(.in0(tmp00_94_8), .in1(tmp00_95_8), .out(tmp01_47_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001064(.in0(tmp00_96_8), .in1(tmp00_97_8), .out(tmp01_48_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001065(.in0(tmp00_98_8), .in1(tmp00_99_8), .out(tmp01_49_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001066(.in0(tmp00_100_8), .in1(tmp00_101_8), .out(tmp01_50_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001067(.in0(tmp00_102_8), .in1(tmp00_103_8), .out(tmp01_51_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001068(.in0(tmp00_104_8), .in1(tmp00_105_8), .out(tmp01_52_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001069(.in0(tmp00_106_8), .in1(tmp00_107_8), .out(tmp01_53_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001070(.in0(tmp00_108_8), .in1(tmp00_109_8), .out(tmp01_54_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001071(.in0(tmp00_110_8), .in1(tmp00_111_8), .out(tmp01_55_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001072(.in0(tmp00_112_8), .in1(tmp00_113_8), .out(tmp01_56_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001073(.in0(tmp00_114_8), .in1(tmp00_115_8), .out(tmp01_57_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001074(.in0(tmp00_116_8), .in1(tmp00_117_8), .out(tmp01_58_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001075(.in0(tmp00_118_8), .in1(tmp00_119_8), .out(tmp01_59_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001076(.in0(tmp00_120_8), .in1(tmp00_121_8), .out(tmp01_60_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001077(.in0(tmp00_122_8), .in1(tmp00_123_8), .out(tmp01_61_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001078(.in0(tmp00_124_8), .in1(tmp00_125_8), .out(tmp01_62_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001079(.in0(tmp00_126_8), .in1(tmp00_127_8), .out(tmp01_63_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001080(.in0(tmp01_0_8), .in1(tmp01_1_8), .out(tmp02_0_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001081(.in0(tmp01_2_8), .in1(tmp01_3_8), .out(tmp02_1_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001082(.in0(tmp01_4_8), .in1(tmp01_5_8), .out(tmp02_2_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001083(.in0(tmp01_6_8), .in1(tmp01_7_8), .out(tmp02_3_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001084(.in0(tmp01_8_8), .in1(tmp01_9_8), .out(tmp02_4_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001085(.in0(tmp01_10_8), .in1(tmp01_11_8), .out(tmp02_5_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001086(.in0(tmp01_12_8), .in1(tmp01_13_8), .out(tmp02_6_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001087(.in0(tmp01_14_8), .in1(tmp01_15_8), .out(tmp02_7_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001088(.in0(tmp01_16_8), .in1(tmp01_17_8), .out(tmp02_8_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001089(.in0(tmp01_18_8), .in1(tmp01_19_8), .out(tmp02_9_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001090(.in0(tmp01_20_8), .in1(tmp01_21_8), .out(tmp02_10_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001091(.in0(tmp01_22_8), .in1(tmp01_23_8), .out(tmp02_11_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001092(.in0(tmp01_24_8), .in1(tmp01_25_8), .out(tmp02_12_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001093(.in0(tmp01_26_8), .in1(tmp01_27_8), .out(tmp02_13_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001094(.in0(tmp01_28_8), .in1(tmp01_29_8), .out(tmp02_14_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001095(.in0(tmp01_30_8), .in1(tmp01_31_8), .out(tmp02_15_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001096(.in0(tmp01_32_8), .in1(tmp01_33_8), .out(tmp02_16_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001097(.in0(tmp01_34_8), .in1(tmp01_35_8), .out(tmp02_17_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001098(.in0(tmp01_36_8), .in1(tmp01_37_8), .out(tmp02_18_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001099(.in0(tmp01_38_8), .in1(tmp01_39_8), .out(tmp02_19_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001100(.in0(tmp01_40_8), .in1(tmp01_41_8), .out(tmp02_20_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001101(.in0(tmp01_42_8), .in1(tmp01_43_8), .out(tmp02_21_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001102(.in0(tmp01_44_8), .in1(tmp01_45_8), .out(tmp02_22_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001103(.in0(tmp01_46_8), .in1(tmp01_47_8), .out(tmp02_23_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001104(.in0(tmp01_48_8), .in1(tmp01_49_8), .out(tmp02_24_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001105(.in0(tmp01_50_8), .in1(tmp01_51_8), .out(tmp02_25_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001106(.in0(tmp01_52_8), .in1(tmp01_53_8), .out(tmp02_26_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001107(.in0(tmp01_54_8), .in1(tmp01_55_8), .out(tmp02_27_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001108(.in0(tmp01_56_8), .in1(tmp01_57_8), .out(tmp02_28_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001109(.in0(tmp01_58_8), .in1(tmp01_59_8), .out(tmp02_29_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001110(.in0(tmp01_60_8), .in1(tmp01_61_8), .out(tmp02_30_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001111(.in0(tmp01_62_8), .in1(tmp01_63_8), .out(tmp02_31_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001112(.in0(tmp02_0_8), .in1(tmp02_1_8), .out(tmp03_0_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001113(.in0(tmp02_2_8), .in1(tmp02_3_8), .out(tmp03_1_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001114(.in0(tmp02_4_8), .in1(tmp02_5_8), .out(tmp03_2_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001115(.in0(tmp02_6_8), .in1(tmp02_7_8), .out(tmp03_3_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001116(.in0(tmp02_8_8), .in1(tmp02_9_8), .out(tmp03_4_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001117(.in0(tmp02_10_8), .in1(tmp02_11_8), .out(tmp03_5_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001118(.in0(tmp02_12_8), .in1(tmp02_13_8), .out(tmp03_6_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001119(.in0(tmp02_14_8), .in1(tmp02_15_8), .out(tmp03_7_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001120(.in0(tmp02_16_8), .in1(tmp02_17_8), .out(tmp03_8_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001121(.in0(tmp02_18_8), .in1(tmp02_19_8), .out(tmp03_9_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001122(.in0(tmp02_20_8), .in1(tmp02_21_8), .out(tmp03_10_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001123(.in0(tmp02_22_8), .in1(tmp02_23_8), .out(tmp03_11_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001124(.in0(tmp02_24_8), .in1(tmp02_25_8), .out(tmp03_12_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001125(.in0(tmp02_26_8), .in1(tmp02_27_8), .out(tmp03_13_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001126(.in0(tmp02_28_8), .in1(tmp02_29_8), .out(tmp03_14_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001127(.in0(tmp02_30_8), .in1(tmp02_31_8), .out(tmp03_15_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001128(.in0(tmp03_0_8), .in1(tmp03_1_8), .out(tmp04_0_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001129(.in0(tmp03_2_8), .in1(tmp03_3_8), .out(tmp04_1_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001130(.in0(tmp03_4_8), .in1(tmp03_5_8), .out(tmp04_2_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001131(.in0(tmp03_6_8), .in1(tmp03_7_8), .out(tmp04_3_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001132(.in0(tmp03_8_8), .in1(tmp03_9_8), .out(tmp04_4_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001133(.in0(tmp03_10_8), .in1(tmp03_11_8), .out(tmp04_5_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001134(.in0(tmp03_12_8), .in1(tmp03_13_8), .out(tmp04_6_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001135(.in0(tmp03_14_8), .in1(tmp03_15_8), .out(tmp04_7_8));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001136(.in0(tmp04_0_8), .in1(tmp04_1_8), .out(tmp05_0_8));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001137(.in0(tmp04_2_8), .in1(tmp04_3_8), .out(tmp05_1_8));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001138(.in0(tmp04_4_8), .in1(tmp04_5_8), .out(tmp05_2_8));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001139(.in0(tmp04_6_8), .in1(tmp04_7_8), .out(tmp05_3_8));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001140(.in0(tmp05_0_8), .in1(tmp05_1_8), .out(tmp06_0_8));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001141(.in0(tmp05_2_8), .in1(tmp05_3_8), .out(tmp06_1_8));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add001142(.in0(tmp06_0_8), .in1(tmp06_1_8), .out(tmp07_0_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001143(.in0(tmp00_0_9), .in1(tmp00_1_9), .out(tmp01_0_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001144(.in0(tmp00_2_9), .in1(tmp00_3_9), .out(tmp01_1_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001145(.in0(tmp00_4_9), .in1(tmp00_5_9), .out(tmp01_2_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001146(.in0(tmp00_6_9), .in1(tmp00_7_9), .out(tmp01_3_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001147(.in0(tmp00_8_9), .in1(tmp00_9_9), .out(tmp01_4_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001148(.in0(tmp00_10_9), .in1(tmp00_11_9), .out(tmp01_5_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001149(.in0(tmp00_12_9), .in1(tmp00_13_9), .out(tmp01_6_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001150(.in0(tmp00_14_9), .in1(tmp00_15_9), .out(tmp01_7_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001151(.in0(tmp00_16_9), .in1(tmp00_17_9), .out(tmp01_8_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001152(.in0(tmp00_18_9), .in1(tmp00_19_9), .out(tmp01_9_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001153(.in0(tmp00_20_9), .in1(tmp00_21_9), .out(tmp01_10_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001154(.in0(tmp00_22_9), .in1(tmp00_23_9), .out(tmp01_11_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001155(.in0(tmp00_24_9), .in1(tmp00_25_9), .out(tmp01_12_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001156(.in0(tmp00_26_9), .in1(tmp00_27_9), .out(tmp01_13_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001157(.in0(tmp00_28_9), .in1(tmp00_29_9), .out(tmp01_14_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001158(.in0(tmp00_30_9), .in1(tmp00_31_9), .out(tmp01_15_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001159(.in0(tmp00_32_9), .in1(tmp00_33_9), .out(tmp01_16_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001160(.in0(tmp00_34_9), .in1(tmp00_35_9), .out(tmp01_17_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001161(.in0(tmp00_36_9), .in1(tmp00_37_9), .out(tmp01_18_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001162(.in0(tmp00_38_9), .in1(tmp00_39_9), .out(tmp01_19_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001163(.in0(tmp00_40_9), .in1(tmp00_41_9), .out(tmp01_20_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001164(.in0(tmp00_42_9), .in1(tmp00_43_9), .out(tmp01_21_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001165(.in0(tmp00_44_9), .in1(tmp00_45_9), .out(tmp01_22_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001166(.in0(tmp00_46_9), .in1(tmp00_47_9), .out(tmp01_23_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001167(.in0(tmp00_48_9), .in1(tmp00_49_9), .out(tmp01_24_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001168(.in0(tmp00_50_9), .in1(tmp00_51_9), .out(tmp01_25_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001169(.in0(tmp00_52_9), .in1(tmp00_53_9), .out(tmp01_26_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001170(.in0(tmp00_54_9), .in1(tmp00_55_9), .out(tmp01_27_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001171(.in0(tmp00_56_9), .in1(tmp00_57_9), .out(tmp01_28_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001172(.in0(tmp00_58_9), .in1(tmp00_59_9), .out(tmp01_29_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001173(.in0(tmp00_60_9), .in1(tmp00_61_9), .out(tmp01_30_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001174(.in0(tmp00_62_9), .in1(tmp00_63_9), .out(tmp01_31_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001175(.in0(tmp00_64_9), .in1(tmp00_65_9), .out(tmp01_32_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001176(.in0(tmp00_66_9), .in1(tmp00_67_9), .out(tmp01_33_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001177(.in0(tmp00_68_9), .in1(tmp00_69_9), .out(tmp01_34_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001178(.in0(tmp00_70_9), .in1(tmp00_71_9), .out(tmp01_35_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001179(.in0(tmp00_72_9), .in1(tmp00_73_9), .out(tmp01_36_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001180(.in0(tmp00_74_9), .in1(tmp00_75_9), .out(tmp01_37_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001181(.in0(tmp00_76_9), .in1(tmp00_77_9), .out(tmp01_38_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001182(.in0(tmp00_78_9), .in1(tmp00_79_9), .out(tmp01_39_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001183(.in0(tmp00_80_9), .in1(tmp00_81_9), .out(tmp01_40_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001184(.in0(tmp00_82_9), .in1(tmp00_83_9), .out(tmp01_41_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001185(.in0(tmp00_84_9), .in1(tmp00_85_9), .out(tmp01_42_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001186(.in0(tmp00_86_9), .in1(tmp00_87_9), .out(tmp01_43_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001187(.in0(tmp00_88_9), .in1(tmp00_89_9), .out(tmp01_44_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001188(.in0(tmp00_90_9), .in1(tmp00_91_9), .out(tmp01_45_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001189(.in0(tmp00_92_9), .in1(tmp00_93_9), .out(tmp01_46_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001190(.in0(tmp00_94_9), .in1(tmp00_95_9), .out(tmp01_47_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001191(.in0(tmp00_96_9), .in1(tmp00_97_9), .out(tmp01_48_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001192(.in0(tmp00_98_9), .in1(tmp00_99_9), .out(tmp01_49_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001193(.in0(tmp00_100_9), .in1(tmp00_101_9), .out(tmp01_50_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001194(.in0(tmp00_102_9), .in1(tmp00_103_9), .out(tmp01_51_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001195(.in0(tmp00_104_9), .in1(tmp00_105_9), .out(tmp01_52_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001196(.in0(tmp00_106_9), .in1(tmp00_107_9), .out(tmp01_53_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001197(.in0(tmp00_108_9), .in1(tmp00_109_9), .out(tmp01_54_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001198(.in0(tmp00_110_9), .in1(tmp00_111_9), .out(tmp01_55_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001199(.in0(tmp00_112_9), .in1(tmp00_113_9), .out(tmp01_56_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001200(.in0(tmp00_114_9), .in1(tmp00_115_9), .out(tmp01_57_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001201(.in0(tmp00_116_9), .in1(tmp00_117_9), .out(tmp01_58_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001202(.in0(tmp00_118_9), .in1(tmp00_119_9), .out(tmp01_59_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001203(.in0(tmp00_120_9), .in1(tmp00_121_9), .out(tmp01_60_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001204(.in0(tmp00_122_9), .in1(tmp00_123_9), .out(tmp01_61_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001205(.in0(tmp00_124_9), .in1(tmp00_125_9), .out(tmp01_62_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001206(.in0(tmp00_126_9), .in1(tmp00_127_9), .out(tmp01_63_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001207(.in0(tmp01_0_9), .in1(tmp01_1_9), .out(tmp02_0_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001208(.in0(tmp01_2_9), .in1(tmp01_3_9), .out(tmp02_1_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001209(.in0(tmp01_4_9), .in1(tmp01_5_9), .out(tmp02_2_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001210(.in0(tmp01_6_9), .in1(tmp01_7_9), .out(tmp02_3_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001211(.in0(tmp01_8_9), .in1(tmp01_9_9), .out(tmp02_4_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001212(.in0(tmp01_10_9), .in1(tmp01_11_9), .out(tmp02_5_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001213(.in0(tmp01_12_9), .in1(tmp01_13_9), .out(tmp02_6_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001214(.in0(tmp01_14_9), .in1(tmp01_15_9), .out(tmp02_7_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001215(.in0(tmp01_16_9), .in1(tmp01_17_9), .out(tmp02_8_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001216(.in0(tmp01_18_9), .in1(tmp01_19_9), .out(tmp02_9_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001217(.in0(tmp01_20_9), .in1(tmp01_21_9), .out(tmp02_10_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001218(.in0(tmp01_22_9), .in1(tmp01_23_9), .out(tmp02_11_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001219(.in0(tmp01_24_9), .in1(tmp01_25_9), .out(tmp02_12_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001220(.in0(tmp01_26_9), .in1(tmp01_27_9), .out(tmp02_13_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001221(.in0(tmp01_28_9), .in1(tmp01_29_9), .out(tmp02_14_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001222(.in0(tmp01_30_9), .in1(tmp01_31_9), .out(tmp02_15_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001223(.in0(tmp01_32_9), .in1(tmp01_33_9), .out(tmp02_16_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001224(.in0(tmp01_34_9), .in1(tmp01_35_9), .out(tmp02_17_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001225(.in0(tmp01_36_9), .in1(tmp01_37_9), .out(tmp02_18_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001226(.in0(tmp01_38_9), .in1(tmp01_39_9), .out(tmp02_19_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001227(.in0(tmp01_40_9), .in1(tmp01_41_9), .out(tmp02_20_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001228(.in0(tmp01_42_9), .in1(tmp01_43_9), .out(tmp02_21_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001229(.in0(tmp01_44_9), .in1(tmp01_45_9), .out(tmp02_22_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001230(.in0(tmp01_46_9), .in1(tmp01_47_9), .out(tmp02_23_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001231(.in0(tmp01_48_9), .in1(tmp01_49_9), .out(tmp02_24_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001232(.in0(tmp01_50_9), .in1(tmp01_51_9), .out(tmp02_25_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001233(.in0(tmp01_52_9), .in1(tmp01_53_9), .out(tmp02_26_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001234(.in0(tmp01_54_9), .in1(tmp01_55_9), .out(tmp02_27_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001235(.in0(tmp01_56_9), .in1(tmp01_57_9), .out(tmp02_28_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001236(.in0(tmp01_58_9), .in1(tmp01_59_9), .out(tmp02_29_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001237(.in0(tmp01_60_9), .in1(tmp01_61_9), .out(tmp02_30_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001238(.in0(tmp01_62_9), .in1(tmp01_63_9), .out(tmp02_31_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001239(.in0(tmp02_0_9), .in1(tmp02_1_9), .out(tmp03_0_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001240(.in0(tmp02_2_9), .in1(tmp02_3_9), .out(tmp03_1_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001241(.in0(tmp02_4_9), .in1(tmp02_5_9), .out(tmp03_2_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001242(.in0(tmp02_6_9), .in1(tmp02_7_9), .out(tmp03_3_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001243(.in0(tmp02_8_9), .in1(tmp02_9_9), .out(tmp03_4_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001244(.in0(tmp02_10_9), .in1(tmp02_11_9), .out(tmp03_5_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001245(.in0(tmp02_12_9), .in1(tmp02_13_9), .out(tmp03_6_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001246(.in0(tmp02_14_9), .in1(tmp02_15_9), .out(tmp03_7_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001247(.in0(tmp02_16_9), .in1(tmp02_17_9), .out(tmp03_8_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001248(.in0(tmp02_18_9), .in1(tmp02_19_9), .out(tmp03_9_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001249(.in0(tmp02_20_9), .in1(tmp02_21_9), .out(tmp03_10_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001250(.in0(tmp02_22_9), .in1(tmp02_23_9), .out(tmp03_11_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001251(.in0(tmp02_24_9), .in1(tmp02_25_9), .out(tmp03_12_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001252(.in0(tmp02_26_9), .in1(tmp02_27_9), .out(tmp03_13_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001253(.in0(tmp02_28_9), .in1(tmp02_29_9), .out(tmp03_14_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001254(.in0(tmp02_30_9), .in1(tmp02_31_9), .out(tmp03_15_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001255(.in0(tmp03_0_9), .in1(tmp03_1_9), .out(tmp04_0_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001256(.in0(tmp03_2_9), .in1(tmp03_3_9), .out(tmp04_1_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001257(.in0(tmp03_4_9), .in1(tmp03_5_9), .out(tmp04_2_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001258(.in0(tmp03_6_9), .in1(tmp03_7_9), .out(tmp04_3_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001259(.in0(tmp03_8_9), .in1(tmp03_9_9), .out(tmp04_4_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001260(.in0(tmp03_10_9), .in1(tmp03_11_9), .out(tmp04_5_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001261(.in0(tmp03_12_9), .in1(tmp03_13_9), .out(tmp04_6_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001262(.in0(tmp03_14_9), .in1(tmp03_15_9), .out(tmp04_7_9));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001263(.in0(tmp04_0_9), .in1(tmp04_1_9), .out(tmp05_0_9));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001264(.in0(tmp04_2_9), .in1(tmp04_3_9), .out(tmp05_1_9));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001265(.in0(tmp04_4_9), .in1(tmp04_5_9), .out(tmp05_2_9));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001266(.in0(tmp04_6_9), .in1(tmp04_7_9), .out(tmp05_3_9));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001267(.in0(tmp05_0_9), .in1(tmp05_1_9), .out(tmp06_0_9));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001268(.in0(tmp05_2_9), .in1(tmp05_3_9), .out(tmp06_1_9));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add001269(.in0(tmp06_0_9), .in1(tmp06_1_9), .out(tmp07_0_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001270(.in0(tmp00_0_10), .in1(tmp00_1_10), .out(tmp01_0_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001271(.in0(tmp00_2_10), .in1(tmp00_3_10), .out(tmp01_1_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001272(.in0(tmp00_4_10), .in1(tmp00_5_10), .out(tmp01_2_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001273(.in0(tmp00_6_10), .in1(tmp00_7_10), .out(tmp01_3_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001274(.in0(tmp00_8_10), .in1(tmp00_9_10), .out(tmp01_4_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001275(.in0(tmp00_10_10), .in1(tmp00_11_10), .out(tmp01_5_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001276(.in0(tmp00_12_10), .in1(tmp00_13_10), .out(tmp01_6_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001277(.in0(tmp00_14_10), .in1(tmp00_15_10), .out(tmp01_7_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001278(.in0(tmp00_16_10), .in1(tmp00_17_10), .out(tmp01_8_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001279(.in0(tmp00_18_10), .in1(tmp00_19_10), .out(tmp01_9_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001280(.in0(tmp00_20_10), .in1(tmp00_21_10), .out(tmp01_10_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001281(.in0(tmp00_22_10), .in1(tmp00_23_10), .out(tmp01_11_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001282(.in0(tmp00_24_10), .in1(tmp00_25_10), .out(tmp01_12_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001283(.in0(tmp00_26_10), .in1(tmp00_27_10), .out(tmp01_13_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001284(.in0(tmp00_28_10), .in1(tmp00_29_10), .out(tmp01_14_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001285(.in0(tmp00_30_10), .in1(tmp00_31_10), .out(tmp01_15_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001286(.in0(tmp00_32_10), .in1(tmp00_33_10), .out(tmp01_16_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001287(.in0(tmp00_34_10), .in1(tmp00_35_10), .out(tmp01_17_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001288(.in0(tmp00_36_10), .in1(tmp00_37_10), .out(tmp01_18_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001289(.in0(tmp00_38_10), .in1(tmp00_39_10), .out(tmp01_19_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001290(.in0(tmp00_40_10), .in1(tmp00_41_10), .out(tmp01_20_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001291(.in0(tmp00_42_10), .in1(tmp00_43_10), .out(tmp01_21_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001292(.in0(tmp00_44_10), .in1(tmp00_45_10), .out(tmp01_22_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001293(.in0(tmp00_46_10), .in1(tmp00_47_10), .out(tmp01_23_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001294(.in0(tmp00_48_10), .in1(tmp00_49_10), .out(tmp01_24_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001295(.in0(tmp00_50_10), .in1(tmp00_51_10), .out(tmp01_25_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001296(.in0(tmp00_52_10), .in1(tmp00_53_10), .out(tmp01_26_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001297(.in0(tmp00_54_10), .in1(tmp00_55_10), .out(tmp01_27_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001298(.in0(tmp00_56_10), .in1(tmp00_57_10), .out(tmp01_28_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001299(.in0(tmp00_58_10), .in1(tmp00_59_10), .out(tmp01_29_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001300(.in0(tmp00_60_10), .in1(tmp00_61_10), .out(tmp01_30_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001301(.in0(tmp00_62_10), .in1(tmp00_63_10), .out(tmp01_31_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001302(.in0(tmp00_64_10), .in1(tmp00_65_10), .out(tmp01_32_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001303(.in0(tmp00_66_10), .in1(tmp00_67_10), .out(tmp01_33_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001304(.in0(tmp00_68_10), .in1(tmp00_69_10), .out(tmp01_34_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001305(.in0(tmp00_70_10), .in1(tmp00_71_10), .out(tmp01_35_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001306(.in0(tmp00_72_10), .in1(tmp00_73_10), .out(tmp01_36_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001307(.in0(tmp00_74_10), .in1(tmp00_75_10), .out(tmp01_37_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001308(.in0(tmp00_76_10), .in1(tmp00_77_10), .out(tmp01_38_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001309(.in0(tmp00_78_10), .in1(tmp00_79_10), .out(tmp01_39_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001310(.in0(tmp00_80_10), .in1(tmp00_81_10), .out(tmp01_40_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001311(.in0(tmp00_82_10), .in1(tmp00_83_10), .out(tmp01_41_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001312(.in0(tmp00_84_10), .in1(tmp00_85_10), .out(tmp01_42_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001313(.in0(tmp00_86_10), .in1(tmp00_87_10), .out(tmp01_43_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001314(.in0(tmp00_88_10), .in1(tmp00_89_10), .out(tmp01_44_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001315(.in0(tmp00_90_10), .in1(tmp00_91_10), .out(tmp01_45_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001316(.in0(tmp00_92_10), .in1(tmp00_93_10), .out(tmp01_46_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001317(.in0(tmp00_94_10), .in1(tmp00_95_10), .out(tmp01_47_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001318(.in0(tmp00_96_10), .in1(tmp00_97_10), .out(tmp01_48_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001319(.in0(tmp00_98_10), .in1(tmp00_99_10), .out(tmp01_49_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001320(.in0(tmp00_100_10), .in1(tmp00_101_10), .out(tmp01_50_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001321(.in0(tmp00_102_10), .in1(tmp00_103_10), .out(tmp01_51_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001322(.in0(tmp00_104_10), .in1(tmp00_105_10), .out(tmp01_52_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001323(.in0(tmp00_106_10), .in1(tmp00_107_10), .out(tmp01_53_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001324(.in0(tmp00_108_10), .in1(tmp00_109_10), .out(tmp01_54_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001325(.in0(tmp00_110_10), .in1(tmp00_111_10), .out(tmp01_55_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001326(.in0(tmp00_112_10), .in1(tmp00_113_10), .out(tmp01_56_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001327(.in0(tmp00_114_10), .in1(tmp00_115_10), .out(tmp01_57_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001328(.in0(tmp00_116_10), .in1(tmp00_117_10), .out(tmp01_58_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001329(.in0(tmp00_118_10), .in1(tmp00_119_10), .out(tmp01_59_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001330(.in0(tmp00_120_10), .in1(tmp00_121_10), .out(tmp01_60_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001331(.in0(tmp00_122_10), .in1(tmp00_123_10), .out(tmp01_61_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001332(.in0(tmp00_124_10), .in1(tmp00_125_10), .out(tmp01_62_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001333(.in0(tmp00_126_10), .in1(tmp00_127_10), .out(tmp01_63_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001334(.in0(tmp01_0_10), .in1(tmp01_1_10), .out(tmp02_0_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001335(.in0(tmp01_2_10), .in1(tmp01_3_10), .out(tmp02_1_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001336(.in0(tmp01_4_10), .in1(tmp01_5_10), .out(tmp02_2_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001337(.in0(tmp01_6_10), .in1(tmp01_7_10), .out(tmp02_3_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001338(.in0(tmp01_8_10), .in1(tmp01_9_10), .out(tmp02_4_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001339(.in0(tmp01_10_10), .in1(tmp01_11_10), .out(tmp02_5_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001340(.in0(tmp01_12_10), .in1(tmp01_13_10), .out(tmp02_6_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001341(.in0(tmp01_14_10), .in1(tmp01_15_10), .out(tmp02_7_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001342(.in0(tmp01_16_10), .in1(tmp01_17_10), .out(tmp02_8_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001343(.in0(tmp01_18_10), .in1(tmp01_19_10), .out(tmp02_9_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001344(.in0(tmp01_20_10), .in1(tmp01_21_10), .out(tmp02_10_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001345(.in0(tmp01_22_10), .in1(tmp01_23_10), .out(tmp02_11_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001346(.in0(tmp01_24_10), .in1(tmp01_25_10), .out(tmp02_12_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001347(.in0(tmp01_26_10), .in1(tmp01_27_10), .out(tmp02_13_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001348(.in0(tmp01_28_10), .in1(tmp01_29_10), .out(tmp02_14_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001349(.in0(tmp01_30_10), .in1(tmp01_31_10), .out(tmp02_15_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001350(.in0(tmp01_32_10), .in1(tmp01_33_10), .out(tmp02_16_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001351(.in0(tmp01_34_10), .in1(tmp01_35_10), .out(tmp02_17_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001352(.in0(tmp01_36_10), .in1(tmp01_37_10), .out(tmp02_18_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001353(.in0(tmp01_38_10), .in1(tmp01_39_10), .out(tmp02_19_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001354(.in0(tmp01_40_10), .in1(tmp01_41_10), .out(tmp02_20_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001355(.in0(tmp01_42_10), .in1(tmp01_43_10), .out(tmp02_21_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001356(.in0(tmp01_44_10), .in1(tmp01_45_10), .out(tmp02_22_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001357(.in0(tmp01_46_10), .in1(tmp01_47_10), .out(tmp02_23_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001358(.in0(tmp01_48_10), .in1(tmp01_49_10), .out(tmp02_24_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001359(.in0(tmp01_50_10), .in1(tmp01_51_10), .out(tmp02_25_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001360(.in0(tmp01_52_10), .in1(tmp01_53_10), .out(tmp02_26_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001361(.in0(tmp01_54_10), .in1(tmp01_55_10), .out(tmp02_27_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001362(.in0(tmp01_56_10), .in1(tmp01_57_10), .out(tmp02_28_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001363(.in0(tmp01_58_10), .in1(tmp01_59_10), .out(tmp02_29_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001364(.in0(tmp01_60_10), .in1(tmp01_61_10), .out(tmp02_30_10));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001365(.in0(tmp01_62_10), .in1(tmp01_63_10), .out(tmp02_31_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001366(.in0(tmp02_0_10), .in1(tmp02_1_10), .out(tmp03_0_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001367(.in0(tmp02_2_10), .in1(tmp02_3_10), .out(tmp03_1_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001368(.in0(tmp02_4_10), .in1(tmp02_5_10), .out(tmp03_2_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001369(.in0(tmp02_6_10), .in1(tmp02_7_10), .out(tmp03_3_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001370(.in0(tmp02_8_10), .in1(tmp02_9_10), .out(tmp03_4_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001371(.in0(tmp02_10_10), .in1(tmp02_11_10), .out(tmp03_5_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001372(.in0(tmp02_12_10), .in1(tmp02_13_10), .out(tmp03_6_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001373(.in0(tmp02_14_10), .in1(tmp02_15_10), .out(tmp03_7_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001374(.in0(tmp02_16_10), .in1(tmp02_17_10), .out(tmp03_8_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001375(.in0(tmp02_18_10), .in1(tmp02_19_10), .out(tmp03_9_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001376(.in0(tmp02_20_10), .in1(tmp02_21_10), .out(tmp03_10_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001377(.in0(tmp02_22_10), .in1(tmp02_23_10), .out(tmp03_11_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001378(.in0(tmp02_24_10), .in1(tmp02_25_10), .out(tmp03_12_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001379(.in0(tmp02_26_10), .in1(tmp02_27_10), .out(tmp03_13_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001380(.in0(tmp02_28_10), .in1(tmp02_29_10), .out(tmp03_14_10));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001381(.in0(tmp02_30_10), .in1(tmp02_31_10), .out(tmp03_15_10));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001382(.in0(tmp03_0_10), .in1(tmp03_1_10), .out(tmp04_0_10));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001383(.in0(tmp03_2_10), .in1(tmp03_3_10), .out(tmp04_1_10));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001384(.in0(tmp03_4_10), .in1(tmp03_5_10), .out(tmp04_2_10));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001385(.in0(tmp03_6_10), .in1(tmp03_7_10), .out(tmp04_3_10));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001386(.in0(tmp03_8_10), .in1(tmp03_9_10), .out(tmp04_4_10));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001387(.in0(tmp03_10_10), .in1(tmp03_11_10), .out(tmp04_5_10));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001388(.in0(tmp03_12_10), .in1(tmp03_13_10), .out(tmp04_6_10));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001389(.in0(tmp03_14_10), .in1(tmp03_15_10), .out(tmp04_7_10));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001390(.in0(tmp04_0_10), .in1(tmp04_1_10), .out(tmp05_0_10));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001391(.in0(tmp04_2_10), .in1(tmp04_3_10), .out(tmp05_1_10));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001392(.in0(tmp04_4_10), .in1(tmp04_5_10), .out(tmp05_2_10));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001393(.in0(tmp04_6_10), .in1(tmp04_7_10), .out(tmp05_3_10));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001394(.in0(tmp05_0_10), .in1(tmp05_1_10), .out(tmp06_0_10));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001395(.in0(tmp05_2_10), .in1(tmp05_3_10), .out(tmp06_1_10));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add001396(.in0(tmp06_0_10), .in1(tmp06_1_10), .out(tmp07_0_10));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001397(.in0(tmp00_0_11), .in1(tmp00_1_11), .out(tmp01_0_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001398(.in0(tmp00_2_11), .in1(tmp00_3_11), .out(tmp01_1_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001399(.in0(tmp00_4_11), .in1(tmp00_5_11), .out(tmp01_2_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001400(.in0(tmp00_6_11), .in1(tmp00_7_11), .out(tmp01_3_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001401(.in0(tmp00_8_11), .in1(tmp00_9_11), .out(tmp01_4_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001402(.in0(tmp00_10_11), .in1(tmp00_11_11), .out(tmp01_5_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001403(.in0(tmp00_12_11), .in1(tmp00_13_11), .out(tmp01_6_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001404(.in0(tmp00_14_11), .in1(tmp00_15_11), .out(tmp01_7_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001405(.in0(tmp00_16_11), .in1(tmp00_17_11), .out(tmp01_8_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001406(.in0(tmp00_18_11), .in1(tmp00_19_11), .out(tmp01_9_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001407(.in0(tmp00_20_11), .in1(tmp00_21_11), .out(tmp01_10_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001408(.in0(tmp00_22_11), .in1(tmp00_23_11), .out(tmp01_11_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001409(.in0(tmp00_24_11), .in1(tmp00_25_11), .out(tmp01_12_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001410(.in0(tmp00_26_11), .in1(tmp00_27_11), .out(tmp01_13_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001411(.in0(tmp00_28_11), .in1(tmp00_29_11), .out(tmp01_14_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001412(.in0(tmp00_30_11), .in1(tmp00_31_11), .out(tmp01_15_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001413(.in0(tmp00_32_11), .in1(tmp00_33_11), .out(tmp01_16_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001414(.in0(tmp00_34_11), .in1(tmp00_35_11), .out(tmp01_17_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001415(.in0(tmp00_36_11), .in1(tmp00_37_11), .out(tmp01_18_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001416(.in0(tmp00_38_11), .in1(tmp00_39_11), .out(tmp01_19_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001417(.in0(tmp00_40_11), .in1(tmp00_41_11), .out(tmp01_20_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001418(.in0(tmp00_42_11), .in1(tmp00_43_11), .out(tmp01_21_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001419(.in0(tmp00_44_11), .in1(tmp00_45_11), .out(tmp01_22_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001420(.in0(tmp00_46_11), .in1(tmp00_47_11), .out(tmp01_23_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001421(.in0(tmp00_48_11), .in1(tmp00_49_11), .out(tmp01_24_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001422(.in0(tmp00_50_11), .in1(tmp00_51_11), .out(tmp01_25_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001423(.in0(tmp00_52_11), .in1(tmp00_53_11), .out(tmp01_26_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001424(.in0(tmp00_54_11), .in1(tmp00_55_11), .out(tmp01_27_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001425(.in0(tmp00_56_11), .in1(tmp00_57_11), .out(tmp01_28_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001426(.in0(tmp00_58_11), .in1(tmp00_59_11), .out(tmp01_29_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001427(.in0(tmp00_60_11), .in1(tmp00_61_11), .out(tmp01_30_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001428(.in0(tmp00_62_11), .in1(tmp00_63_11), .out(tmp01_31_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001429(.in0(tmp00_64_11), .in1(tmp00_65_11), .out(tmp01_32_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001430(.in0(tmp00_66_11), .in1(tmp00_67_11), .out(tmp01_33_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001431(.in0(tmp00_68_11), .in1(tmp00_69_11), .out(tmp01_34_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001432(.in0(tmp00_70_11), .in1(tmp00_71_11), .out(tmp01_35_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001433(.in0(tmp00_72_11), .in1(tmp00_73_11), .out(tmp01_36_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001434(.in0(tmp00_74_11), .in1(tmp00_75_11), .out(tmp01_37_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001435(.in0(tmp00_76_11), .in1(tmp00_77_11), .out(tmp01_38_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001436(.in0(tmp00_78_11), .in1(tmp00_79_11), .out(tmp01_39_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001437(.in0(tmp00_80_11), .in1(tmp00_81_11), .out(tmp01_40_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001438(.in0(tmp00_82_11), .in1(tmp00_83_11), .out(tmp01_41_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001439(.in0(tmp00_84_11), .in1(tmp00_85_11), .out(tmp01_42_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001440(.in0(tmp00_86_11), .in1(tmp00_87_11), .out(tmp01_43_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001441(.in0(tmp00_88_11), .in1(tmp00_89_11), .out(tmp01_44_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001442(.in0(tmp00_90_11), .in1(tmp00_91_11), .out(tmp01_45_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001443(.in0(tmp00_92_11), .in1(tmp00_93_11), .out(tmp01_46_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001444(.in0(tmp00_94_11), .in1(tmp00_95_11), .out(tmp01_47_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001445(.in0(tmp00_96_11), .in1(tmp00_97_11), .out(tmp01_48_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001446(.in0(tmp00_98_11), .in1(tmp00_99_11), .out(tmp01_49_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001447(.in0(tmp00_100_11), .in1(tmp00_101_11), .out(tmp01_50_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001448(.in0(tmp00_102_11), .in1(tmp00_103_11), .out(tmp01_51_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001449(.in0(tmp00_104_11), .in1(tmp00_105_11), .out(tmp01_52_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001450(.in0(tmp00_106_11), .in1(tmp00_107_11), .out(tmp01_53_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001451(.in0(tmp00_108_11), .in1(tmp00_109_11), .out(tmp01_54_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001452(.in0(tmp00_110_11), .in1(tmp00_111_11), .out(tmp01_55_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001453(.in0(tmp00_112_11), .in1(tmp00_113_11), .out(tmp01_56_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001454(.in0(tmp00_114_11), .in1(tmp00_115_11), .out(tmp01_57_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001455(.in0(tmp00_116_11), .in1(tmp00_117_11), .out(tmp01_58_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001456(.in0(tmp00_118_11), .in1(tmp00_119_11), .out(tmp01_59_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001457(.in0(tmp00_120_11), .in1(tmp00_121_11), .out(tmp01_60_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001458(.in0(tmp00_122_11), .in1(tmp00_123_11), .out(tmp01_61_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001459(.in0(tmp00_124_11), .in1(tmp00_125_11), .out(tmp01_62_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001460(.in0(tmp00_126_11), .in1(tmp00_127_11), .out(tmp01_63_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001461(.in0(tmp01_0_11), .in1(tmp01_1_11), .out(tmp02_0_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001462(.in0(tmp01_2_11), .in1(tmp01_3_11), .out(tmp02_1_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001463(.in0(tmp01_4_11), .in1(tmp01_5_11), .out(tmp02_2_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001464(.in0(tmp01_6_11), .in1(tmp01_7_11), .out(tmp02_3_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001465(.in0(tmp01_8_11), .in1(tmp01_9_11), .out(tmp02_4_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001466(.in0(tmp01_10_11), .in1(tmp01_11_11), .out(tmp02_5_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001467(.in0(tmp01_12_11), .in1(tmp01_13_11), .out(tmp02_6_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001468(.in0(tmp01_14_11), .in1(tmp01_15_11), .out(tmp02_7_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001469(.in0(tmp01_16_11), .in1(tmp01_17_11), .out(tmp02_8_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001470(.in0(tmp01_18_11), .in1(tmp01_19_11), .out(tmp02_9_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001471(.in0(tmp01_20_11), .in1(tmp01_21_11), .out(tmp02_10_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001472(.in0(tmp01_22_11), .in1(tmp01_23_11), .out(tmp02_11_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001473(.in0(tmp01_24_11), .in1(tmp01_25_11), .out(tmp02_12_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001474(.in0(tmp01_26_11), .in1(tmp01_27_11), .out(tmp02_13_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001475(.in0(tmp01_28_11), .in1(tmp01_29_11), .out(tmp02_14_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001476(.in0(tmp01_30_11), .in1(tmp01_31_11), .out(tmp02_15_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001477(.in0(tmp01_32_11), .in1(tmp01_33_11), .out(tmp02_16_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001478(.in0(tmp01_34_11), .in1(tmp01_35_11), .out(tmp02_17_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001479(.in0(tmp01_36_11), .in1(tmp01_37_11), .out(tmp02_18_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001480(.in0(tmp01_38_11), .in1(tmp01_39_11), .out(tmp02_19_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001481(.in0(tmp01_40_11), .in1(tmp01_41_11), .out(tmp02_20_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001482(.in0(tmp01_42_11), .in1(tmp01_43_11), .out(tmp02_21_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001483(.in0(tmp01_44_11), .in1(tmp01_45_11), .out(tmp02_22_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001484(.in0(tmp01_46_11), .in1(tmp01_47_11), .out(tmp02_23_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001485(.in0(tmp01_48_11), .in1(tmp01_49_11), .out(tmp02_24_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001486(.in0(tmp01_50_11), .in1(tmp01_51_11), .out(tmp02_25_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001487(.in0(tmp01_52_11), .in1(tmp01_53_11), .out(tmp02_26_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001488(.in0(tmp01_54_11), .in1(tmp01_55_11), .out(tmp02_27_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001489(.in0(tmp01_56_11), .in1(tmp01_57_11), .out(tmp02_28_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001490(.in0(tmp01_58_11), .in1(tmp01_59_11), .out(tmp02_29_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001491(.in0(tmp01_60_11), .in1(tmp01_61_11), .out(tmp02_30_11));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001492(.in0(tmp01_62_11), .in1(tmp01_63_11), .out(tmp02_31_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001493(.in0(tmp02_0_11), .in1(tmp02_1_11), .out(tmp03_0_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001494(.in0(tmp02_2_11), .in1(tmp02_3_11), .out(tmp03_1_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001495(.in0(tmp02_4_11), .in1(tmp02_5_11), .out(tmp03_2_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001496(.in0(tmp02_6_11), .in1(tmp02_7_11), .out(tmp03_3_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001497(.in0(tmp02_8_11), .in1(tmp02_9_11), .out(tmp03_4_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001498(.in0(tmp02_10_11), .in1(tmp02_11_11), .out(tmp03_5_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001499(.in0(tmp02_12_11), .in1(tmp02_13_11), .out(tmp03_6_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001500(.in0(tmp02_14_11), .in1(tmp02_15_11), .out(tmp03_7_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001501(.in0(tmp02_16_11), .in1(tmp02_17_11), .out(tmp03_8_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001502(.in0(tmp02_18_11), .in1(tmp02_19_11), .out(tmp03_9_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001503(.in0(tmp02_20_11), .in1(tmp02_21_11), .out(tmp03_10_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001504(.in0(tmp02_22_11), .in1(tmp02_23_11), .out(tmp03_11_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001505(.in0(tmp02_24_11), .in1(tmp02_25_11), .out(tmp03_12_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001506(.in0(tmp02_26_11), .in1(tmp02_27_11), .out(tmp03_13_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001507(.in0(tmp02_28_11), .in1(tmp02_29_11), .out(tmp03_14_11));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001508(.in0(tmp02_30_11), .in1(tmp02_31_11), .out(tmp03_15_11));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001509(.in0(tmp03_0_11), .in1(tmp03_1_11), .out(tmp04_0_11));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001510(.in0(tmp03_2_11), .in1(tmp03_3_11), .out(tmp04_1_11));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001511(.in0(tmp03_4_11), .in1(tmp03_5_11), .out(tmp04_2_11));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001512(.in0(tmp03_6_11), .in1(tmp03_7_11), .out(tmp04_3_11));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001513(.in0(tmp03_8_11), .in1(tmp03_9_11), .out(tmp04_4_11));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001514(.in0(tmp03_10_11), .in1(tmp03_11_11), .out(tmp04_5_11));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001515(.in0(tmp03_12_11), .in1(tmp03_13_11), .out(tmp04_6_11));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001516(.in0(tmp03_14_11), .in1(tmp03_15_11), .out(tmp04_7_11));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001517(.in0(tmp04_0_11), .in1(tmp04_1_11), .out(tmp05_0_11));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001518(.in0(tmp04_2_11), .in1(tmp04_3_11), .out(tmp05_1_11));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001519(.in0(tmp04_4_11), .in1(tmp04_5_11), .out(tmp05_2_11));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001520(.in0(tmp04_6_11), .in1(tmp04_7_11), .out(tmp05_3_11));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001521(.in0(tmp05_0_11), .in1(tmp05_1_11), .out(tmp06_0_11));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001522(.in0(tmp05_2_11), .in1(tmp05_3_11), .out(tmp06_1_11));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add001523(.in0(tmp06_0_11), .in1(tmp06_1_11), .out(tmp07_0_11));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001524(.in0(tmp00_0_12), .in1(tmp00_1_12), .out(tmp01_0_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001525(.in0(tmp00_2_12), .in1(tmp00_3_12), .out(tmp01_1_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001526(.in0(tmp00_4_12), .in1(tmp00_5_12), .out(tmp01_2_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001527(.in0(tmp00_6_12), .in1(tmp00_7_12), .out(tmp01_3_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001528(.in0(tmp00_8_12), .in1(tmp00_9_12), .out(tmp01_4_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001529(.in0(tmp00_10_12), .in1(tmp00_11_12), .out(tmp01_5_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001530(.in0(tmp00_12_12), .in1(tmp00_13_12), .out(tmp01_6_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001531(.in0(tmp00_14_12), .in1(tmp00_15_12), .out(tmp01_7_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001532(.in0(tmp00_16_12), .in1(tmp00_17_12), .out(tmp01_8_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001533(.in0(tmp00_18_12), .in1(tmp00_19_12), .out(tmp01_9_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001534(.in0(tmp00_20_12), .in1(tmp00_21_12), .out(tmp01_10_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001535(.in0(tmp00_22_12), .in1(tmp00_23_12), .out(tmp01_11_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001536(.in0(tmp00_24_12), .in1(tmp00_25_12), .out(tmp01_12_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001537(.in0(tmp00_26_12), .in1(tmp00_27_12), .out(tmp01_13_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001538(.in0(tmp00_28_12), .in1(tmp00_29_12), .out(tmp01_14_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001539(.in0(tmp00_30_12), .in1(tmp00_31_12), .out(tmp01_15_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001540(.in0(tmp00_32_12), .in1(tmp00_33_12), .out(tmp01_16_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001541(.in0(tmp00_34_12), .in1(tmp00_35_12), .out(tmp01_17_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001542(.in0(tmp00_36_12), .in1(tmp00_37_12), .out(tmp01_18_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001543(.in0(tmp00_38_12), .in1(tmp00_39_12), .out(tmp01_19_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001544(.in0(tmp00_40_12), .in1(tmp00_41_12), .out(tmp01_20_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001545(.in0(tmp00_42_12), .in1(tmp00_43_12), .out(tmp01_21_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001546(.in0(tmp00_44_12), .in1(tmp00_45_12), .out(tmp01_22_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001547(.in0(tmp00_46_12), .in1(tmp00_47_12), .out(tmp01_23_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001548(.in0(tmp00_48_12), .in1(tmp00_49_12), .out(tmp01_24_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001549(.in0(tmp00_50_12), .in1(tmp00_51_12), .out(tmp01_25_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001550(.in0(tmp00_52_12), .in1(tmp00_53_12), .out(tmp01_26_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001551(.in0(tmp00_54_12), .in1(tmp00_55_12), .out(tmp01_27_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001552(.in0(tmp00_56_12), .in1(tmp00_57_12), .out(tmp01_28_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001553(.in0(tmp00_58_12), .in1(tmp00_59_12), .out(tmp01_29_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001554(.in0(tmp00_60_12), .in1(tmp00_61_12), .out(tmp01_30_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001555(.in0(tmp00_62_12), .in1(tmp00_63_12), .out(tmp01_31_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001556(.in0(tmp00_64_12), .in1(tmp00_65_12), .out(tmp01_32_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001557(.in0(tmp00_66_12), .in1(tmp00_67_12), .out(tmp01_33_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001558(.in0(tmp00_68_12), .in1(tmp00_69_12), .out(tmp01_34_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001559(.in0(tmp00_70_12), .in1(tmp00_71_12), .out(tmp01_35_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001560(.in0(tmp00_72_12), .in1(tmp00_73_12), .out(tmp01_36_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001561(.in0(tmp00_74_12), .in1(tmp00_75_12), .out(tmp01_37_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001562(.in0(tmp00_76_12), .in1(tmp00_77_12), .out(tmp01_38_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001563(.in0(tmp00_78_12), .in1(tmp00_79_12), .out(tmp01_39_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001564(.in0(tmp00_80_12), .in1(tmp00_81_12), .out(tmp01_40_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001565(.in0(tmp00_82_12), .in1(tmp00_83_12), .out(tmp01_41_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001566(.in0(tmp00_84_12), .in1(tmp00_85_12), .out(tmp01_42_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001567(.in0(tmp00_86_12), .in1(tmp00_87_12), .out(tmp01_43_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001568(.in0(tmp00_88_12), .in1(tmp00_89_12), .out(tmp01_44_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001569(.in0(tmp00_90_12), .in1(tmp00_91_12), .out(tmp01_45_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001570(.in0(tmp00_92_12), .in1(tmp00_93_12), .out(tmp01_46_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001571(.in0(tmp00_94_12), .in1(tmp00_95_12), .out(tmp01_47_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001572(.in0(tmp00_96_12), .in1(tmp00_97_12), .out(tmp01_48_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001573(.in0(tmp00_98_12), .in1(tmp00_99_12), .out(tmp01_49_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001574(.in0(tmp00_100_12), .in1(tmp00_101_12), .out(tmp01_50_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001575(.in0(tmp00_102_12), .in1(tmp00_103_12), .out(tmp01_51_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001576(.in0(tmp00_104_12), .in1(tmp00_105_12), .out(tmp01_52_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001577(.in0(tmp00_106_12), .in1(tmp00_107_12), .out(tmp01_53_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001578(.in0(tmp00_108_12), .in1(tmp00_109_12), .out(tmp01_54_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001579(.in0(tmp00_110_12), .in1(tmp00_111_12), .out(tmp01_55_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001580(.in0(tmp00_112_12), .in1(tmp00_113_12), .out(tmp01_56_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001581(.in0(tmp00_114_12), .in1(tmp00_115_12), .out(tmp01_57_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001582(.in0(tmp00_116_12), .in1(tmp00_117_12), .out(tmp01_58_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001583(.in0(tmp00_118_12), .in1(tmp00_119_12), .out(tmp01_59_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001584(.in0(tmp00_120_12), .in1(tmp00_121_12), .out(tmp01_60_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001585(.in0(tmp00_122_12), .in1(tmp00_123_12), .out(tmp01_61_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001586(.in0(tmp00_124_12), .in1(tmp00_125_12), .out(tmp01_62_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001587(.in0(tmp00_126_12), .in1(tmp00_127_12), .out(tmp01_63_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001588(.in0(tmp01_0_12), .in1(tmp01_1_12), .out(tmp02_0_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001589(.in0(tmp01_2_12), .in1(tmp01_3_12), .out(tmp02_1_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001590(.in0(tmp01_4_12), .in1(tmp01_5_12), .out(tmp02_2_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001591(.in0(tmp01_6_12), .in1(tmp01_7_12), .out(tmp02_3_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001592(.in0(tmp01_8_12), .in1(tmp01_9_12), .out(tmp02_4_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001593(.in0(tmp01_10_12), .in1(tmp01_11_12), .out(tmp02_5_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001594(.in0(tmp01_12_12), .in1(tmp01_13_12), .out(tmp02_6_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001595(.in0(tmp01_14_12), .in1(tmp01_15_12), .out(tmp02_7_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001596(.in0(tmp01_16_12), .in1(tmp01_17_12), .out(tmp02_8_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001597(.in0(tmp01_18_12), .in1(tmp01_19_12), .out(tmp02_9_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001598(.in0(tmp01_20_12), .in1(tmp01_21_12), .out(tmp02_10_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001599(.in0(tmp01_22_12), .in1(tmp01_23_12), .out(tmp02_11_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001600(.in0(tmp01_24_12), .in1(tmp01_25_12), .out(tmp02_12_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001601(.in0(tmp01_26_12), .in1(tmp01_27_12), .out(tmp02_13_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001602(.in0(tmp01_28_12), .in1(tmp01_29_12), .out(tmp02_14_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001603(.in0(tmp01_30_12), .in1(tmp01_31_12), .out(tmp02_15_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001604(.in0(tmp01_32_12), .in1(tmp01_33_12), .out(tmp02_16_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001605(.in0(tmp01_34_12), .in1(tmp01_35_12), .out(tmp02_17_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001606(.in0(tmp01_36_12), .in1(tmp01_37_12), .out(tmp02_18_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001607(.in0(tmp01_38_12), .in1(tmp01_39_12), .out(tmp02_19_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001608(.in0(tmp01_40_12), .in1(tmp01_41_12), .out(tmp02_20_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001609(.in0(tmp01_42_12), .in1(tmp01_43_12), .out(tmp02_21_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001610(.in0(tmp01_44_12), .in1(tmp01_45_12), .out(tmp02_22_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001611(.in0(tmp01_46_12), .in1(tmp01_47_12), .out(tmp02_23_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001612(.in0(tmp01_48_12), .in1(tmp01_49_12), .out(tmp02_24_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001613(.in0(tmp01_50_12), .in1(tmp01_51_12), .out(tmp02_25_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001614(.in0(tmp01_52_12), .in1(tmp01_53_12), .out(tmp02_26_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001615(.in0(tmp01_54_12), .in1(tmp01_55_12), .out(tmp02_27_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001616(.in0(tmp01_56_12), .in1(tmp01_57_12), .out(tmp02_28_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001617(.in0(tmp01_58_12), .in1(tmp01_59_12), .out(tmp02_29_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001618(.in0(tmp01_60_12), .in1(tmp01_61_12), .out(tmp02_30_12));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001619(.in0(tmp01_62_12), .in1(tmp01_63_12), .out(tmp02_31_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001620(.in0(tmp02_0_12), .in1(tmp02_1_12), .out(tmp03_0_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001621(.in0(tmp02_2_12), .in1(tmp02_3_12), .out(tmp03_1_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001622(.in0(tmp02_4_12), .in1(tmp02_5_12), .out(tmp03_2_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001623(.in0(tmp02_6_12), .in1(tmp02_7_12), .out(tmp03_3_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001624(.in0(tmp02_8_12), .in1(tmp02_9_12), .out(tmp03_4_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001625(.in0(tmp02_10_12), .in1(tmp02_11_12), .out(tmp03_5_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001626(.in0(tmp02_12_12), .in1(tmp02_13_12), .out(tmp03_6_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001627(.in0(tmp02_14_12), .in1(tmp02_15_12), .out(tmp03_7_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001628(.in0(tmp02_16_12), .in1(tmp02_17_12), .out(tmp03_8_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001629(.in0(tmp02_18_12), .in1(tmp02_19_12), .out(tmp03_9_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001630(.in0(tmp02_20_12), .in1(tmp02_21_12), .out(tmp03_10_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001631(.in0(tmp02_22_12), .in1(tmp02_23_12), .out(tmp03_11_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001632(.in0(tmp02_24_12), .in1(tmp02_25_12), .out(tmp03_12_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001633(.in0(tmp02_26_12), .in1(tmp02_27_12), .out(tmp03_13_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001634(.in0(tmp02_28_12), .in1(tmp02_29_12), .out(tmp03_14_12));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001635(.in0(tmp02_30_12), .in1(tmp02_31_12), .out(tmp03_15_12));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001636(.in0(tmp03_0_12), .in1(tmp03_1_12), .out(tmp04_0_12));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001637(.in0(tmp03_2_12), .in1(tmp03_3_12), .out(tmp04_1_12));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001638(.in0(tmp03_4_12), .in1(tmp03_5_12), .out(tmp04_2_12));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001639(.in0(tmp03_6_12), .in1(tmp03_7_12), .out(tmp04_3_12));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001640(.in0(tmp03_8_12), .in1(tmp03_9_12), .out(tmp04_4_12));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001641(.in0(tmp03_10_12), .in1(tmp03_11_12), .out(tmp04_5_12));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001642(.in0(tmp03_12_12), .in1(tmp03_13_12), .out(tmp04_6_12));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001643(.in0(tmp03_14_12), .in1(tmp03_15_12), .out(tmp04_7_12));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001644(.in0(tmp04_0_12), .in1(tmp04_1_12), .out(tmp05_0_12));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001645(.in0(tmp04_2_12), .in1(tmp04_3_12), .out(tmp05_1_12));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001646(.in0(tmp04_4_12), .in1(tmp04_5_12), .out(tmp05_2_12));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001647(.in0(tmp04_6_12), .in1(tmp04_7_12), .out(tmp05_3_12));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001648(.in0(tmp05_0_12), .in1(tmp05_1_12), .out(tmp06_0_12));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001649(.in0(tmp05_2_12), .in1(tmp05_3_12), .out(tmp06_1_12));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add001650(.in0(tmp06_0_12), .in1(tmp06_1_12), .out(tmp07_0_12));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001651(.in0(tmp00_0_13), .in1(tmp00_1_13), .out(tmp01_0_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001652(.in0(tmp00_2_13), .in1(tmp00_3_13), .out(tmp01_1_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001653(.in0(tmp00_4_13), .in1(tmp00_5_13), .out(tmp01_2_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001654(.in0(tmp00_6_13), .in1(tmp00_7_13), .out(tmp01_3_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001655(.in0(tmp00_8_13), .in1(tmp00_9_13), .out(tmp01_4_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001656(.in0(tmp00_10_13), .in1(tmp00_11_13), .out(tmp01_5_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001657(.in0(tmp00_12_13), .in1(tmp00_13_13), .out(tmp01_6_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001658(.in0(tmp00_14_13), .in1(tmp00_15_13), .out(tmp01_7_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001659(.in0(tmp00_16_13), .in1(tmp00_17_13), .out(tmp01_8_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001660(.in0(tmp00_18_13), .in1(tmp00_19_13), .out(tmp01_9_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001661(.in0(tmp00_20_13), .in1(tmp00_21_13), .out(tmp01_10_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001662(.in0(tmp00_22_13), .in1(tmp00_23_13), .out(tmp01_11_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001663(.in0(tmp00_24_13), .in1(tmp00_25_13), .out(tmp01_12_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001664(.in0(tmp00_26_13), .in1(tmp00_27_13), .out(tmp01_13_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001665(.in0(tmp00_28_13), .in1(tmp00_29_13), .out(tmp01_14_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001666(.in0(tmp00_30_13), .in1(tmp00_31_13), .out(tmp01_15_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001667(.in0(tmp00_32_13), .in1(tmp00_33_13), .out(tmp01_16_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001668(.in0(tmp00_34_13), .in1(tmp00_35_13), .out(tmp01_17_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001669(.in0(tmp00_36_13), .in1(tmp00_37_13), .out(tmp01_18_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001670(.in0(tmp00_38_13), .in1(tmp00_39_13), .out(tmp01_19_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001671(.in0(tmp00_40_13), .in1(tmp00_41_13), .out(tmp01_20_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001672(.in0(tmp00_42_13), .in1(tmp00_43_13), .out(tmp01_21_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001673(.in0(tmp00_44_13), .in1(tmp00_45_13), .out(tmp01_22_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001674(.in0(tmp00_46_13), .in1(tmp00_47_13), .out(tmp01_23_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001675(.in0(tmp00_48_13), .in1(tmp00_49_13), .out(tmp01_24_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001676(.in0(tmp00_50_13), .in1(tmp00_51_13), .out(tmp01_25_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001677(.in0(tmp00_52_13), .in1(tmp00_53_13), .out(tmp01_26_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001678(.in0(tmp00_54_13), .in1(tmp00_55_13), .out(tmp01_27_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001679(.in0(tmp00_56_13), .in1(tmp00_57_13), .out(tmp01_28_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001680(.in0(tmp00_58_13), .in1(tmp00_59_13), .out(tmp01_29_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001681(.in0(tmp00_60_13), .in1(tmp00_61_13), .out(tmp01_30_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001682(.in0(tmp00_62_13), .in1(tmp00_63_13), .out(tmp01_31_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001683(.in0(tmp00_64_13), .in1(tmp00_65_13), .out(tmp01_32_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001684(.in0(tmp00_66_13), .in1(tmp00_67_13), .out(tmp01_33_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001685(.in0(tmp00_68_13), .in1(tmp00_69_13), .out(tmp01_34_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001686(.in0(tmp00_70_13), .in1(tmp00_71_13), .out(tmp01_35_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001687(.in0(tmp00_72_13), .in1(tmp00_73_13), .out(tmp01_36_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001688(.in0(tmp00_74_13), .in1(tmp00_75_13), .out(tmp01_37_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001689(.in0(tmp00_76_13), .in1(tmp00_77_13), .out(tmp01_38_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001690(.in0(tmp00_78_13), .in1(tmp00_79_13), .out(tmp01_39_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001691(.in0(tmp00_80_13), .in1(tmp00_81_13), .out(tmp01_40_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001692(.in0(tmp00_82_13), .in1(tmp00_83_13), .out(tmp01_41_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001693(.in0(tmp00_84_13), .in1(tmp00_85_13), .out(tmp01_42_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001694(.in0(tmp00_86_13), .in1(tmp00_87_13), .out(tmp01_43_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001695(.in0(tmp00_88_13), .in1(tmp00_89_13), .out(tmp01_44_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001696(.in0(tmp00_90_13), .in1(tmp00_91_13), .out(tmp01_45_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001697(.in0(tmp00_92_13), .in1(tmp00_93_13), .out(tmp01_46_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001698(.in0(tmp00_94_13), .in1(tmp00_95_13), .out(tmp01_47_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001699(.in0(tmp00_96_13), .in1(tmp00_97_13), .out(tmp01_48_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001700(.in0(tmp00_98_13), .in1(tmp00_99_13), .out(tmp01_49_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001701(.in0(tmp00_100_13), .in1(tmp00_101_13), .out(tmp01_50_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001702(.in0(tmp00_102_13), .in1(tmp00_103_13), .out(tmp01_51_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001703(.in0(tmp00_104_13), .in1(tmp00_105_13), .out(tmp01_52_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001704(.in0(tmp00_106_13), .in1(tmp00_107_13), .out(tmp01_53_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001705(.in0(tmp00_108_13), .in1(tmp00_109_13), .out(tmp01_54_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001706(.in0(tmp00_110_13), .in1(tmp00_111_13), .out(tmp01_55_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001707(.in0(tmp00_112_13), .in1(tmp00_113_13), .out(tmp01_56_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001708(.in0(tmp00_114_13), .in1(tmp00_115_13), .out(tmp01_57_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001709(.in0(tmp00_116_13), .in1(tmp00_117_13), .out(tmp01_58_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001710(.in0(tmp00_118_13), .in1(tmp00_119_13), .out(tmp01_59_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001711(.in0(tmp00_120_13), .in1(tmp00_121_13), .out(tmp01_60_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001712(.in0(tmp00_122_13), .in1(tmp00_123_13), .out(tmp01_61_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001713(.in0(tmp00_124_13), .in1(tmp00_125_13), .out(tmp01_62_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001714(.in0(tmp00_126_13), .in1(tmp00_127_13), .out(tmp01_63_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001715(.in0(tmp01_0_13), .in1(tmp01_1_13), .out(tmp02_0_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001716(.in0(tmp01_2_13), .in1(tmp01_3_13), .out(tmp02_1_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001717(.in0(tmp01_4_13), .in1(tmp01_5_13), .out(tmp02_2_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001718(.in0(tmp01_6_13), .in1(tmp01_7_13), .out(tmp02_3_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001719(.in0(tmp01_8_13), .in1(tmp01_9_13), .out(tmp02_4_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001720(.in0(tmp01_10_13), .in1(tmp01_11_13), .out(tmp02_5_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001721(.in0(tmp01_12_13), .in1(tmp01_13_13), .out(tmp02_6_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001722(.in0(tmp01_14_13), .in1(tmp01_15_13), .out(tmp02_7_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001723(.in0(tmp01_16_13), .in1(tmp01_17_13), .out(tmp02_8_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001724(.in0(tmp01_18_13), .in1(tmp01_19_13), .out(tmp02_9_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001725(.in0(tmp01_20_13), .in1(tmp01_21_13), .out(tmp02_10_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001726(.in0(tmp01_22_13), .in1(tmp01_23_13), .out(tmp02_11_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001727(.in0(tmp01_24_13), .in1(tmp01_25_13), .out(tmp02_12_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001728(.in0(tmp01_26_13), .in1(tmp01_27_13), .out(tmp02_13_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001729(.in0(tmp01_28_13), .in1(tmp01_29_13), .out(tmp02_14_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001730(.in0(tmp01_30_13), .in1(tmp01_31_13), .out(tmp02_15_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001731(.in0(tmp01_32_13), .in1(tmp01_33_13), .out(tmp02_16_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001732(.in0(tmp01_34_13), .in1(tmp01_35_13), .out(tmp02_17_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001733(.in0(tmp01_36_13), .in1(tmp01_37_13), .out(tmp02_18_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001734(.in0(tmp01_38_13), .in1(tmp01_39_13), .out(tmp02_19_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001735(.in0(tmp01_40_13), .in1(tmp01_41_13), .out(tmp02_20_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001736(.in0(tmp01_42_13), .in1(tmp01_43_13), .out(tmp02_21_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001737(.in0(tmp01_44_13), .in1(tmp01_45_13), .out(tmp02_22_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001738(.in0(tmp01_46_13), .in1(tmp01_47_13), .out(tmp02_23_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001739(.in0(tmp01_48_13), .in1(tmp01_49_13), .out(tmp02_24_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001740(.in0(tmp01_50_13), .in1(tmp01_51_13), .out(tmp02_25_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001741(.in0(tmp01_52_13), .in1(tmp01_53_13), .out(tmp02_26_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001742(.in0(tmp01_54_13), .in1(tmp01_55_13), .out(tmp02_27_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001743(.in0(tmp01_56_13), .in1(tmp01_57_13), .out(tmp02_28_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001744(.in0(tmp01_58_13), .in1(tmp01_59_13), .out(tmp02_29_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001745(.in0(tmp01_60_13), .in1(tmp01_61_13), .out(tmp02_30_13));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001746(.in0(tmp01_62_13), .in1(tmp01_63_13), .out(tmp02_31_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001747(.in0(tmp02_0_13), .in1(tmp02_1_13), .out(tmp03_0_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001748(.in0(tmp02_2_13), .in1(tmp02_3_13), .out(tmp03_1_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001749(.in0(tmp02_4_13), .in1(tmp02_5_13), .out(tmp03_2_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001750(.in0(tmp02_6_13), .in1(tmp02_7_13), .out(tmp03_3_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001751(.in0(tmp02_8_13), .in1(tmp02_9_13), .out(tmp03_4_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001752(.in0(tmp02_10_13), .in1(tmp02_11_13), .out(tmp03_5_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001753(.in0(tmp02_12_13), .in1(tmp02_13_13), .out(tmp03_6_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001754(.in0(tmp02_14_13), .in1(tmp02_15_13), .out(tmp03_7_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001755(.in0(tmp02_16_13), .in1(tmp02_17_13), .out(tmp03_8_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001756(.in0(tmp02_18_13), .in1(tmp02_19_13), .out(tmp03_9_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001757(.in0(tmp02_20_13), .in1(tmp02_21_13), .out(tmp03_10_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001758(.in0(tmp02_22_13), .in1(tmp02_23_13), .out(tmp03_11_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001759(.in0(tmp02_24_13), .in1(tmp02_25_13), .out(tmp03_12_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001760(.in0(tmp02_26_13), .in1(tmp02_27_13), .out(tmp03_13_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001761(.in0(tmp02_28_13), .in1(tmp02_29_13), .out(tmp03_14_13));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001762(.in0(tmp02_30_13), .in1(tmp02_31_13), .out(tmp03_15_13));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001763(.in0(tmp03_0_13), .in1(tmp03_1_13), .out(tmp04_0_13));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001764(.in0(tmp03_2_13), .in1(tmp03_3_13), .out(tmp04_1_13));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001765(.in0(tmp03_4_13), .in1(tmp03_5_13), .out(tmp04_2_13));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001766(.in0(tmp03_6_13), .in1(tmp03_7_13), .out(tmp04_3_13));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001767(.in0(tmp03_8_13), .in1(tmp03_9_13), .out(tmp04_4_13));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001768(.in0(tmp03_10_13), .in1(tmp03_11_13), .out(tmp04_5_13));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001769(.in0(tmp03_12_13), .in1(tmp03_13_13), .out(tmp04_6_13));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001770(.in0(tmp03_14_13), .in1(tmp03_15_13), .out(tmp04_7_13));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001771(.in0(tmp04_0_13), .in1(tmp04_1_13), .out(tmp05_0_13));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001772(.in0(tmp04_2_13), .in1(tmp04_3_13), .out(tmp05_1_13));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001773(.in0(tmp04_4_13), .in1(tmp04_5_13), .out(tmp05_2_13));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001774(.in0(tmp04_6_13), .in1(tmp04_7_13), .out(tmp05_3_13));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001775(.in0(tmp05_0_13), .in1(tmp05_1_13), .out(tmp06_0_13));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001776(.in0(tmp05_2_13), .in1(tmp05_3_13), .out(tmp06_1_13));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add001777(.in0(tmp06_0_13), .in1(tmp06_1_13), .out(tmp07_0_13));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001778(.in0(tmp00_0_14), .in1(tmp00_1_14), .out(tmp01_0_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001779(.in0(tmp00_2_14), .in1(tmp00_3_14), .out(tmp01_1_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001780(.in0(tmp00_4_14), .in1(tmp00_5_14), .out(tmp01_2_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001781(.in0(tmp00_6_14), .in1(tmp00_7_14), .out(tmp01_3_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001782(.in0(tmp00_8_14), .in1(tmp00_9_14), .out(tmp01_4_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001783(.in0(tmp00_10_14), .in1(tmp00_11_14), .out(tmp01_5_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001784(.in0(tmp00_12_14), .in1(tmp00_13_14), .out(tmp01_6_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001785(.in0(tmp00_14_14), .in1(tmp00_15_14), .out(tmp01_7_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001786(.in0(tmp00_16_14), .in1(tmp00_17_14), .out(tmp01_8_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001787(.in0(tmp00_18_14), .in1(tmp00_19_14), .out(tmp01_9_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001788(.in0(tmp00_20_14), .in1(tmp00_21_14), .out(tmp01_10_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001789(.in0(tmp00_22_14), .in1(tmp00_23_14), .out(tmp01_11_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001790(.in0(tmp00_24_14), .in1(tmp00_25_14), .out(tmp01_12_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001791(.in0(tmp00_26_14), .in1(tmp00_27_14), .out(tmp01_13_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001792(.in0(tmp00_28_14), .in1(tmp00_29_14), .out(tmp01_14_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001793(.in0(tmp00_30_14), .in1(tmp00_31_14), .out(tmp01_15_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001794(.in0(tmp00_32_14), .in1(tmp00_33_14), .out(tmp01_16_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001795(.in0(tmp00_34_14), .in1(tmp00_35_14), .out(tmp01_17_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001796(.in0(tmp00_36_14), .in1(tmp00_37_14), .out(tmp01_18_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001797(.in0(tmp00_38_14), .in1(tmp00_39_14), .out(tmp01_19_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001798(.in0(tmp00_40_14), .in1(tmp00_41_14), .out(tmp01_20_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001799(.in0(tmp00_42_14), .in1(tmp00_43_14), .out(tmp01_21_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001800(.in0(tmp00_44_14), .in1(tmp00_45_14), .out(tmp01_22_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001801(.in0(tmp00_46_14), .in1(tmp00_47_14), .out(tmp01_23_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001802(.in0(tmp00_48_14), .in1(tmp00_49_14), .out(tmp01_24_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001803(.in0(tmp00_50_14), .in1(tmp00_51_14), .out(tmp01_25_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001804(.in0(tmp00_52_14), .in1(tmp00_53_14), .out(tmp01_26_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001805(.in0(tmp00_54_14), .in1(tmp00_55_14), .out(tmp01_27_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001806(.in0(tmp00_56_14), .in1(tmp00_57_14), .out(tmp01_28_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001807(.in0(tmp00_58_14), .in1(tmp00_59_14), .out(tmp01_29_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001808(.in0(tmp00_60_14), .in1(tmp00_61_14), .out(tmp01_30_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001809(.in0(tmp00_62_14), .in1(tmp00_63_14), .out(tmp01_31_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001810(.in0(tmp00_64_14), .in1(tmp00_65_14), .out(tmp01_32_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001811(.in0(tmp00_66_14), .in1(tmp00_67_14), .out(tmp01_33_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001812(.in0(tmp00_68_14), .in1(tmp00_69_14), .out(tmp01_34_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001813(.in0(tmp00_70_14), .in1(tmp00_71_14), .out(tmp01_35_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001814(.in0(tmp00_72_14), .in1(tmp00_73_14), .out(tmp01_36_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001815(.in0(tmp00_74_14), .in1(tmp00_75_14), .out(tmp01_37_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001816(.in0(tmp00_76_14), .in1(tmp00_77_14), .out(tmp01_38_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001817(.in0(tmp00_78_14), .in1(tmp00_79_14), .out(tmp01_39_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001818(.in0(tmp00_80_14), .in1(tmp00_81_14), .out(tmp01_40_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001819(.in0(tmp00_82_14), .in1(tmp00_83_14), .out(tmp01_41_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001820(.in0(tmp00_84_14), .in1(tmp00_85_14), .out(tmp01_42_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001821(.in0(tmp00_86_14), .in1(tmp00_87_14), .out(tmp01_43_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001822(.in0(tmp00_88_14), .in1(tmp00_89_14), .out(tmp01_44_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001823(.in0(tmp00_90_14), .in1(tmp00_91_14), .out(tmp01_45_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001824(.in0(tmp00_92_14), .in1(tmp00_93_14), .out(tmp01_46_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001825(.in0(tmp00_94_14), .in1(tmp00_95_14), .out(tmp01_47_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001826(.in0(tmp00_96_14), .in1(tmp00_97_14), .out(tmp01_48_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001827(.in0(tmp00_98_14), .in1(tmp00_99_14), .out(tmp01_49_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001828(.in0(tmp00_100_14), .in1(tmp00_101_14), .out(tmp01_50_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001829(.in0(tmp00_102_14), .in1(tmp00_103_14), .out(tmp01_51_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001830(.in0(tmp00_104_14), .in1(tmp00_105_14), .out(tmp01_52_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001831(.in0(tmp00_106_14), .in1(tmp00_107_14), .out(tmp01_53_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001832(.in0(tmp00_108_14), .in1(tmp00_109_14), .out(tmp01_54_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001833(.in0(tmp00_110_14), .in1(tmp00_111_14), .out(tmp01_55_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001834(.in0(tmp00_112_14), .in1(tmp00_113_14), .out(tmp01_56_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001835(.in0(tmp00_114_14), .in1(tmp00_115_14), .out(tmp01_57_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001836(.in0(tmp00_116_14), .in1(tmp00_117_14), .out(tmp01_58_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001837(.in0(tmp00_118_14), .in1(tmp00_119_14), .out(tmp01_59_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001838(.in0(tmp00_120_14), .in1(tmp00_121_14), .out(tmp01_60_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001839(.in0(tmp00_122_14), .in1(tmp00_123_14), .out(tmp01_61_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001840(.in0(tmp00_124_14), .in1(tmp00_125_14), .out(tmp01_62_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001841(.in0(tmp00_126_14), .in1(tmp00_127_14), .out(tmp01_63_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001842(.in0(tmp01_0_14), .in1(tmp01_1_14), .out(tmp02_0_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001843(.in0(tmp01_2_14), .in1(tmp01_3_14), .out(tmp02_1_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001844(.in0(tmp01_4_14), .in1(tmp01_5_14), .out(tmp02_2_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001845(.in0(tmp01_6_14), .in1(tmp01_7_14), .out(tmp02_3_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001846(.in0(tmp01_8_14), .in1(tmp01_9_14), .out(tmp02_4_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001847(.in0(tmp01_10_14), .in1(tmp01_11_14), .out(tmp02_5_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001848(.in0(tmp01_12_14), .in1(tmp01_13_14), .out(tmp02_6_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001849(.in0(tmp01_14_14), .in1(tmp01_15_14), .out(tmp02_7_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001850(.in0(tmp01_16_14), .in1(tmp01_17_14), .out(tmp02_8_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001851(.in0(tmp01_18_14), .in1(tmp01_19_14), .out(tmp02_9_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001852(.in0(tmp01_20_14), .in1(tmp01_21_14), .out(tmp02_10_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001853(.in0(tmp01_22_14), .in1(tmp01_23_14), .out(tmp02_11_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001854(.in0(tmp01_24_14), .in1(tmp01_25_14), .out(tmp02_12_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001855(.in0(tmp01_26_14), .in1(tmp01_27_14), .out(tmp02_13_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001856(.in0(tmp01_28_14), .in1(tmp01_29_14), .out(tmp02_14_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001857(.in0(tmp01_30_14), .in1(tmp01_31_14), .out(tmp02_15_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001858(.in0(tmp01_32_14), .in1(tmp01_33_14), .out(tmp02_16_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001859(.in0(tmp01_34_14), .in1(tmp01_35_14), .out(tmp02_17_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001860(.in0(tmp01_36_14), .in1(tmp01_37_14), .out(tmp02_18_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001861(.in0(tmp01_38_14), .in1(tmp01_39_14), .out(tmp02_19_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001862(.in0(tmp01_40_14), .in1(tmp01_41_14), .out(tmp02_20_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001863(.in0(tmp01_42_14), .in1(tmp01_43_14), .out(tmp02_21_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001864(.in0(tmp01_44_14), .in1(tmp01_45_14), .out(tmp02_22_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001865(.in0(tmp01_46_14), .in1(tmp01_47_14), .out(tmp02_23_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001866(.in0(tmp01_48_14), .in1(tmp01_49_14), .out(tmp02_24_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001867(.in0(tmp01_50_14), .in1(tmp01_51_14), .out(tmp02_25_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001868(.in0(tmp01_52_14), .in1(tmp01_53_14), .out(tmp02_26_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001869(.in0(tmp01_54_14), .in1(tmp01_55_14), .out(tmp02_27_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001870(.in0(tmp01_56_14), .in1(tmp01_57_14), .out(tmp02_28_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001871(.in0(tmp01_58_14), .in1(tmp01_59_14), .out(tmp02_29_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001872(.in0(tmp01_60_14), .in1(tmp01_61_14), .out(tmp02_30_14));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001873(.in0(tmp01_62_14), .in1(tmp01_63_14), .out(tmp02_31_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001874(.in0(tmp02_0_14), .in1(tmp02_1_14), .out(tmp03_0_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001875(.in0(tmp02_2_14), .in1(tmp02_3_14), .out(tmp03_1_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001876(.in0(tmp02_4_14), .in1(tmp02_5_14), .out(tmp03_2_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001877(.in0(tmp02_6_14), .in1(tmp02_7_14), .out(tmp03_3_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001878(.in0(tmp02_8_14), .in1(tmp02_9_14), .out(tmp03_4_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001879(.in0(tmp02_10_14), .in1(tmp02_11_14), .out(tmp03_5_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001880(.in0(tmp02_12_14), .in1(tmp02_13_14), .out(tmp03_6_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001881(.in0(tmp02_14_14), .in1(tmp02_15_14), .out(tmp03_7_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001882(.in0(tmp02_16_14), .in1(tmp02_17_14), .out(tmp03_8_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001883(.in0(tmp02_18_14), .in1(tmp02_19_14), .out(tmp03_9_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001884(.in0(tmp02_20_14), .in1(tmp02_21_14), .out(tmp03_10_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001885(.in0(tmp02_22_14), .in1(tmp02_23_14), .out(tmp03_11_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001886(.in0(tmp02_24_14), .in1(tmp02_25_14), .out(tmp03_12_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001887(.in0(tmp02_26_14), .in1(tmp02_27_14), .out(tmp03_13_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001888(.in0(tmp02_28_14), .in1(tmp02_29_14), .out(tmp03_14_14));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add001889(.in0(tmp02_30_14), .in1(tmp02_31_14), .out(tmp03_15_14));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001890(.in0(tmp03_0_14), .in1(tmp03_1_14), .out(tmp04_0_14));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001891(.in0(tmp03_2_14), .in1(tmp03_3_14), .out(tmp04_1_14));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001892(.in0(tmp03_4_14), .in1(tmp03_5_14), .out(tmp04_2_14));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001893(.in0(tmp03_6_14), .in1(tmp03_7_14), .out(tmp04_3_14));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001894(.in0(tmp03_8_14), .in1(tmp03_9_14), .out(tmp04_4_14));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001895(.in0(tmp03_10_14), .in1(tmp03_11_14), .out(tmp04_5_14));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001896(.in0(tmp03_12_14), .in1(tmp03_13_14), .out(tmp04_6_14));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add001897(.in0(tmp03_14_14), .in1(tmp03_15_14), .out(tmp04_7_14));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001898(.in0(tmp04_0_14), .in1(tmp04_1_14), .out(tmp05_0_14));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001899(.in0(tmp04_2_14), .in1(tmp04_3_14), .out(tmp05_1_14));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001900(.in0(tmp04_4_14), .in1(tmp04_5_14), .out(tmp05_2_14));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add001901(.in0(tmp04_6_14), .in1(tmp04_7_14), .out(tmp05_3_14));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001902(.in0(tmp05_0_14), .in1(tmp05_1_14), .out(tmp06_0_14));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add001903(.in0(tmp05_2_14), .in1(tmp05_3_14), .out(tmp06_1_14));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add001904(.in0(tmp06_0_14), .in1(tmp06_1_14), .out(tmp07_0_14));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001905(.in0(tmp00_0_15), .in1(tmp00_1_15), .out(tmp01_0_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001906(.in0(tmp00_2_15), .in1(tmp00_3_15), .out(tmp01_1_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001907(.in0(tmp00_4_15), .in1(tmp00_5_15), .out(tmp01_2_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001908(.in0(tmp00_6_15), .in1(tmp00_7_15), .out(tmp01_3_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001909(.in0(tmp00_8_15), .in1(tmp00_9_15), .out(tmp01_4_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001910(.in0(tmp00_10_15), .in1(tmp00_11_15), .out(tmp01_5_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001911(.in0(tmp00_12_15), .in1(tmp00_13_15), .out(tmp01_6_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001912(.in0(tmp00_14_15), .in1(tmp00_15_15), .out(tmp01_7_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001913(.in0(tmp00_16_15), .in1(tmp00_17_15), .out(tmp01_8_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001914(.in0(tmp00_18_15), .in1(tmp00_19_15), .out(tmp01_9_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001915(.in0(tmp00_20_15), .in1(tmp00_21_15), .out(tmp01_10_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001916(.in0(tmp00_22_15), .in1(tmp00_23_15), .out(tmp01_11_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001917(.in0(tmp00_24_15), .in1(tmp00_25_15), .out(tmp01_12_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001918(.in0(tmp00_26_15), .in1(tmp00_27_15), .out(tmp01_13_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001919(.in0(tmp00_28_15), .in1(tmp00_29_15), .out(tmp01_14_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001920(.in0(tmp00_30_15), .in1(tmp00_31_15), .out(tmp01_15_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001921(.in0(tmp00_32_15), .in1(tmp00_33_15), .out(tmp01_16_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001922(.in0(tmp00_34_15), .in1(tmp00_35_15), .out(tmp01_17_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001923(.in0(tmp00_36_15), .in1(tmp00_37_15), .out(tmp01_18_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001924(.in0(tmp00_38_15), .in1(tmp00_39_15), .out(tmp01_19_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001925(.in0(tmp00_40_15), .in1(tmp00_41_15), .out(tmp01_20_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001926(.in0(tmp00_42_15), .in1(tmp00_43_15), .out(tmp01_21_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001927(.in0(tmp00_44_15), .in1(tmp00_45_15), .out(tmp01_22_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001928(.in0(tmp00_46_15), .in1(tmp00_47_15), .out(tmp01_23_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001929(.in0(tmp00_48_15), .in1(tmp00_49_15), .out(tmp01_24_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001930(.in0(tmp00_50_15), .in1(tmp00_51_15), .out(tmp01_25_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001931(.in0(tmp00_52_15), .in1(tmp00_53_15), .out(tmp01_26_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001932(.in0(tmp00_54_15), .in1(tmp00_55_15), .out(tmp01_27_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001933(.in0(tmp00_56_15), .in1(tmp00_57_15), .out(tmp01_28_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001934(.in0(tmp00_58_15), .in1(tmp00_59_15), .out(tmp01_29_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001935(.in0(tmp00_60_15), .in1(tmp00_61_15), .out(tmp01_30_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001936(.in0(tmp00_62_15), .in1(tmp00_63_15), .out(tmp01_31_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001937(.in0(tmp00_64_15), .in1(tmp00_65_15), .out(tmp01_32_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001938(.in0(tmp00_66_15), .in1(tmp00_67_15), .out(tmp01_33_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001939(.in0(tmp00_68_15), .in1(tmp00_69_15), .out(tmp01_34_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001940(.in0(tmp00_70_15), .in1(tmp00_71_15), .out(tmp01_35_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001941(.in0(tmp00_72_15), .in1(tmp00_73_15), .out(tmp01_36_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001942(.in0(tmp00_74_15), .in1(tmp00_75_15), .out(tmp01_37_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001943(.in0(tmp00_76_15), .in1(tmp00_77_15), .out(tmp01_38_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001944(.in0(tmp00_78_15), .in1(tmp00_79_15), .out(tmp01_39_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001945(.in0(tmp00_80_15), .in1(tmp00_81_15), .out(tmp01_40_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001946(.in0(tmp00_82_15), .in1(tmp00_83_15), .out(tmp01_41_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001947(.in0(tmp00_84_15), .in1(tmp00_85_15), .out(tmp01_42_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001948(.in0(tmp00_86_15), .in1(tmp00_87_15), .out(tmp01_43_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001949(.in0(tmp00_88_15), .in1(tmp00_89_15), .out(tmp01_44_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001950(.in0(tmp00_90_15), .in1(tmp00_91_15), .out(tmp01_45_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001951(.in0(tmp00_92_15), .in1(tmp00_93_15), .out(tmp01_46_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001952(.in0(tmp00_94_15), .in1(tmp00_95_15), .out(tmp01_47_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001953(.in0(tmp00_96_15), .in1(tmp00_97_15), .out(tmp01_48_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001954(.in0(tmp00_98_15), .in1(tmp00_99_15), .out(tmp01_49_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001955(.in0(tmp00_100_15), .in1(tmp00_101_15), .out(tmp01_50_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001956(.in0(tmp00_102_15), .in1(tmp00_103_15), .out(tmp01_51_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001957(.in0(tmp00_104_15), .in1(tmp00_105_15), .out(tmp01_52_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001958(.in0(tmp00_106_15), .in1(tmp00_107_15), .out(tmp01_53_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001959(.in0(tmp00_108_15), .in1(tmp00_109_15), .out(tmp01_54_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001960(.in0(tmp00_110_15), .in1(tmp00_111_15), .out(tmp01_55_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001961(.in0(tmp00_112_15), .in1(tmp00_113_15), .out(tmp01_56_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001962(.in0(tmp00_114_15), .in1(tmp00_115_15), .out(tmp01_57_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001963(.in0(tmp00_116_15), .in1(tmp00_117_15), .out(tmp01_58_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001964(.in0(tmp00_118_15), .in1(tmp00_119_15), .out(tmp01_59_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001965(.in0(tmp00_120_15), .in1(tmp00_121_15), .out(tmp01_60_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001966(.in0(tmp00_122_15), .in1(tmp00_123_15), .out(tmp01_61_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001967(.in0(tmp00_124_15), .in1(tmp00_125_15), .out(tmp01_62_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add001968(.in0(tmp00_126_15), .in1(tmp00_127_15), .out(tmp01_63_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001969(.in0(tmp01_0_15), .in1(tmp01_1_15), .out(tmp02_0_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001970(.in0(tmp01_2_15), .in1(tmp01_3_15), .out(tmp02_1_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001971(.in0(tmp01_4_15), .in1(tmp01_5_15), .out(tmp02_2_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001972(.in0(tmp01_6_15), .in1(tmp01_7_15), .out(tmp02_3_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001973(.in0(tmp01_8_15), .in1(tmp01_9_15), .out(tmp02_4_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001974(.in0(tmp01_10_15), .in1(tmp01_11_15), .out(tmp02_5_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001975(.in0(tmp01_12_15), .in1(tmp01_13_15), .out(tmp02_6_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001976(.in0(tmp01_14_15), .in1(tmp01_15_15), .out(tmp02_7_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001977(.in0(tmp01_16_15), .in1(tmp01_17_15), .out(tmp02_8_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001978(.in0(tmp01_18_15), .in1(tmp01_19_15), .out(tmp02_9_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001979(.in0(tmp01_20_15), .in1(tmp01_21_15), .out(tmp02_10_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001980(.in0(tmp01_22_15), .in1(tmp01_23_15), .out(tmp02_11_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001981(.in0(tmp01_24_15), .in1(tmp01_25_15), .out(tmp02_12_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001982(.in0(tmp01_26_15), .in1(tmp01_27_15), .out(tmp02_13_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001983(.in0(tmp01_28_15), .in1(tmp01_29_15), .out(tmp02_14_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001984(.in0(tmp01_30_15), .in1(tmp01_31_15), .out(tmp02_15_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001985(.in0(tmp01_32_15), .in1(tmp01_33_15), .out(tmp02_16_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001986(.in0(tmp01_34_15), .in1(tmp01_35_15), .out(tmp02_17_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001987(.in0(tmp01_36_15), .in1(tmp01_37_15), .out(tmp02_18_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001988(.in0(tmp01_38_15), .in1(tmp01_39_15), .out(tmp02_19_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001989(.in0(tmp01_40_15), .in1(tmp01_41_15), .out(tmp02_20_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001990(.in0(tmp01_42_15), .in1(tmp01_43_15), .out(tmp02_21_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001991(.in0(tmp01_44_15), .in1(tmp01_45_15), .out(tmp02_22_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001992(.in0(tmp01_46_15), .in1(tmp01_47_15), .out(tmp02_23_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001993(.in0(tmp01_48_15), .in1(tmp01_49_15), .out(tmp02_24_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001994(.in0(tmp01_50_15), .in1(tmp01_51_15), .out(tmp02_25_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001995(.in0(tmp01_52_15), .in1(tmp01_53_15), .out(tmp02_26_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001996(.in0(tmp01_54_15), .in1(tmp01_55_15), .out(tmp02_27_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001997(.in0(tmp01_56_15), .in1(tmp01_57_15), .out(tmp02_28_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001998(.in0(tmp01_58_15), .in1(tmp01_59_15), .out(tmp02_29_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add001999(.in0(tmp01_60_15), .in1(tmp01_61_15), .out(tmp02_30_15));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002000(.in0(tmp01_62_15), .in1(tmp01_63_15), .out(tmp02_31_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002001(.in0(tmp02_0_15), .in1(tmp02_1_15), .out(tmp03_0_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002002(.in0(tmp02_2_15), .in1(tmp02_3_15), .out(tmp03_1_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002003(.in0(tmp02_4_15), .in1(tmp02_5_15), .out(tmp03_2_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002004(.in0(tmp02_6_15), .in1(tmp02_7_15), .out(tmp03_3_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002005(.in0(tmp02_8_15), .in1(tmp02_9_15), .out(tmp03_4_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002006(.in0(tmp02_10_15), .in1(tmp02_11_15), .out(tmp03_5_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002007(.in0(tmp02_12_15), .in1(tmp02_13_15), .out(tmp03_6_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002008(.in0(tmp02_14_15), .in1(tmp02_15_15), .out(tmp03_7_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002009(.in0(tmp02_16_15), .in1(tmp02_17_15), .out(tmp03_8_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002010(.in0(tmp02_18_15), .in1(tmp02_19_15), .out(tmp03_9_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002011(.in0(tmp02_20_15), .in1(tmp02_21_15), .out(tmp03_10_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002012(.in0(tmp02_22_15), .in1(tmp02_23_15), .out(tmp03_11_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002013(.in0(tmp02_24_15), .in1(tmp02_25_15), .out(tmp03_12_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002014(.in0(tmp02_26_15), .in1(tmp02_27_15), .out(tmp03_13_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002015(.in0(tmp02_28_15), .in1(tmp02_29_15), .out(tmp03_14_15));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002016(.in0(tmp02_30_15), .in1(tmp02_31_15), .out(tmp03_15_15));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002017(.in0(tmp03_0_15), .in1(tmp03_1_15), .out(tmp04_0_15));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002018(.in0(tmp03_2_15), .in1(tmp03_3_15), .out(tmp04_1_15));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002019(.in0(tmp03_4_15), .in1(tmp03_5_15), .out(tmp04_2_15));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002020(.in0(tmp03_6_15), .in1(tmp03_7_15), .out(tmp04_3_15));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002021(.in0(tmp03_8_15), .in1(tmp03_9_15), .out(tmp04_4_15));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002022(.in0(tmp03_10_15), .in1(tmp03_11_15), .out(tmp04_5_15));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002023(.in0(tmp03_12_15), .in1(tmp03_13_15), .out(tmp04_6_15));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002024(.in0(tmp03_14_15), .in1(tmp03_15_15), .out(tmp04_7_15));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002025(.in0(tmp04_0_15), .in1(tmp04_1_15), .out(tmp05_0_15));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002026(.in0(tmp04_2_15), .in1(tmp04_3_15), .out(tmp05_1_15));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002027(.in0(tmp04_4_15), .in1(tmp04_5_15), .out(tmp05_2_15));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002028(.in0(tmp04_6_15), .in1(tmp04_7_15), .out(tmp05_3_15));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002029(.in0(tmp05_0_15), .in1(tmp05_1_15), .out(tmp06_0_15));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002030(.in0(tmp05_2_15), .in1(tmp05_3_15), .out(tmp06_1_15));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add002031(.in0(tmp06_0_15), .in1(tmp06_1_15), .out(tmp07_0_15));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002032(.in0(tmp00_0_16), .in1(tmp00_1_16), .out(tmp01_0_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002033(.in0(tmp00_2_16), .in1(tmp00_3_16), .out(tmp01_1_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002034(.in0(tmp00_4_16), .in1(tmp00_5_16), .out(tmp01_2_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002035(.in0(tmp00_6_16), .in1(tmp00_7_16), .out(tmp01_3_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002036(.in0(tmp00_8_16), .in1(tmp00_9_16), .out(tmp01_4_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002037(.in0(tmp00_10_16), .in1(tmp00_11_16), .out(tmp01_5_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002038(.in0(tmp00_12_16), .in1(tmp00_13_16), .out(tmp01_6_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002039(.in0(tmp00_14_16), .in1(tmp00_15_16), .out(tmp01_7_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002040(.in0(tmp00_16_16), .in1(tmp00_17_16), .out(tmp01_8_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002041(.in0(tmp00_18_16), .in1(tmp00_19_16), .out(tmp01_9_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002042(.in0(tmp00_20_16), .in1(tmp00_21_16), .out(tmp01_10_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002043(.in0(tmp00_22_16), .in1(tmp00_23_16), .out(tmp01_11_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002044(.in0(tmp00_24_16), .in1(tmp00_25_16), .out(tmp01_12_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002045(.in0(tmp00_26_16), .in1(tmp00_27_16), .out(tmp01_13_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002046(.in0(tmp00_28_16), .in1(tmp00_29_16), .out(tmp01_14_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002047(.in0(tmp00_30_16), .in1(tmp00_31_16), .out(tmp01_15_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002048(.in0(tmp00_32_16), .in1(tmp00_33_16), .out(tmp01_16_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002049(.in0(tmp00_34_16), .in1(tmp00_35_16), .out(tmp01_17_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002050(.in0(tmp00_36_16), .in1(tmp00_37_16), .out(tmp01_18_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002051(.in0(tmp00_38_16), .in1(tmp00_39_16), .out(tmp01_19_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002052(.in0(tmp00_40_16), .in1(tmp00_41_16), .out(tmp01_20_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002053(.in0(tmp00_42_16), .in1(tmp00_43_16), .out(tmp01_21_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002054(.in0(tmp00_44_16), .in1(tmp00_45_16), .out(tmp01_22_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002055(.in0(tmp00_46_16), .in1(tmp00_47_16), .out(tmp01_23_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002056(.in0(tmp00_48_16), .in1(tmp00_49_16), .out(tmp01_24_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002057(.in0(tmp00_50_16), .in1(tmp00_51_16), .out(tmp01_25_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002058(.in0(tmp00_52_16), .in1(tmp00_53_16), .out(tmp01_26_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002059(.in0(tmp00_54_16), .in1(tmp00_55_16), .out(tmp01_27_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002060(.in0(tmp00_56_16), .in1(tmp00_57_16), .out(tmp01_28_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002061(.in0(tmp00_58_16), .in1(tmp00_59_16), .out(tmp01_29_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002062(.in0(tmp00_60_16), .in1(tmp00_61_16), .out(tmp01_30_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002063(.in0(tmp00_62_16), .in1(tmp00_63_16), .out(tmp01_31_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002064(.in0(tmp00_64_16), .in1(tmp00_65_16), .out(tmp01_32_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002065(.in0(tmp00_66_16), .in1(tmp00_67_16), .out(tmp01_33_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002066(.in0(tmp00_68_16), .in1(tmp00_69_16), .out(tmp01_34_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002067(.in0(tmp00_70_16), .in1(tmp00_71_16), .out(tmp01_35_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002068(.in0(tmp00_72_16), .in1(tmp00_73_16), .out(tmp01_36_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002069(.in0(tmp00_74_16), .in1(tmp00_75_16), .out(tmp01_37_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002070(.in0(tmp00_76_16), .in1(tmp00_77_16), .out(tmp01_38_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002071(.in0(tmp00_78_16), .in1(tmp00_79_16), .out(tmp01_39_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002072(.in0(tmp00_80_16), .in1(tmp00_81_16), .out(tmp01_40_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002073(.in0(tmp00_82_16), .in1(tmp00_83_16), .out(tmp01_41_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002074(.in0(tmp00_84_16), .in1(tmp00_85_16), .out(tmp01_42_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002075(.in0(tmp00_86_16), .in1(tmp00_87_16), .out(tmp01_43_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002076(.in0(tmp00_88_16), .in1(tmp00_89_16), .out(tmp01_44_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002077(.in0(tmp00_90_16), .in1(tmp00_91_16), .out(tmp01_45_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002078(.in0(tmp00_92_16), .in1(tmp00_93_16), .out(tmp01_46_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002079(.in0(tmp00_94_16), .in1(tmp00_95_16), .out(tmp01_47_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002080(.in0(tmp00_96_16), .in1(tmp00_97_16), .out(tmp01_48_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002081(.in0(tmp00_98_16), .in1(tmp00_99_16), .out(tmp01_49_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002082(.in0(tmp00_100_16), .in1(tmp00_101_16), .out(tmp01_50_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002083(.in0(tmp00_102_16), .in1(tmp00_103_16), .out(tmp01_51_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002084(.in0(tmp00_104_16), .in1(tmp00_105_16), .out(tmp01_52_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002085(.in0(tmp00_106_16), .in1(tmp00_107_16), .out(tmp01_53_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002086(.in0(tmp00_108_16), .in1(tmp00_109_16), .out(tmp01_54_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002087(.in0(tmp00_110_16), .in1(tmp00_111_16), .out(tmp01_55_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002088(.in0(tmp00_112_16), .in1(tmp00_113_16), .out(tmp01_56_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002089(.in0(tmp00_114_16), .in1(tmp00_115_16), .out(tmp01_57_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002090(.in0(tmp00_116_16), .in1(tmp00_117_16), .out(tmp01_58_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002091(.in0(tmp00_118_16), .in1(tmp00_119_16), .out(tmp01_59_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002092(.in0(tmp00_120_16), .in1(tmp00_121_16), .out(tmp01_60_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002093(.in0(tmp00_122_16), .in1(tmp00_123_16), .out(tmp01_61_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002094(.in0(tmp00_124_16), .in1(tmp00_125_16), .out(tmp01_62_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002095(.in0(tmp00_126_16), .in1(tmp00_127_16), .out(tmp01_63_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002096(.in0(tmp01_0_16), .in1(tmp01_1_16), .out(tmp02_0_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002097(.in0(tmp01_2_16), .in1(tmp01_3_16), .out(tmp02_1_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002098(.in0(tmp01_4_16), .in1(tmp01_5_16), .out(tmp02_2_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002099(.in0(tmp01_6_16), .in1(tmp01_7_16), .out(tmp02_3_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002100(.in0(tmp01_8_16), .in1(tmp01_9_16), .out(tmp02_4_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002101(.in0(tmp01_10_16), .in1(tmp01_11_16), .out(tmp02_5_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002102(.in0(tmp01_12_16), .in1(tmp01_13_16), .out(tmp02_6_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002103(.in0(tmp01_14_16), .in1(tmp01_15_16), .out(tmp02_7_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002104(.in0(tmp01_16_16), .in1(tmp01_17_16), .out(tmp02_8_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002105(.in0(tmp01_18_16), .in1(tmp01_19_16), .out(tmp02_9_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002106(.in0(tmp01_20_16), .in1(tmp01_21_16), .out(tmp02_10_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002107(.in0(tmp01_22_16), .in1(tmp01_23_16), .out(tmp02_11_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002108(.in0(tmp01_24_16), .in1(tmp01_25_16), .out(tmp02_12_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002109(.in0(tmp01_26_16), .in1(tmp01_27_16), .out(tmp02_13_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002110(.in0(tmp01_28_16), .in1(tmp01_29_16), .out(tmp02_14_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002111(.in0(tmp01_30_16), .in1(tmp01_31_16), .out(tmp02_15_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002112(.in0(tmp01_32_16), .in1(tmp01_33_16), .out(tmp02_16_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002113(.in0(tmp01_34_16), .in1(tmp01_35_16), .out(tmp02_17_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002114(.in0(tmp01_36_16), .in1(tmp01_37_16), .out(tmp02_18_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002115(.in0(tmp01_38_16), .in1(tmp01_39_16), .out(tmp02_19_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002116(.in0(tmp01_40_16), .in1(tmp01_41_16), .out(tmp02_20_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002117(.in0(tmp01_42_16), .in1(tmp01_43_16), .out(tmp02_21_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002118(.in0(tmp01_44_16), .in1(tmp01_45_16), .out(tmp02_22_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002119(.in0(tmp01_46_16), .in1(tmp01_47_16), .out(tmp02_23_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002120(.in0(tmp01_48_16), .in1(tmp01_49_16), .out(tmp02_24_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002121(.in0(tmp01_50_16), .in1(tmp01_51_16), .out(tmp02_25_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002122(.in0(tmp01_52_16), .in1(tmp01_53_16), .out(tmp02_26_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002123(.in0(tmp01_54_16), .in1(tmp01_55_16), .out(tmp02_27_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002124(.in0(tmp01_56_16), .in1(tmp01_57_16), .out(tmp02_28_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002125(.in0(tmp01_58_16), .in1(tmp01_59_16), .out(tmp02_29_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002126(.in0(tmp01_60_16), .in1(tmp01_61_16), .out(tmp02_30_16));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002127(.in0(tmp01_62_16), .in1(tmp01_63_16), .out(tmp02_31_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002128(.in0(tmp02_0_16), .in1(tmp02_1_16), .out(tmp03_0_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002129(.in0(tmp02_2_16), .in1(tmp02_3_16), .out(tmp03_1_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002130(.in0(tmp02_4_16), .in1(tmp02_5_16), .out(tmp03_2_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002131(.in0(tmp02_6_16), .in1(tmp02_7_16), .out(tmp03_3_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002132(.in0(tmp02_8_16), .in1(tmp02_9_16), .out(tmp03_4_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002133(.in0(tmp02_10_16), .in1(tmp02_11_16), .out(tmp03_5_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002134(.in0(tmp02_12_16), .in1(tmp02_13_16), .out(tmp03_6_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002135(.in0(tmp02_14_16), .in1(tmp02_15_16), .out(tmp03_7_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002136(.in0(tmp02_16_16), .in1(tmp02_17_16), .out(tmp03_8_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002137(.in0(tmp02_18_16), .in1(tmp02_19_16), .out(tmp03_9_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002138(.in0(tmp02_20_16), .in1(tmp02_21_16), .out(tmp03_10_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002139(.in0(tmp02_22_16), .in1(tmp02_23_16), .out(tmp03_11_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002140(.in0(tmp02_24_16), .in1(tmp02_25_16), .out(tmp03_12_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002141(.in0(tmp02_26_16), .in1(tmp02_27_16), .out(tmp03_13_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002142(.in0(tmp02_28_16), .in1(tmp02_29_16), .out(tmp03_14_16));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002143(.in0(tmp02_30_16), .in1(tmp02_31_16), .out(tmp03_15_16));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002144(.in0(tmp03_0_16), .in1(tmp03_1_16), .out(tmp04_0_16));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002145(.in0(tmp03_2_16), .in1(tmp03_3_16), .out(tmp04_1_16));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002146(.in0(tmp03_4_16), .in1(tmp03_5_16), .out(tmp04_2_16));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002147(.in0(tmp03_6_16), .in1(tmp03_7_16), .out(tmp04_3_16));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002148(.in0(tmp03_8_16), .in1(tmp03_9_16), .out(tmp04_4_16));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002149(.in0(tmp03_10_16), .in1(tmp03_11_16), .out(tmp04_5_16));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002150(.in0(tmp03_12_16), .in1(tmp03_13_16), .out(tmp04_6_16));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002151(.in0(tmp03_14_16), .in1(tmp03_15_16), .out(tmp04_7_16));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002152(.in0(tmp04_0_16), .in1(tmp04_1_16), .out(tmp05_0_16));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002153(.in0(tmp04_2_16), .in1(tmp04_3_16), .out(tmp05_1_16));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002154(.in0(tmp04_4_16), .in1(tmp04_5_16), .out(tmp05_2_16));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002155(.in0(tmp04_6_16), .in1(tmp04_7_16), .out(tmp05_3_16));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002156(.in0(tmp05_0_16), .in1(tmp05_1_16), .out(tmp06_0_16));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002157(.in0(tmp05_2_16), .in1(tmp05_3_16), .out(tmp06_1_16));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add002158(.in0(tmp06_0_16), .in1(tmp06_1_16), .out(tmp07_0_16));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002159(.in0(tmp00_0_17), .in1(tmp00_1_17), .out(tmp01_0_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002160(.in0(tmp00_2_17), .in1(tmp00_3_17), .out(tmp01_1_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002161(.in0(tmp00_4_17), .in1(tmp00_5_17), .out(tmp01_2_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002162(.in0(tmp00_6_17), .in1(tmp00_7_17), .out(tmp01_3_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002163(.in0(tmp00_8_17), .in1(tmp00_9_17), .out(tmp01_4_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002164(.in0(tmp00_10_17), .in1(tmp00_11_17), .out(tmp01_5_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002165(.in0(tmp00_12_17), .in1(tmp00_13_17), .out(tmp01_6_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002166(.in0(tmp00_14_17), .in1(tmp00_15_17), .out(tmp01_7_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002167(.in0(tmp00_16_17), .in1(tmp00_17_17), .out(tmp01_8_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002168(.in0(tmp00_18_17), .in1(tmp00_19_17), .out(tmp01_9_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002169(.in0(tmp00_20_17), .in1(tmp00_21_17), .out(tmp01_10_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002170(.in0(tmp00_22_17), .in1(tmp00_23_17), .out(tmp01_11_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002171(.in0(tmp00_24_17), .in1(tmp00_25_17), .out(tmp01_12_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002172(.in0(tmp00_26_17), .in1(tmp00_27_17), .out(tmp01_13_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002173(.in0(tmp00_28_17), .in1(tmp00_29_17), .out(tmp01_14_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002174(.in0(tmp00_30_17), .in1(tmp00_31_17), .out(tmp01_15_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002175(.in0(tmp00_32_17), .in1(tmp00_33_17), .out(tmp01_16_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002176(.in0(tmp00_34_17), .in1(tmp00_35_17), .out(tmp01_17_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002177(.in0(tmp00_36_17), .in1(tmp00_37_17), .out(tmp01_18_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002178(.in0(tmp00_38_17), .in1(tmp00_39_17), .out(tmp01_19_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002179(.in0(tmp00_40_17), .in1(tmp00_41_17), .out(tmp01_20_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002180(.in0(tmp00_42_17), .in1(tmp00_43_17), .out(tmp01_21_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002181(.in0(tmp00_44_17), .in1(tmp00_45_17), .out(tmp01_22_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002182(.in0(tmp00_46_17), .in1(tmp00_47_17), .out(tmp01_23_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002183(.in0(tmp00_48_17), .in1(tmp00_49_17), .out(tmp01_24_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002184(.in0(tmp00_50_17), .in1(tmp00_51_17), .out(tmp01_25_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002185(.in0(tmp00_52_17), .in1(tmp00_53_17), .out(tmp01_26_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002186(.in0(tmp00_54_17), .in1(tmp00_55_17), .out(tmp01_27_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002187(.in0(tmp00_56_17), .in1(tmp00_57_17), .out(tmp01_28_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002188(.in0(tmp00_58_17), .in1(tmp00_59_17), .out(tmp01_29_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002189(.in0(tmp00_60_17), .in1(tmp00_61_17), .out(tmp01_30_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002190(.in0(tmp00_62_17), .in1(tmp00_63_17), .out(tmp01_31_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002191(.in0(tmp00_64_17), .in1(tmp00_65_17), .out(tmp01_32_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002192(.in0(tmp00_66_17), .in1(tmp00_67_17), .out(tmp01_33_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002193(.in0(tmp00_68_17), .in1(tmp00_69_17), .out(tmp01_34_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002194(.in0(tmp00_70_17), .in1(tmp00_71_17), .out(tmp01_35_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002195(.in0(tmp00_72_17), .in1(tmp00_73_17), .out(tmp01_36_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002196(.in0(tmp00_74_17), .in1(tmp00_75_17), .out(tmp01_37_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002197(.in0(tmp00_76_17), .in1(tmp00_77_17), .out(tmp01_38_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002198(.in0(tmp00_78_17), .in1(tmp00_79_17), .out(tmp01_39_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002199(.in0(tmp00_80_17), .in1(tmp00_81_17), .out(tmp01_40_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002200(.in0(tmp00_82_17), .in1(tmp00_83_17), .out(tmp01_41_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002201(.in0(tmp00_84_17), .in1(tmp00_85_17), .out(tmp01_42_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002202(.in0(tmp00_86_17), .in1(tmp00_87_17), .out(tmp01_43_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002203(.in0(tmp00_88_17), .in1(tmp00_89_17), .out(tmp01_44_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002204(.in0(tmp00_90_17), .in1(tmp00_91_17), .out(tmp01_45_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002205(.in0(tmp00_92_17), .in1(tmp00_93_17), .out(tmp01_46_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002206(.in0(tmp00_94_17), .in1(tmp00_95_17), .out(tmp01_47_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002207(.in0(tmp00_96_17), .in1(tmp00_97_17), .out(tmp01_48_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002208(.in0(tmp00_98_17), .in1(tmp00_99_17), .out(tmp01_49_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002209(.in0(tmp00_100_17), .in1(tmp00_101_17), .out(tmp01_50_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002210(.in0(tmp00_102_17), .in1(tmp00_103_17), .out(tmp01_51_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002211(.in0(tmp00_104_17), .in1(tmp00_105_17), .out(tmp01_52_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002212(.in0(tmp00_106_17), .in1(tmp00_107_17), .out(tmp01_53_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002213(.in0(tmp00_108_17), .in1(tmp00_109_17), .out(tmp01_54_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002214(.in0(tmp00_110_17), .in1(tmp00_111_17), .out(tmp01_55_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002215(.in0(tmp00_112_17), .in1(tmp00_113_17), .out(tmp01_56_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002216(.in0(tmp00_114_17), .in1(tmp00_115_17), .out(tmp01_57_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002217(.in0(tmp00_116_17), .in1(tmp00_117_17), .out(tmp01_58_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002218(.in0(tmp00_118_17), .in1(tmp00_119_17), .out(tmp01_59_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002219(.in0(tmp00_120_17), .in1(tmp00_121_17), .out(tmp01_60_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002220(.in0(tmp00_122_17), .in1(tmp00_123_17), .out(tmp01_61_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002221(.in0(tmp00_124_17), .in1(tmp00_125_17), .out(tmp01_62_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002222(.in0(tmp00_126_17), .in1(tmp00_127_17), .out(tmp01_63_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002223(.in0(tmp01_0_17), .in1(tmp01_1_17), .out(tmp02_0_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002224(.in0(tmp01_2_17), .in1(tmp01_3_17), .out(tmp02_1_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002225(.in0(tmp01_4_17), .in1(tmp01_5_17), .out(tmp02_2_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002226(.in0(tmp01_6_17), .in1(tmp01_7_17), .out(tmp02_3_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002227(.in0(tmp01_8_17), .in1(tmp01_9_17), .out(tmp02_4_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002228(.in0(tmp01_10_17), .in1(tmp01_11_17), .out(tmp02_5_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002229(.in0(tmp01_12_17), .in1(tmp01_13_17), .out(tmp02_6_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002230(.in0(tmp01_14_17), .in1(tmp01_15_17), .out(tmp02_7_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002231(.in0(tmp01_16_17), .in1(tmp01_17_17), .out(tmp02_8_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002232(.in0(tmp01_18_17), .in1(tmp01_19_17), .out(tmp02_9_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002233(.in0(tmp01_20_17), .in1(tmp01_21_17), .out(tmp02_10_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002234(.in0(tmp01_22_17), .in1(tmp01_23_17), .out(tmp02_11_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002235(.in0(tmp01_24_17), .in1(tmp01_25_17), .out(tmp02_12_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002236(.in0(tmp01_26_17), .in1(tmp01_27_17), .out(tmp02_13_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002237(.in0(tmp01_28_17), .in1(tmp01_29_17), .out(tmp02_14_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002238(.in0(tmp01_30_17), .in1(tmp01_31_17), .out(tmp02_15_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002239(.in0(tmp01_32_17), .in1(tmp01_33_17), .out(tmp02_16_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002240(.in0(tmp01_34_17), .in1(tmp01_35_17), .out(tmp02_17_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002241(.in0(tmp01_36_17), .in1(tmp01_37_17), .out(tmp02_18_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002242(.in0(tmp01_38_17), .in1(tmp01_39_17), .out(tmp02_19_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002243(.in0(tmp01_40_17), .in1(tmp01_41_17), .out(tmp02_20_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002244(.in0(tmp01_42_17), .in1(tmp01_43_17), .out(tmp02_21_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002245(.in0(tmp01_44_17), .in1(tmp01_45_17), .out(tmp02_22_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002246(.in0(tmp01_46_17), .in1(tmp01_47_17), .out(tmp02_23_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002247(.in0(tmp01_48_17), .in1(tmp01_49_17), .out(tmp02_24_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002248(.in0(tmp01_50_17), .in1(tmp01_51_17), .out(tmp02_25_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002249(.in0(tmp01_52_17), .in1(tmp01_53_17), .out(tmp02_26_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002250(.in0(tmp01_54_17), .in1(tmp01_55_17), .out(tmp02_27_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002251(.in0(tmp01_56_17), .in1(tmp01_57_17), .out(tmp02_28_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002252(.in0(tmp01_58_17), .in1(tmp01_59_17), .out(tmp02_29_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002253(.in0(tmp01_60_17), .in1(tmp01_61_17), .out(tmp02_30_17));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002254(.in0(tmp01_62_17), .in1(tmp01_63_17), .out(tmp02_31_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002255(.in0(tmp02_0_17), .in1(tmp02_1_17), .out(tmp03_0_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002256(.in0(tmp02_2_17), .in1(tmp02_3_17), .out(tmp03_1_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002257(.in0(tmp02_4_17), .in1(tmp02_5_17), .out(tmp03_2_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002258(.in0(tmp02_6_17), .in1(tmp02_7_17), .out(tmp03_3_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002259(.in0(tmp02_8_17), .in1(tmp02_9_17), .out(tmp03_4_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002260(.in0(tmp02_10_17), .in1(tmp02_11_17), .out(tmp03_5_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002261(.in0(tmp02_12_17), .in1(tmp02_13_17), .out(tmp03_6_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002262(.in0(tmp02_14_17), .in1(tmp02_15_17), .out(tmp03_7_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002263(.in0(tmp02_16_17), .in1(tmp02_17_17), .out(tmp03_8_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002264(.in0(tmp02_18_17), .in1(tmp02_19_17), .out(tmp03_9_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002265(.in0(tmp02_20_17), .in1(tmp02_21_17), .out(tmp03_10_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002266(.in0(tmp02_22_17), .in1(tmp02_23_17), .out(tmp03_11_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002267(.in0(tmp02_24_17), .in1(tmp02_25_17), .out(tmp03_12_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002268(.in0(tmp02_26_17), .in1(tmp02_27_17), .out(tmp03_13_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002269(.in0(tmp02_28_17), .in1(tmp02_29_17), .out(tmp03_14_17));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002270(.in0(tmp02_30_17), .in1(tmp02_31_17), .out(tmp03_15_17));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002271(.in0(tmp03_0_17), .in1(tmp03_1_17), .out(tmp04_0_17));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002272(.in0(tmp03_2_17), .in1(tmp03_3_17), .out(tmp04_1_17));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002273(.in0(tmp03_4_17), .in1(tmp03_5_17), .out(tmp04_2_17));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002274(.in0(tmp03_6_17), .in1(tmp03_7_17), .out(tmp04_3_17));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002275(.in0(tmp03_8_17), .in1(tmp03_9_17), .out(tmp04_4_17));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002276(.in0(tmp03_10_17), .in1(tmp03_11_17), .out(tmp04_5_17));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002277(.in0(tmp03_12_17), .in1(tmp03_13_17), .out(tmp04_6_17));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002278(.in0(tmp03_14_17), .in1(tmp03_15_17), .out(tmp04_7_17));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002279(.in0(tmp04_0_17), .in1(tmp04_1_17), .out(tmp05_0_17));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002280(.in0(tmp04_2_17), .in1(tmp04_3_17), .out(tmp05_1_17));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002281(.in0(tmp04_4_17), .in1(tmp04_5_17), .out(tmp05_2_17));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002282(.in0(tmp04_6_17), .in1(tmp04_7_17), .out(tmp05_3_17));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002283(.in0(tmp05_0_17), .in1(tmp05_1_17), .out(tmp06_0_17));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002284(.in0(tmp05_2_17), .in1(tmp05_3_17), .out(tmp06_1_17));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add002285(.in0(tmp06_0_17), .in1(tmp06_1_17), .out(tmp07_0_17));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002286(.in0(tmp00_0_18), .in1(tmp00_1_18), .out(tmp01_0_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002287(.in0(tmp00_2_18), .in1(tmp00_3_18), .out(tmp01_1_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002288(.in0(tmp00_4_18), .in1(tmp00_5_18), .out(tmp01_2_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002289(.in0(tmp00_6_18), .in1(tmp00_7_18), .out(tmp01_3_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002290(.in0(tmp00_8_18), .in1(tmp00_9_18), .out(tmp01_4_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002291(.in0(tmp00_10_18), .in1(tmp00_11_18), .out(tmp01_5_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002292(.in0(tmp00_12_18), .in1(tmp00_13_18), .out(tmp01_6_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002293(.in0(tmp00_14_18), .in1(tmp00_15_18), .out(tmp01_7_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002294(.in0(tmp00_16_18), .in1(tmp00_17_18), .out(tmp01_8_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002295(.in0(tmp00_18_18), .in1(tmp00_19_18), .out(tmp01_9_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002296(.in0(tmp00_20_18), .in1(tmp00_21_18), .out(tmp01_10_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002297(.in0(tmp00_22_18), .in1(tmp00_23_18), .out(tmp01_11_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002298(.in0(tmp00_24_18), .in1(tmp00_25_18), .out(tmp01_12_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002299(.in0(tmp00_26_18), .in1(tmp00_27_18), .out(tmp01_13_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002300(.in0(tmp00_28_18), .in1(tmp00_29_18), .out(tmp01_14_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002301(.in0(tmp00_30_18), .in1(tmp00_31_18), .out(tmp01_15_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002302(.in0(tmp00_32_18), .in1(tmp00_33_18), .out(tmp01_16_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002303(.in0(tmp00_34_18), .in1(tmp00_35_18), .out(tmp01_17_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002304(.in0(tmp00_36_18), .in1(tmp00_37_18), .out(tmp01_18_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002305(.in0(tmp00_38_18), .in1(tmp00_39_18), .out(tmp01_19_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002306(.in0(tmp00_40_18), .in1(tmp00_41_18), .out(tmp01_20_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002307(.in0(tmp00_42_18), .in1(tmp00_43_18), .out(tmp01_21_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002308(.in0(tmp00_44_18), .in1(tmp00_45_18), .out(tmp01_22_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002309(.in0(tmp00_46_18), .in1(tmp00_47_18), .out(tmp01_23_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002310(.in0(tmp00_48_18), .in1(tmp00_49_18), .out(tmp01_24_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002311(.in0(tmp00_50_18), .in1(tmp00_51_18), .out(tmp01_25_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002312(.in0(tmp00_52_18), .in1(tmp00_53_18), .out(tmp01_26_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002313(.in0(tmp00_54_18), .in1(tmp00_55_18), .out(tmp01_27_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002314(.in0(tmp00_56_18), .in1(tmp00_57_18), .out(tmp01_28_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002315(.in0(tmp00_58_18), .in1(tmp00_59_18), .out(tmp01_29_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002316(.in0(tmp00_60_18), .in1(tmp00_61_18), .out(tmp01_30_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002317(.in0(tmp00_62_18), .in1(tmp00_63_18), .out(tmp01_31_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002318(.in0(tmp00_64_18), .in1(tmp00_65_18), .out(tmp01_32_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002319(.in0(tmp00_66_18), .in1(tmp00_67_18), .out(tmp01_33_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002320(.in0(tmp00_68_18), .in1(tmp00_69_18), .out(tmp01_34_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002321(.in0(tmp00_70_18), .in1(tmp00_71_18), .out(tmp01_35_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002322(.in0(tmp00_72_18), .in1(tmp00_73_18), .out(tmp01_36_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002323(.in0(tmp00_74_18), .in1(tmp00_75_18), .out(tmp01_37_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002324(.in0(tmp00_76_18), .in1(tmp00_77_18), .out(tmp01_38_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002325(.in0(tmp00_78_18), .in1(tmp00_79_18), .out(tmp01_39_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002326(.in0(tmp00_80_18), .in1(tmp00_81_18), .out(tmp01_40_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002327(.in0(tmp00_82_18), .in1(tmp00_83_18), .out(tmp01_41_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002328(.in0(tmp00_84_18), .in1(tmp00_85_18), .out(tmp01_42_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002329(.in0(tmp00_86_18), .in1(tmp00_87_18), .out(tmp01_43_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002330(.in0(tmp00_88_18), .in1(tmp00_89_18), .out(tmp01_44_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002331(.in0(tmp00_90_18), .in1(tmp00_91_18), .out(tmp01_45_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002332(.in0(tmp00_92_18), .in1(tmp00_93_18), .out(tmp01_46_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002333(.in0(tmp00_94_18), .in1(tmp00_95_18), .out(tmp01_47_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002334(.in0(tmp00_96_18), .in1(tmp00_97_18), .out(tmp01_48_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002335(.in0(tmp00_98_18), .in1(tmp00_99_18), .out(tmp01_49_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002336(.in0(tmp00_100_18), .in1(tmp00_101_18), .out(tmp01_50_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002337(.in0(tmp00_102_18), .in1(tmp00_103_18), .out(tmp01_51_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002338(.in0(tmp00_104_18), .in1(tmp00_105_18), .out(tmp01_52_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002339(.in0(tmp00_106_18), .in1(tmp00_107_18), .out(tmp01_53_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002340(.in0(tmp00_108_18), .in1(tmp00_109_18), .out(tmp01_54_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002341(.in0(tmp00_110_18), .in1(tmp00_111_18), .out(tmp01_55_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002342(.in0(tmp00_112_18), .in1(tmp00_113_18), .out(tmp01_56_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002343(.in0(tmp00_114_18), .in1(tmp00_115_18), .out(tmp01_57_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002344(.in0(tmp00_116_18), .in1(tmp00_117_18), .out(tmp01_58_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002345(.in0(tmp00_118_18), .in1(tmp00_119_18), .out(tmp01_59_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002346(.in0(tmp00_120_18), .in1(tmp00_121_18), .out(tmp01_60_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002347(.in0(tmp00_122_18), .in1(tmp00_123_18), .out(tmp01_61_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002348(.in0(tmp00_124_18), .in1(tmp00_125_18), .out(tmp01_62_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002349(.in0(tmp00_126_18), .in1(tmp00_127_18), .out(tmp01_63_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002350(.in0(tmp01_0_18), .in1(tmp01_1_18), .out(tmp02_0_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002351(.in0(tmp01_2_18), .in1(tmp01_3_18), .out(tmp02_1_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002352(.in0(tmp01_4_18), .in1(tmp01_5_18), .out(tmp02_2_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002353(.in0(tmp01_6_18), .in1(tmp01_7_18), .out(tmp02_3_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002354(.in0(tmp01_8_18), .in1(tmp01_9_18), .out(tmp02_4_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002355(.in0(tmp01_10_18), .in1(tmp01_11_18), .out(tmp02_5_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002356(.in0(tmp01_12_18), .in1(tmp01_13_18), .out(tmp02_6_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002357(.in0(tmp01_14_18), .in1(tmp01_15_18), .out(tmp02_7_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002358(.in0(tmp01_16_18), .in1(tmp01_17_18), .out(tmp02_8_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002359(.in0(tmp01_18_18), .in1(tmp01_19_18), .out(tmp02_9_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002360(.in0(tmp01_20_18), .in1(tmp01_21_18), .out(tmp02_10_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002361(.in0(tmp01_22_18), .in1(tmp01_23_18), .out(tmp02_11_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002362(.in0(tmp01_24_18), .in1(tmp01_25_18), .out(tmp02_12_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002363(.in0(tmp01_26_18), .in1(tmp01_27_18), .out(tmp02_13_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002364(.in0(tmp01_28_18), .in1(tmp01_29_18), .out(tmp02_14_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002365(.in0(tmp01_30_18), .in1(tmp01_31_18), .out(tmp02_15_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002366(.in0(tmp01_32_18), .in1(tmp01_33_18), .out(tmp02_16_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002367(.in0(tmp01_34_18), .in1(tmp01_35_18), .out(tmp02_17_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002368(.in0(tmp01_36_18), .in1(tmp01_37_18), .out(tmp02_18_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002369(.in0(tmp01_38_18), .in1(tmp01_39_18), .out(tmp02_19_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002370(.in0(tmp01_40_18), .in1(tmp01_41_18), .out(tmp02_20_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002371(.in0(tmp01_42_18), .in1(tmp01_43_18), .out(tmp02_21_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002372(.in0(tmp01_44_18), .in1(tmp01_45_18), .out(tmp02_22_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002373(.in0(tmp01_46_18), .in1(tmp01_47_18), .out(tmp02_23_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002374(.in0(tmp01_48_18), .in1(tmp01_49_18), .out(tmp02_24_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002375(.in0(tmp01_50_18), .in1(tmp01_51_18), .out(tmp02_25_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002376(.in0(tmp01_52_18), .in1(tmp01_53_18), .out(tmp02_26_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002377(.in0(tmp01_54_18), .in1(tmp01_55_18), .out(tmp02_27_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002378(.in0(tmp01_56_18), .in1(tmp01_57_18), .out(tmp02_28_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002379(.in0(tmp01_58_18), .in1(tmp01_59_18), .out(tmp02_29_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002380(.in0(tmp01_60_18), .in1(tmp01_61_18), .out(tmp02_30_18));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002381(.in0(tmp01_62_18), .in1(tmp01_63_18), .out(tmp02_31_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002382(.in0(tmp02_0_18), .in1(tmp02_1_18), .out(tmp03_0_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002383(.in0(tmp02_2_18), .in1(tmp02_3_18), .out(tmp03_1_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002384(.in0(tmp02_4_18), .in1(tmp02_5_18), .out(tmp03_2_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002385(.in0(tmp02_6_18), .in1(tmp02_7_18), .out(tmp03_3_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002386(.in0(tmp02_8_18), .in1(tmp02_9_18), .out(tmp03_4_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002387(.in0(tmp02_10_18), .in1(tmp02_11_18), .out(tmp03_5_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002388(.in0(tmp02_12_18), .in1(tmp02_13_18), .out(tmp03_6_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002389(.in0(tmp02_14_18), .in1(tmp02_15_18), .out(tmp03_7_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002390(.in0(tmp02_16_18), .in1(tmp02_17_18), .out(tmp03_8_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002391(.in0(tmp02_18_18), .in1(tmp02_19_18), .out(tmp03_9_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002392(.in0(tmp02_20_18), .in1(tmp02_21_18), .out(tmp03_10_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002393(.in0(tmp02_22_18), .in1(tmp02_23_18), .out(tmp03_11_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002394(.in0(tmp02_24_18), .in1(tmp02_25_18), .out(tmp03_12_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002395(.in0(tmp02_26_18), .in1(tmp02_27_18), .out(tmp03_13_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002396(.in0(tmp02_28_18), .in1(tmp02_29_18), .out(tmp03_14_18));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002397(.in0(tmp02_30_18), .in1(tmp02_31_18), .out(tmp03_15_18));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002398(.in0(tmp03_0_18), .in1(tmp03_1_18), .out(tmp04_0_18));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002399(.in0(tmp03_2_18), .in1(tmp03_3_18), .out(tmp04_1_18));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002400(.in0(tmp03_4_18), .in1(tmp03_5_18), .out(tmp04_2_18));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002401(.in0(tmp03_6_18), .in1(tmp03_7_18), .out(tmp04_3_18));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002402(.in0(tmp03_8_18), .in1(tmp03_9_18), .out(tmp04_4_18));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002403(.in0(tmp03_10_18), .in1(tmp03_11_18), .out(tmp04_5_18));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002404(.in0(tmp03_12_18), .in1(tmp03_13_18), .out(tmp04_6_18));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002405(.in0(tmp03_14_18), .in1(tmp03_15_18), .out(tmp04_7_18));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002406(.in0(tmp04_0_18), .in1(tmp04_1_18), .out(tmp05_0_18));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002407(.in0(tmp04_2_18), .in1(tmp04_3_18), .out(tmp05_1_18));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002408(.in0(tmp04_4_18), .in1(tmp04_5_18), .out(tmp05_2_18));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002409(.in0(tmp04_6_18), .in1(tmp04_7_18), .out(tmp05_3_18));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002410(.in0(tmp05_0_18), .in1(tmp05_1_18), .out(tmp06_0_18));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002411(.in0(tmp05_2_18), .in1(tmp05_3_18), .out(tmp06_1_18));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add002412(.in0(tmp06_0_18), .in1(tmp06_1_18), .out(tmp07_0_18));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002413(.in0(tmp00_0_19), .in1(tmp00_1_19), .out(tmp01_0_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002414(.in0(tmp00_2_19), .in1(tmp00_3_19), .out(tmp01_1_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002415(.in0(tmp00_4_19), .in1(tmp00_5_19), .out(tmp01_2_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002416(.in0(tmp00_6_19), .in1(tmp00_7_19), .out(tmp01_3_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002417(.in0(tmp00_8_19), .in1(tmp00_9_19), .out(tmp01_4_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002418(.in0(tmp00_10_19), .in1(tmp00_11_19), .out(tmp01_5_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002419(.in0(tmp00_12_19), .in1(tmp00_13_19), .out(tmp01_6_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002420(.in0(tmp00_14_19), .in1(tmp00_15_19), .out(tmp01_7_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002421(.in0(tmp00_16_19), .in1(tmp00_17_19), .out(tmp01_8_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002422(.in0(tmp00_18_19), .in1(tmp00_19_19), .out(tmp01_9_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002423(.in0(tmp00_20_19), .in1(tmp00_21_19), .out(tmp01_10_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002424(.in0(tmp00_22_19), .in1(tmp00_23_19), .out(tmp01_11_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002425(.in0(tmp00_24_19), .in1(tmp00_25_19), .out(tmp01_12_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002426(.in0(tmp00_26_19), .in1(tmp00_27_19), .out(tmp01_13_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002427(.in0(tmp00_28_19), .in1(tmp00_29_19), .out(tmp01_14_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002428(.in0(tmp00_30_19), .in1(tmp00_31_19), .out(tmp01_15_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002429(.in0(tmp00_32_19), .in1(tmp00_33_19), .out(tmp01_16_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002430(.in0(tmp00_34_19), .in1(tmp00_35_19), .out(tmp01_17_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002431(.in0(tmp00_36_19), .in1(tmp00_37_19), .out(tmp01_18_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002432(.in0(tmp00_38_19), .in1(tmp00_39_19), .out(tmp01_19_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002433(.in0(tmp00_40_19), .in1(tmp00_41_19), .out(tmp01_20_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002434(.in0(tmp00_42_19), .in1(tmp00_43_19), .out(tmp01_21_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002435(.in0(tmp00_44_19), .in1(tmp00_45_19), .out(tmp01_22_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002436(.in0(tmp00_46_19), .in1(tmp00_47_19), .out(tmp01_23_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002437(.in0(tmp00_48_19), .in1(tmp00_49_19), .out(tmp01_24_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002438(.in0(tmp00_50_19), .in1(tmp00_51_19), .out(tmp01_25_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002439(.in0(tmp00_52_19), .in1(tmp00_53_19), .out(tmp01_26_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002440(.in0(tmp00_54_19), .in1(tmp00_55_19), .out(tmp01_27_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002441(.in0(tmp00_56_19), .in1(tmp00_57_19), .out(tmp01_28_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002442(.in0(tmp00_58_19), .in1(tmp00_59_19), .out(tmp01_29_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002443(.in0(tmp00_60_19), .in1(tmp00_61_19), .out(tmp01_30_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002444(.in0(tmp00_62_19), .in1(tmp00_63_19), .out(tmp01_31_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002445(.in0(tmp00_64_19), .in1(tmp00_65_19), .out(tmp01_32_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002446(.in0(tmp00_66_19), .in1(tmp00_67_19), .out(tmp01_33_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002447(.in0(tmp00_68_19), .in1(tmp00_69_19), .out(tmp01_34_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002448(.in0(tmp00_70_19), .in1(tmp00_71_19), .out(tmp01_35_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002449(.in0(tmp00_72_19), .in1(tmp00_73_19), .out(tmp01_36_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002450(.in0(tmp00_74_19), .in1(tmp00_75_19), .out(tmp01_37_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002451(.in0(tmp00_76_19), .in1(tmp00_77_19), .out(tmp01_38_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002452(.in0(tmp00_78_19), .in1(tmp00_79_19), .out(tmp01_39_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002453(.in0(tmp00_80_19), .in1(tmp00_81_19), .out(tmp01_40_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002454(.in0(tmp00_82_19), .in1(tmp00_83_19), .out(tmp01_41_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002455(.in0(tmp00_84_19), .in1(tmp00_85_19), .out(tmp01_42_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002456(.in0(tmp00_86_19), .in1(tmp00_87_19), .out(tmp01_43_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002457(.in0(tmp00_88_19), .in1(tmp00_89_19), .out(tmp01_44_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002458(.in0(tmp00_90_19), .in1(tmp00_91_19), .out(tmp01_45_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002459(.in0(tmp00_92_19), .in1(tmp00_93_19), .out(tmp01_46_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002460(.in0(tmp00_94_19), .in1(tmp00_95_19), .out(tmp01_47_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002461(.in0(tmp00_96_19), .in1(tmp00_97_19), .out(tmp01_48_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002462(.in0(tmp00_98_19), .in1(tmp00_99_19), .out(tmp01_49_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002463(.in0(tmp00_100_19), .in1(tmp00_101_19), .out(tmp01_50_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002464(.in0(tmp00_102_19), .in1(tmp00_103_19), .out(tmp01_51_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002465(.in0(tmp00_104_19), .in1(tmp00_105_19), .out(tmp01_52_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002466(.in0(tmp00_106_19), .in1(tmp00_107_19), .out(tmp01_53_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002467(.in0(tmp00_108_19), .in1(tmp00_109_19), .out(tmp01_54_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002468(.in0(tmp00_110_19), .in1(tmp00_111_19), .out(tmp01_55_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002469(.in0(tmp00_112_19), .in1(tmp00_113_19), .out(tmp01_56_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002470(.in0(tmp00_114_19), .in1(tmp00_115_19), .out(tmp01_57_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002471(.in0(tmp00_116_19), .in1(tmp00_117_19), .out(tmp01_58_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002472(.in0(tmp00_118_19), .in1(tmp00_119_19), .out(tmp01_59_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002473(.in0(tmp00_120_19), .in1(tmp00_121_19), .out(tmp01_60_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002474(.in0(tmp00_122_19), .in1(tmp00_123_19), .out(tmp01_61_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002475(.in0(tmp00_124_19), .in1(tmp00_125_19), .out(tmp01_62_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002476(.in0(tmp00_126_19), .in1(tmp00_127_19), .out(tmp01_63_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002477(.in0(tmp01_0_19), .in1(tmp01_1_19), .out(tmp02_0_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002478(.in0(tmp01_2_19), .in1(tmp01_3_19), .out(tmp02_1_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002479(.in0(tmp01_4_19), .in1(tmp01_5_19), .out(tmp02_2_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002480(.in0(tmp01_6_19), .in1(tmp01_7_19), .out(tmp02_3_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002481(.in0(tmp01_8_19), .in1(tmp01_9_19), .out(tmp02_4_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002482(.in0(tmp01_10_19), .in1(tmp01_11_19), .out(tmp02_5_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002483(.in0(tmp01_12_19), .in1(tmp01_13_19), .out(tmp02_6_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002484(.in0(tmp01_14_19), .in1(tmp01_15_19), .out(tmp02_7_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002485(.in0(tmp01_16_19), .in1(tmp01_17_19), .out(tmp02_8_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002486(.in0(tmp01_18_19), .in1(tmp01_19_19), .out(tmp02_9_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002487(.in0(tmp01_20_19), .in1(tmp01_21_19), .out(tmp02_10_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002488(.in0(tmp01_22_19), .in1(tmp01_23_19), .out(tmp02_11_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002489(.in0(tmp01_24_19), .in1(tmp01_25_19), .out(tmp02_12_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002490(.in0(tmp01_26_19), .in1(tmp01_27_19), .out(tmp02_13_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002491(.in0(tmp01_28_19), .in1(tmp01_29_19), .out(tmp02_14_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002492(.in0(tmp01_30_19), .in1(tmp01_31_19), .out(tmp02_15_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002493(.in0(tmp01_32_19), .in1(tmp01_33_19), .out(tmp02_16_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002494(.in0(tmp01_34_19), .in1(tmp01_35_19), .out(tmp02_17_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002495(.in0(tmp01_36_19), .in1(tmp01_37_19), .out(tmp02_18_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002496(.in0(tmp01_38_19), .in1(tmp01_39_19), .out(tmp02_19_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002497(.in0(tmp01_40_19), .in1(tmp01_41_19), .out(tmp02_20_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002498(.in0(tmp01_42_19), .in1(tmp01_43_19), .out(tmp02_21_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002499(.in0(tmp01_44_19), .in1(tmp01_45_19), .out(tmp02_22_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002500(.in0(tmp01_46_19), .in1(tmp01_47_19), .out(tmp02_23_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002501(.in0(tmp01_48_19), .in1(tmp01_49_19), .out(tmp02_24_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002502(.in0(tmp01_50_19), .in1(tmp01_51_19), .out(tmp02_25_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002503(.in0(tmp01_52_19), .in1(tmp01_53_19), .out(tmp02_26_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002504(.in0(tmp01_54_19), .in1(tmp01_55_19), .out(tmp02_27_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002505(.in0(tmp01_56_19), .in1(tmp01_57_19), .out(tmp02_28_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002506(.in0(tmp01_58_19), .in1(tmp01_59_19), .out(tmp02_29_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002507(.in0(tmp01_60_19), .in1(tmp01_61_19), .out(tmp02_30_19));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002508(.in0(tmp01_62_19), .in1(tmp01_63_19), .out(tmp02_31_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002509(.in0(tmp02_0_19), .in1(tmp02_1_19), .out(tmp03_0_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002510(.in0(tmp02_2_19), .in1(tmp02_3_19), .out(tmp03_1_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002511(.in0(tmp02_4_19), .in1(tmp02_5_19), .out(tmp03_2_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002512(.in0(tmp02_6_19), .in1(tmp02_7_19), .out(tmp03_3_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002513(.in0(tmp02_8_19), .in1(tmp02_9_19), .out(tmp03_4_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002514(.in0(tmp02_10_19), .in1(tmp02_11_19), .out(tmp03_5_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002515(.in0(tmp02_12_19), .in1(tmp02_13_19), .out(tmp03_6_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002516(.in0(tmp02_14_19), .in1(tmp02_15_19), .out(tmp03_7_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002517(.in0(tmp02_16_19), .in1(tmp02_17_19), .out(tmp03_8_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002518(.in0(tmp02_18_19), .in1(tmp02_19_19), .out(tmp03_9_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002519(.in0(tmp02_20_19), .in1(tmp02_21_19), .out(tmp03_10_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002520(.in0(tmp02_22_19), .in1(tmp02_23_19), .out(tmp03_11_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002521(.in0(tmp02_24_19), .in1(tmp02_25_19), .out(tmp03_12_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002522(.in0(tmp02_26_19), .in1(tmp02_27_19), .out(tmp03_13_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002523(.in0(tmp02_28_19), .in1(tmp02_29_19), .out(tmp03_14_19));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002524(.in0(tmp02_30_19), .in1(tmp02_31_19), .out(tmp03_15_19));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002525(.in0(tmp03_0_19), .in1(tmp03_1_19), .out(tmp04_0_19));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002526(.in0(tmp03_2_19), .in1(tmp03_3_19), .out(tmp04_1_19));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002527(.in0(tmp03_4_19), .in1(tmp03_5_19), .out(tmp04_2_19));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002528(.in0(tmp03_6_19), .in1(tmp03_7_19), .out(tmp04_3_19));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002529(.in0(tmp03_8_19), .in1(tmp03_9_19), .out(tmp04_4_19));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002530(.in0(tmp03_10_19), .in1(tmp03_11_19), .out(tmp04_5_19));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002531(.in0(tmp03_12_19), .in1(tmp03_13_19), .out(tmp04_6_19));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002532(.in0(tmp03_14_19), .in1(tmp03_15_19), .out(tmp04_7_19));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002533(.in0(tmp04_0_19), .in1(tmp04_1_19), .out(tmp05_0_19));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002534(.in0(tmp04_2_19), .in1(tmp04_3_19), .out(tmp05_1_19));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002535(.in0(tmp04_4_19), .in1(tmp04_5_19), .out(tmp05_2_19));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002536(.in0(tmp04_6_19), .in1(tmp04_7_19), .out(tmp05_3_19));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002537(.in0(tmp05_0_19), .in1(tmp05_1_19), .out(tmp06_0_19));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002538(.in0(tmp05_2_19), .in1(tmp05_3_19), .out(tmp06_1_19));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add002539(.in0(tmp06_0_19), .in1(tmp06_1_19), .out(tmp07_0_19));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002540(.in0(tmp00_0_20), .in1(tmp00_1_20), .out(tmp01_0_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002541(.in0(tmp00_2_20), .in1(tmp00_3_20), .out(tmp01_1_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002542(.in0(tmp00_4_20), .in1(tmp00_5_20), .out(tmp01_2_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002543(.in0(tmp00_6_20), .in1(tmp00_7_20), .out(tmp01_3_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002544(.in0(tmp00_8_20), .in1(tmp00_9_20), .out(tmp01_4_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002545(.in0(tmp00_10_20), .in1(tmp00_11_20), .out(tmp01_5_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002546(.in0(tmp00_12_20), .in1(tmp00_13_20), .out(tmp01_6_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002547(.in0(tmp00_14_20), .in1(tmp00_15_20), .out(tmp01_7_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002548(.in0(tmp00_16_20), .in1(tmp00_17_20), .out(tmp01_8_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002549(.in0(tmp00_18_20), .in1(tmp00_19_20), .out(tmp01_9_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002550(.in0(tmp00_20_20), .in1(tmp00_21_20), .out(tmp01_10_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002551(.in0(tmp00_22_20), .in1(tmp00_23_20), .out(tmp01_11_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002552(.in0(tmp00_24_20), .in1(tmp00_25_20), .out(tmp01_12_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002553(.in0(tmp00_26_20), .in1(tmp00_27_20), .out(tmp01_13_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002554(.in0(tmp00_28_20), .in1(tmp00_29_20), .out(tmp01_14_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002555(.in0(tmp00_30_20), .in1(tmp00_31_20), .out(tmp01_15_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002556(.in0(tmp00_32_20), .in1(tmp00_33_20), .out(tmp01_16_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002557(.in0(tmp00_34_20), .in1(tmp00_35_20), .out(tmp01_17_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002558(.in0(tmp00_36_20), .in1(tmp00_37_20), .out(tmp01_18_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002559(.in0(tmp00_38_20), .in1(tmp00_39_20), .out(tmp01_19_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002560(.in0(tmp00_40_20), .in1(tmp00_41_20), .out(tmp01_20_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002561(.in0(tmp00_42_20), .in1(tmp00_43_20), .out(tmp01_21_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002562(.in0(tmp00_44_20), .in1(tmp00_45_20), .out(tmp01_22_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002563(.in0(tmp00_46_20), .in1(tmp00_47_20), .out(tmp01_23_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002564(.in0(tmp00_48_20), .in1(tmp00_49_20), .out(tmp01_24_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002565(.in0(tmp00_50_20), .in1(tmp00_51_20), .out(tmp01_25_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002566(.in0(tmp00_52_20), .in1(tmp00_53_20), .out(tmp01_26_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002567(.in0(tmp00_54_20), .in1(tmp00_55_20), .out(tmp01_27_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002568(.in0(tmp00_56_20), .in1(tmp00_57_20), .out(tmp01_28_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002569(.in0(tmp00_58_20), .in1(tmp00_59_20), .out(tmp01_29_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002570(.in0(tmp00_60_20), .in1(tmp00_61_20), .out(tmp01_30_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002571(.in0(tmp00_62_20), .in1(tmp00_63_20), .out(tmp01_31_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002572(.in0(tmp00_64_20), .in1(tmp00_65_20), .out(tmp01_32_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002573(.in0(tmp00_66_20), .in1(tmp00_67_20), .out(tmp01_33_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002574(.in0(tmp00_68_20), .in1(tmp00_69_20), .out(tmp01_34_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002575(.in0(tmp00_70_20), .in1(tmp00_71_20), .out(tmp01_35_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002576(.in0(tmp00_72_20), .in1(tmp00_73_20), .out(tmp01_36_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002577(.in0(tmp00_74_20), .in1(tmp00_75_20), .out(tmp01_37_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002578(.in0(tmp00_76_20), .in1(tmp00_77_20), .out(tmp01_38_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002579(.in0(tmp00_78_20), .in1(tmp00_79_20), .out(tmp01_39_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002580(.in0(tmp00_80_20), .in1(tmp00_81_20), .out(tmp01_40_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002581(.in0(tmp00_82_20), .in1(tmp00_83_20), .out(tmp01_41_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002582(.in0(tmp00_84_20), .in1(tmp00_85_20), .out(tmp01_42_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002583(.in0(tmp00_86_20), .in1(tmp00_87_20), .out(tmp01_43_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002584(.in0(tmp00_88_20), .in1(tmp00_89_20), .out(tmp01_44_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002585(.in0(tmp00_90_20), .in1(tmp00_91_20), .out(tmp01_45_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002586(.in0(tmp00_92_20), .in1(tmp00_93_20), .out(tmp01_46_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002587(.in0(tmp00_94_20), .in1(tmp00_95_20), .out(tmp01_47_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002588(.in0(tmp00_96_20), .in1(tmp00_97_20), .out(tmp01_48_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002589(.in0(tmp00_98_20), .in1(tmp00_99_20), .out(tmp01_49_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002590(.in0(tmp00_100_20), .in1(tmp00_101_20), .out(tmp01_50_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002591(.in0(tmp00_102_20), .in1(tmp00_103_20), .out(tmp01_51_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002592(.in0(tmp00_104_20), .in1(tmp00_105_20), .out(tmp01_52_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002593(.in0(tmp00_106_20), .in1(tmp00_107_20), .out(tmp01_53_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002594(.in0(tmp00_108_20), .in1(tmp00_109_20), .out(tmp01_54_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002595(.in0(tmp00_110_20), .in1(tmp00_111_20), .out(tmp01_55_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002596(.in0(tmp00_112_20), .in1(tmp00_113_20), .out(tmp01_56_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002597(.in0(tmp00_114_20), .in1(tmp00_115_20), .out(tmp01_57_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002598(.in0(tmp00_116_20), .in1(tmp00_117_20), .out(tmp01_58_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002599(.in0(tmp00_118_20), .in1(tmp00_119_20), .out(tmp01_59_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002600(.in0(tmp00_120_20), .in1(tmp00_121_20), .out(tmp01_60_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002601(.in0(tmp00_122_20), .in1(tmp00_123_20), .out(tmp01_61_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002602(.in0(tmp00_124_20), .in1(tmp00_125_20), .out(tmp01_62_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002603(.in0(tmp00_126_20), .in1(tmp00_127_20), .out(tmp01_63_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002604(.in0(tmp01_0_20), .in1(tmp01_1_20), .out(tmp02_0_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002605(.in0(tmp01_2_20), .in1(tmp01_3_20), .out(tmp02_1_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002606(.in0(tmp01_4_20), .in1(tmp01_5_20), .out(tmp02_2_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002607(.in0(tmp01_6_20), .in1(tmp01_7_20), .out(tmp02_3_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002608(.in0(tmp01_8_20), .in1(tmp01_9_20), .out(tmp02_4_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002609(.in0(tmp01_10_20), .in1(tmp01_11_20), .out(tmp02_5_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002610(.in0(tmp01_12_20), .in1(tmp01_13_20), .out(tmp02_6_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002611(.in0(tmp01_14_20), .in1(tmp01_15_20), .out(tmp02_7_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002612(.in0(tmp01_16_20), .in1(tmp01_17_20), .out(tmp02_8_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002613(.in0(tmp01_18_20), .in1(tmp01_19_20), .out(tmp02_9_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002614(.in0(tmp01_20_20), .in1(tmp01_21_20), .out(tmp02_10_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002615(.in0(tmp01_22_20), .in1(tmp01_23_20), .out(tmp02_11_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002616(.in0(tmp01_24_20), .in1(tmp01_25_20), .out(tmp02_12_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002617(.in0(tmp01_26_20), .in1(tmp01_27_20), .out(tmp02_13_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002618(.in0(tmp01_28_20), .in1(tmp01_29_20), .out(tmp02_14_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002619(.in0(tmp01_30_20), .in1(tmp01_31_20), .out(tmp02_15_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002620(.in0(tmp01_32_20), .in1(tmp01_33_20), .out(tmp02_16_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002621(.in0(tmp01_34_20), .in1(tmp01_35_20), .out(tmp02_17_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002622(.in0(tmp01_36_20), .in1(tmp01_37_20), .out(tmp02_18_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002623(.in0(tmp01_38_20), .in1(tmp01_39_20), .out(tmp02_19_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002624(.in0(tmp01_40_20), .in1(tmp01_41_20), .out(tmp02_20_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002625(.in0(tmp01_42_20), .in1(tmp01_43_20), .out(tmp02_21_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002626(.in0(tmp01_44_20), .in1(tmp01_45_20), .out(tmp02_22_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002627(.in0(tmp01_46_20), .in1(tmp01_47_20), .out(tmp02_23_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002628(.in0(tmp01_48_20), .in1(tmp01_49_20), .out(tmp02_24_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002629(.in0(tmp01_50_20), .in1(tmp01_51_20), .out(tmp02_25_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002630(.in0(tmp01_52_20), .in1(tmp01_53_20), .out(tmp02_26_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002631(.in0(tmp01_54_20), .in1(tmp01_55_20), .out(tmp02_27_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002632(.in0(tmp01_56_20), .in1(tmp01_57_20), .out(tmp02_28_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002633(.in0(tmp01_58_20), .in1(tmp01_59_20), .out(tmp02_29_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002634(.in0(tmp01_60_20), .in1(tmp01_61_20), .out(tmp02_30_20));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002635(.in0(tmp01_62_20), .in1(tmp01_63_20), .out(tmp02_31_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002636(.in0(tmp02_0_20), .in1(tmp02_1_20), .out(tmp03_0_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002637(.in0(tmp02_2_20), .in1(tmp02_3_20), .out(tmp03_1_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002638(.in0(tmp02_4_20), .in1(tmp02_5_20), .out(tmp03_2_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002639(.in0(tmp02_6_20), .in1(tmp02_7_20), .out(tmp03_3_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002640(.in0(tmp02_8_20), .in1(tmp02_9_20), .out(tmp03_4_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002641(.in0(tmp02_10_20), .in1(tmp02_11_20), .out(tmp03_5_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002642(.in0(tmp02_12_20), .in1(tmp02_13_20), .out(tmp03_6_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002643(.in0(tmp02_14_20), .in1(tmp02_15_20), .out(tmp03_7_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002644(.in0(tmp02_16_20), .in1(tmp02_17_20), .out(tmp03_8_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002645(.in0(tmp02_18_20), .in1(tmp02_19_20), .out(tmp03_9_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002646(.in0(tmp02_20_20), .in1(tmp02_21_20), .out(tmp03_10_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002647(.in0(tmp02_22_20), .in1(tmp02_23_20), .out(tmp03_11_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002648(.in0(tmp02_24_20), .in1(tmp02_25_20), .out(tmp03_12_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002649(.in0(tmp02_26_20), .in1(tmp02_27_20), .out(tmp03_13_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002650(.in0(tmp02_28_20), .in1(tmp02_29_20), .out(tmp03_14_20));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002651(.in0(tmp02_30_20), .in1(tmp02_31_20), .out(tmp03_15_20));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002652(.in0(tmp03_0_20), .in1(tmp03_1_20), .out(tmp04_0_20));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002653(.in0(tmp03_2_20), .in1(tmp03_3_20), .out(tmp04_1_20));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002654(.in0(tmp03_4_20), .in1(tmp03_5_20), .out(tmp04_2_20));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002655(.in0(tmp03_6_20), .in1(tmp03_7_20), .out(tmp04_3_20));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002656(.in0(tmp03_8_20), .in1(tmp03_9_20), .out(tmp04_4_20));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002657(.in0(tmp03_10_20), .in1(tmp03_11_20), .out(tmp04_5_20));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002658(.in0(tmp03_12_20), .in1(tmp03_13_20), .out(tmp04_6_20));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002659(.in0(tmp03_14_20), .in1(tmp03_15_20), .out(tmp04_7_20));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002660(.in0(tmp04_0_20), .in1(tmp04_1_20), .out(tmp05_0_20));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002661(.in0(tmp04_2_20), .in1(tmp04_3_20), .out(tmp05_1_20));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002662(.in0(tmp04_4_20), .in1(tmp04_5_20), .out(tmp05_2_20));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002663(.in0(tmp04_6_20), .in1(tmp04_7_20), .out(tmp05_3_20));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002664(.in0(tmp05_0_20), .in1(tmp05_1_20), .out(tmp06_0_20));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002665(.in0(tmp05_2_20), .in1(tmp05_3_20), .out(tmp06_1_20));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add002666(.in0(tmp06_0_20), .in1(tmp06_1_20), .out(tmp07_0_20));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002667(.in0(tmp00_0_21), .in1(tmp00_1_21), .out(tmp01_0_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002668(.in0(tmp00_2_21), .in1(tmp00_3_21), .out(tmp01_1_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002669(.in0(tmp00_4_21), .in1(tmp00_5_21), .out(tmp01_2_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002670(.in0(tmp00_6_21), .in1(tmp00_7_21), .out(tmp01_3_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002671(.in0(tmp00_8_21), .in1(tmp00_9_21), .out(tmp01_4_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002672(.in0(tmp00_10_21), .in1(tmp00_11_21), .out(tmp01_5_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002673(.in0(tmp00_12_21), .in1(tmp00_13_21), .out(tmp01_6_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002674(.in0(tmp00_14_21), .in1(tmp00_15_21), .out(tmp01_7_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002675(.in0(tmp00_16_21), .in1(tmp00_17_21), .out(tmp01_8_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002676(.in0(tmp00_18_21), .in1(tmp00_19_21), .out(tmp01_9_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002677(.in0(tmp00_20_21), .in1(tmp00_21_21), .out(tmp01_10_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002678(.in0(tmp00_22_21), .in1(tmp00_23_21), .out(tmp01_11_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002679(.in0(tmp00_24_21), .in1(tmp00_25_21), .out(tmp01_12_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002680(.in0(tmp00_26_21), .in1(tmp00_27_21), .out(tmp01_13_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002681(.in0(tmp00_28_21), .in1(tmp00_29_21), .out(tmp01_14_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002682(.in0(tmp00_30_21), .in1(tmp00_31_21), .out(tmp01_15_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002683(.in0(tmp00_32_21), .in1(tmp00_33_21), .out(tmp01_16_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002684(.in0(tmp00_34_21), .in1(tmp00_35_21), .out(tmp01_17_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002685(.in0(tmp00_36_21), .in1(tmp00_37_21), .out(tmp01_18_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002686(.in0(tmp00_38_21), .in1(tmp00_39_21), .out(tmp01_19_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002687(.in0(tmp00_40_21), .in1(tmp00_41_21), .out(tmp01_20_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002688(.in0(tmp00_42_21), .in1(tmp00_43_21), .out(tmp01_21_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002689(.in0(tmp00_44_21), .in1(tmp00_45_21), .out(tmp01_22_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002690(.in0(tmp00_46_21), .in1(tmp00_47_21), .out(tmp01_23_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002691(.in0(tmp00_48_21), .in1(tmp00_49_21), .out(tmp01_24_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002692(.in0(tmp00_50_21), .in1(tmp00_51_21), .out(tmp01_25_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002693(.in0(tmp00_52_21), .in1(tmp00_53_21), .out(tmp01_26_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002694(.in0(tmp00_54_21), .in1(tmp00_55_21), .out(tmp01_27_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002695(.in0(tmp00_56_21), .in1(tmp00_57_21), .out(tmp01_28_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002696(.in0(tmp00_58_21), .in1(tmp00_59_21), .out(tmp01_29_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002697(.in0(tmp00_60_21), .in1(tmp00_61_21), .out(tmp01_30_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002698(.in0(tmp00_62_21), .in1(tmp00_63_21), .out(tmp01_31_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002699(.in0(tmp00_64_21), .in1(tmp00_65_21), .out(tmp01_32_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002700(.in0(tmp00_66_21), .in1(tmp00_67_21), .out(tmp01_33_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002701(.in0(tmp00_68_21), .in1(tmp00_69_21), .out(tmp01_34_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002702(.in0(tmp00_70_21), .in1(tmp00_71_21), .out(tmp01_35_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002703(.in0(tmp00_72_21), .in1(tmp00_73_21), .out(tmp01_36_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002704(.in0(tmp00_74_21), .in1(tmp00_75_21), .out(tmp01_37_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002705(.in0(tmp00_76_21), .in1(tmp00_77_21), .out(tmp01_38_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002706(.in0(tmp00_78_21), .in1(tmp00_79_21), .out(tmp01_39_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002707(.in0(tmp00_80_21), .in1(tmp00_81_21), .out(tmp01_40_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002708(.in0(tmp00_82_21), .in1(tmp00_83_21), .out(tmp01_41_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002709(.in0(tmp00_84_21), .in1(tmp00_85_21), .out(tmp01_42_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002710(.in0(tmp00_86_21), .in1(tmp00_87_21), .out(tmp01_43_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002711(.in0(tmp00_88_21), .in1(tmp00_89_21), .out(tmp01_44_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002712(.in0(tmp00_90_21), .in1(tmp00_91_21), .out(tmp01_45_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002713(.in0(tmp00_92_21), .in1(tmp00_93_21), .out(tmp01_46_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002714(.in0(tmp00_94_21), .in1(tmp00_95_21), .out(tmp01_47_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002715(.in0(tmp00_96_21), .in1(tmp00_97_21), .out(tmp01_48_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002716(.in0(tmp00_98_21), .in1(tmp00_99_21), .out(tmp01_49_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002717(.in0(tmp00_100_21), .in1(tmp00_101_21), .out(tmp01_50_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002718(.in0(tmp00_102_21), .in1(tmp00_103_21), .out(tmp01_51_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002719(.in0(tmp00_104_21), .in1(tmp00_105_21), .out(tmp01_52_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002720(.in0(tmp00_106_21), .in1(tmp00_107_21), .out(tmp01_53_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002721(.in0(tmp00_108_21), .in1(tmp00_109_21), .out(tmp01_54_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002722(.in0(tmp00_110_21), .in1(tmp00_111_21), .out(tmp01_55_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002723(.in0(tmp00_112_21), .in1(tmp00_113_21), .out(tmp01_56_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002724(.in0(tmp00_114_21), .in1(tmp00_115_21), .out(tmp01_57_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002725(.in0(tmp00_116_21), .in1(tmp00_117_21), .out(tmp01_58_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002726(.in0(tmp00_118_21), .in1(tmp00_119_21), .out(tmp01_59_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002727(.in0(tmp00_120_21), .in1(tmp00_121_21), .out(tmp01_60_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002728(.in0(tmp00_122_21), .in1(tmp00_123_21), .out(tmp01_61_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002729(.in0(tmp00_124_21), .in1(tmp00_125_21), .out(tmp01_62_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002730(.in0(tmp00_126_21), .in1(tmp00_127_21), .out(tmp01_63_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002731(.in0(tmp01_0_21), .in1(tmp01_1_21), .out(tmp02_0_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002732(.in0(tmp01_2_21), .in1(tmp01_3_21), .out(tmp02_1_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002733(.in0(tmp01_4_21), .in1(tmp01_5_21), .out(tmp02_2_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002734(.in0(tmp01_6_21), .in1(tmp01_7_21), .out(tmp02_3_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002735(.in0(tmp01_8_21), .in1(tmp01_9_21), .out(tmp02_4_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002736(.in0(tmp01_10_21), .in1(tmp01_11_21), .out(tmp02_5_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002737(.in0(tmp01_12_21), .in1(tmp01_13_21), .out(tmp02_6_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002738(.in0(tmp01_14_21), .in1(tmp01_15_21), .out(tmp02_7_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002739(.in0(tmp01_16_21), .in1(tmp01_17_21), .out(tmp02_8_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002740(.in0(tmp01_18_21), .in1(tmp01_19_21), .out(tmp02_9_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002741(.in0(tmp01_20_21), .in1(tmp01_21_21), .out(tmp02_10_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002742(.in0(tmp01_22_21), .in1(tmp01_23_21), .out(tmp02_11_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002743(.in0(tmp01_24_21), .in1(tmp01_25_21), .out(tmp02_12_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002744(.in0(tmp01_26_21), .in1(tmp01_27_21), .out(tmp02_13_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002745(.in0(tmp01_28_21), .in1(tmp01_29_21), .out(tmp02_14_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002746(.in0(tmp01_30_21), .in1(tmp01_31_21), .out(tmp02_15_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002747(.in0(tmp01_32_21), .in1(tmp01_33_21), .out(tmp02_16_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002748(.in0(tmp01_34_21), .in1(tmp01_35_21), .out(tmp02_17_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002749(.in0(tmp01_36_21), .in1(tmp01_37_21), .out(tmp02_18_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002750(.in0(tmp01_38_21), .in1(tmp01_39_21), .out(tmp02_19_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002751(.in0(tmp01_40_21), .in1(tmp01_41_21), .out(tmp02_20_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002752(.in0(tmp01_42_21), .in1(tmp01_43_21), .out(tmp02_21_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002753(.in0(tmp01_44_21), .in1(tmp01_45_21), .out(tmp02_22_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002754(.in0(tmp01_46_21), .in1(tmp01_47_21), .out(tmp02_23_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002755(.in0(tmp01_48_21), .in1(tmp01_49_21), .out(tmp02_24_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002756(.in0(tmp01_50_21), .in1(tmp01_51_21), .out(tmp02_25_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002757(.in0(tmp01_52_21), .in1(tmp01_53_21), .out(tmp02_26_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002758(.in0(tmp01_54_21), .in1(tmp01_55_21), .out(tmp02_27_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002759(.in0(tmp01_56_21), .in1(tmp01_57_21), .out(tmp02_28_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002760(.in0(tmp01_58_21), .in1(tmp01_59_21), .out(tmp02_29_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002761(.in0(tmp01_60_21), .in1(tmp01_61_21), .out(tmp02_30_21));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002762(.in0(tmp01_62_21), .in1(tmp01_63_21), .out(tmp02_31_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002763(.in0(tmp02_0_21), .in1(tmp02_1_21), .out(tmp03_0_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002764(.in0(tmp02_2_21), .in1(tmp02_3_21), .out(tmp03_1_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002765(.in0(tmp02_4_21), .in1(tmp02_5_21), .out(tmp03_2_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002766(.in0(tmp02_6_21), .in1(tmp02_7_21), .out(tmp03_3_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002767(.in0(tmp02_8_21), .in1(tmp02_9_21), .out(tmp03_4_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002768(.in0(tmp02_10_21), .in1(tmp02_11_21), .out(tmp03_5_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002769(.in0(tmp02_12_21), .in1(tmp02_13_21), .out(tmp03_6_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002770(.in0(tmp02_14_21), .in1(tmp02_15_21), .out(tmp03_7_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002771(.in0(tmp02_16_21), .in1(tmp02_17_21), .out(tmp03_8_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002772(.in0(tmp02_18_21), .in1(tmp02_19_21), .out(tmp03_9_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002773(.in0(tmp02_20_21), .in1(tmp02_21_21), .out(tmp03_10_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002774(.in0(tmp02_22_21), .in1(tmp02_23_21), .out(tmp03_11_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002775(.in0(tmp02_24_21), .in1(tmp02_25_21), .out(tmp03_12_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002776(.in0(tmp02_26_21), .in1(tmp02_27_21), .out(tmp03_13_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002777(.in0(tmp02_28_21), .in1(tmp02_29_21), .out(tmp03_14_21));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002778(.in0(tmp02_30_21), .in1(tmp02_31_21), .out(tmp03_15_21));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002779(.in0(tmp03_0_21), .in1(tmp03_1_21), .out(tmp04_0_21));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002780(.in0(tmp03_2_21), .in1(tmp03_3_21), .out(tmp04_1_21));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002781(.in0(tmp03_4_21), .in1(tmp03_5_21), .out(tmp04_2_21));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002782(.in0(tmp03_6_21), .in1(tmp03_7_21), .out(tmp04_3_21));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002783(.in0(tmp03_8_21), .in1(tmp03_9_21), .out(tmp04_4_21));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002784(.in0(tmp03_10_21), .in1(tmp03_11_21), .out(tmp04_5_21));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002785(.in0(tmp03_12_21), .in1(tmp03_13_21), .out(tmp04_6_21));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002786(.in0(tmp03_14_21), .in1(tmp03_15_21), .out(tmp04_7_21));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002787(.in0(tmp04_0_21), .in1(tmp04_1_21), .out(tmp05_0_21));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002788(.in0(tmp04_2_21), .in1(tmp04_3_21), .out(tmp05_1_21));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002789(.in0(tmp04_4_21), .in1(tmp04_5_21), .out(tmp05_2_21));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002790(.in0(tmp04_6_21), .in1(tmp04_7_21), .out(tmp05_3_21));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002791(.in0(tmp05_0_21), .in1(tmp05_1_21), .out(tmp06_0_21));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002792(.in0(tmp05_2_21), .in1(tmp05_3_21), .out(tmp06_1_21));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add002793(.in0(tmp06_0_21), .in1(tmp06_1_21), .out(tmp07_0_21));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002794(.in0(tmp00_0_22), .in1(tmp00_1_22), .out(tmp01_0_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002795(.in0(tmp00_2_22), .in1(tmp00_3_22), .out(tmp01_1_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002796(.in0(tmp00_4_22), .in1(tmp00_5_22), .out(tmp01_2_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002797(.in0(tmp00_6_22), .in1(tmp00_7_22), .out(tmp01_3_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002798(.in0(tmp00_8_22), .in1(tmp00_9_22), .out(tmp01_4_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002799(.in0(tmp00_10_22), .in1(tmp00_11_22), .out(tmp01_5_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002800(.in0(tmp00_12_22), .in1(tmp00_13_22), .out(tmp01_6_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002801(.in0(tmp00_14_22), .in1(tmp00_15_22), .out(tmp01_7_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002802(.in0(tmp00_16_22), .in1(tmp00_17_22), .out(tmp01_8_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002803(.in0(tmp00_18_22), .in1(tmp00_19_22), .out(tmp01_9_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002804(.in0(tmp00_20_22), .in1(tmp00_21_22), .out(tmp01_10_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002805(.in0(tmp00_22_22), .in1(tmp00_23_22), .out(tmp01_11_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002806(.in0(tmp00_24_22), .in1(tmp00_25_22), .out(tmp01_12_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002807(.in0(tmp00_26_22), .in1(tmp00_27_22), .out(tmp01_13_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002808(.in0(tmp00_28_22), .in1(tmp00_29_22), .out(tmp01_14_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002809(.in0(tmp00_30_22), .in1(tmp00_31_22), .out(tmp01_15_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002810(.in0(tmp00_32_22), .in1(tmp00_33_22), .out(tmp01_16_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002811(.in0(tmp00_34_22), .in1(tmp00_35_22), .out(tmp01_17_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002812(.in0(tmp00_36_22), .in1(tmp00_37_22), .out(tmp01_18_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002813(.in0(tmp00_38_22), .in1(tmp00_39_22), .out(tmp01_19_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002814(.in0(tmp00_40_22), .in1(tmp00_41_22), .out(tmp01_20_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002815(.in0(tmp00_42_22), .in1(tmp00_43_22), .out(tmp01_21_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002816(.in0(tmp00_44_22), .in1(tmp00_45_22), .out(tmp01_22_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002817(.in0(tmp00_46_22), .in1(tmp00_47_22), .out(tmp01_23_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002818(.in0(tmp00_48_22), .in1(tmp00_49_22), .out(tmp01_24_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002819(.in0(tmp00_50_22), .in1(tmp00_51_22), .out(tmp01_25_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002820(.in0(tmp00_52_22), .in1(tmp00_53_22), .out(tmp01_26_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002821(.in0(tmp00_54_22), .in1(tmp00_55_22), .out(tmp01_27_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002822(.in0(tmp00_56_22), .in1(tmp00_57_22), .out(tmp01_28_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002823(.in0(tmp00_58_22), .in1(tmp00_59_22), .out(tmp01_29_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002824(.in0(tmp00_60_22), .in1(tmp00_61_22), .out(tmp01_30_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002825(.in0(tmp00_62_22), .in1(tmp00_63_22), .out(tmp01_31_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002826(.in0(tmp00_64_22), .in1(tmp00_65_22), .out(tmp01_32_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002827(.in0(tmp00_66_22), .in1(tmp00_67_22), .out(tmp01_33_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002828(.in0(tmp00_68_22), .in1(tmp00_69_22), .out(tmp01_34_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002829(.in0(tmp00_70_22), .in1(tmp00_71_22), .out(tmp01_35_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002830(.in0(tmp00_72_22), .in1(tmp00_73_22), .out(tmp01_36_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002831(.in0(tmp00_74_22), .in1(tmp00_75_22), .out(tmp01_37_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002832(.in0(tmp00_76_22), .in1(tmp00_77_22), .out(tmp01_38_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002833(.in0(tmp00_78_22), .in1(tmp00_79_22), .out(tmp01_39_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002834(.in0(tmp00_80_22), .in1(tmp00_81_22), .out(tmp01_40_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002835(.in0(tmp00_82_22), .in1(tmp00_83_22), .out(tmp01_41_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002836(.in0(tmp00_84_22), .in1(tmp00_85_22), .out(tmp01_42_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002837(.in0(tmp00_86_22), .in1(tmp00_87_22), .out(tmp01_43_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002838(.in0(tmp00_88_22), .in1(tmp00_89_22), .out(tmp01_44_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002839(.in0(tmp00_90_22), .in1(tmp00_91_22), .out(tmp01_45_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002840(.in0(tmp00_92_22), .in1(tmp00_93_22), .out(tmp01_46_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002841(.in0(tmp00_94_22), .in1(tmp00_95_22), .out(tmp01_47_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002842(.in0(tmp00_96_22), .in1(tmp00_97_22), .out(tmp01_48_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002843(.in0(tmp00_98_22), .in1(tmp00_99_22), .out(tmp01_49_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002844(.in0(tmp00_100_22), .in1(tmp00_101_22), .out(tmp01_50_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002845(.in0(tmp00_102_22), .in1(tmp00_103_22), .out(tmp01_51_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002846(.in0(tmp00_104_22), .in1(tmp00_105_22), .out(tmp01_52_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002847(.in0(tmp00_106_22), .in1(tmp00_107_22), .out(tmp01_53_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002848(.in0(tmp00_108_22), .in1(tmp00_109_22), .out(tmp01_54_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002849(.in0(tmp00_110_22), .in1(tmp00_111_22), .out(tmp01_55_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002850(.in0(tmp00_112_22), .in1(tmp00_113_22), .out(tmp01_56_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002851(.in0(tmp00_114_22), .in1(tmp00_115_22), .out(tmp01_57_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002852(.in0(tmp00_116_22), .in1(tmp00_117_22), .out(tmp01_58_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002853(.in0(tmp00_118_22), .in1(tmp00_119_22), .out(tmp01_59_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002854(.in0(tmp00_120_22), .in1(tmp00_121_22), .out(tmp01_60_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002855(.in0(tmp00_122_22), .in1(tmp00_123_22), .out(tmp01_61_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002856(.in0(tmp00_124_22), .in1(tmp00_125_22), .out(tmp01_62_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002857(.in0(tmp00_126_22), .in1(tmp00_127_22), .out(tmp01_63_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002858(.in0(tmp01_0_22), .in1(tmp01_1_22), .out(tmp02_0_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002859(.in0(tmp01_2_22), .in1(tmp01_3_22), .out(tmp02_1_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002860(.in0(tmp01_4_22), .in1(tmp01_5_22), .out(tmp02_2_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002861(.in0(tmp01_6_22), .in1(tmp01_7_22), .out(tmp02_3_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002862(.in0(tmp01_8_22), .in1(tmp01_9_22), .out(tmp02_4_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002863(.in0(tmp01_10_22), .in1(tmp01_11_22), .out(tmp02_5_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002864(.in0(tmp01_12_22), .in1(tmp01_13_22), .out(tmp02_6_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002865(.in0(tmp01_14_22), .in1(tmp01_15_22), .out(tmp02_7_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002866(.in0(tmp01_16_22), .in1(tmp01_17_22), .out(tmp02_8_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002867(.in0(tmp01_18_22), .in1(tmp01_19_22), .out(tmp02_9_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002868(.in0(tmp01_20_22), .in1(tmp01_21_22), .out(tmp02_10_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002869(.in0(tmp01_22_22), .in1(tmp01_23_22), .out(tmp02_11_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002870(.in0(tmp01_24_22), .in1(tmp01_25_22), .out(tmp02_12_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002871(.in0(tmp01_26_22), .in1(tmp01_27_22), .out(tmp02_13_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002872(.in0(tmp01_28_22), .in1(tmp01_29_22), .out(tmp02_14_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002873(.in0(tmp01_30_22), .in1(tmp01_31_22), .out(tmp02_15_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002874(.in0(tmp01_32_22), .in1(tmp01_33_22), .out(tmp02_16_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002875(.in0(tmp01_34_22), .in1(tmp01_35_22), .out(tmp02_17_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002876(.in0(tmp01_36_22), .in1(tmp01_37_22), .out(tmp02_18_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002877(.in0(tmp01_38_22), .in1(tmp01_39_22), .out(tmp02_19_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002878(.in0(tmp01_40_22), .in1(tmp01_41_22), .out(tmp02_20_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002879(.in0(tmp01_42_22), .in1(tmp01_43_22), .out(tmp02_21_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002880(.in0(tmp01_44_22), .in1(tmp01_45_22), .out(tmp02_22_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002881(.in0(tmp01_46_22), .in1(tmp01_47_22), .out(tmp02_23_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002882(.in0(tmp01_48_22), .in1(tmp01_49_22), .out(tmp02_24_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002883(.in0(tmp01_50_22), .in1(tmp01_51_22), .out(tmp02_25_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002884(.in0(tmp01_52_22), .in1(tmp01_53_22), .out(tmp02_26_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002885(.in0(tmp01_54_22), .in1(tmp01_55_22), .out(tmp02_27_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002886(.in0(tmp01_56_22), .in1(tmp01_57_22), .out(tmp02_28_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002887(.in0(tmp01_58_22), .in1(tmp01_59_22), .out(tmp02_29_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002888(.in0(tmp01_60_22), .in1(tmp01_61_22), .out(tmp02_30_22));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002889(.in0(tmp01_62_22), .in1(tmp01_63_22), .out(tmp02_31_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002890(.in0(tmp02_0_22), .in1(tmp02_1_22), .out(tmp03_0_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002891(.in0(tmp02_2_22), .in1(tmp02_3_22), .out(tmp03_1_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002892(.in0(tmp02_4_22), .in1(tmp02_5_22), .out(tmp03_2_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002893(.in0(tmp02_6_22), .in1(tmp02_7_22), .out(tmp03_3_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002894(.in0(tmp02_8_22), .in1(tmp02_9_22), .out(tmp03_4_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002895(.in0(tmp02_10_22), .in1(tmp02_11_22), .out(tmp03_5_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002896(.in0(tmp02_12_22), .in1(tmp02_13_22), .out(tmp03_6_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002897(.in0(tmp02_14_22), .in1(tmp02_15_22), .out(tmp03_7_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002898(.in0(tmp02_16_22), .in1(tmp02_17_22), .out(tmp03_8_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002899(.in0(tmp02_18_22), .in1(tmp02_19_22), .out(tmp03_9_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002900(.in0(tmp02_20_22), .in1(tmp02_21_22), .out(tmp03_10_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002901(.in0(tmp02_22_22), .in1(tmp02_23_22), .out(tmp03_11_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002902(.in0(tmp02_24_22), .in1(tmp02_25_22), .out(tmp03_12_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002903(.in0(tmp02_26_22), .in1(tmp02_27_22), .out(tmp03_13_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002904(.in0(tmp02_28_22), .in1(tmp02_29_22), .out(tmp03_14_22));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add002905(.in0(tmp02_30_22), .in1(tmp02_31_22), .out(tmp03_15_22));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002906(.in0(tmp03_0_22), .in1(tmp03_1_22), .out(tmp04_0_22));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002907(.in0(tmp03_2_22), .in1(tmp03_3_22), .out(tmp04_1_22));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002908(.in0(tmp03_4_22), .in1(tmp03_5_22), .out(tmp04_2_22));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002909(.in0(tmp03_6_22), .in1(tmp03_7_22), .out(tmp04_3_22));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002910(.in0(tmp03_8_22), .in1(tmp03_9_22), .out(tmp04_4_22));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002911(.in0(tmp03_10_22), .in1(tmp03_11_22), .out(tmp04_5_22));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002912(.in0(tmp03_12_22), .in1(tmp03_13_22), .out(tmp04_6_22));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add002913(.in0(tmp03_14_22), .in1(tmp03_15_22), .out(tmp04_7_22));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002914(.in0(tmp04_0_22), .in1(tmp04_1_22), .out(tmp05_0_22));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002915(.in0(tmp04_2_22), .in1(tmp04_3_22), .out(tmp05_1_22));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002916(.in0(tmp04_4_22), .in1(tmp04_5_22), .out(tmp05_2_22));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add002917(.in0(tmp04_6_22), .in1(tmp04_7_22), .out(tmp05_3_22));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002918(.in0(tmp05_0_22), .in1(tmp05_1_22), .out(tmp06_0_22));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add002919(.in0(tmp05_2_22), .in1(tmp05_3_22), .out(tmp06_1_22));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add002920(.in0(tmp06_0_22), .in1(tmp06_1_22), .out(tmp07_0_22));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002921(.in0(tmp00_0_23), .in1(tmp00_1_23), .out(tmp01_0_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002922(.in0(tmp00_2_23), .in1(tmp00_3_23), .out(tmp01_1_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002923(.in0(tmp00_4_23), .in1(tmp00_5_23), .out(tmp01_2_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002924(.in0(tmp00_6_23), .in1(tmp00_7_23), .out(tmp01_3_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002925(.in0(tmp00_8_23), .in1(tmp00_9_23), .out(tmp01_4_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002926(.in0(tmp00_10_23), .in1(tmp00_11_23), .out(tmp01_5_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002927(.in0(tmp00_12_23), .in1(tmp00_13_23), .out(tmp01_6_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002928(.in0(tmp00_14_23), .in1(tmp00_15_23), .out(tmp01_7_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002929(.in0(tmp00_16_23), .in1(tmp00_17_23), .out(tmp01_8_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002930(.in0(tmp00_18_23), .in1(tmp00_19_23), .out(tmp01_9_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002931(.in0(tmp00_20_23), .in1(tmp00_21_23), .out(tmp01_10_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002932(.in0(tmp00_22_23), .in1(tmp00_23_23), .out(tmp01_11_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002933(.in0(tmp00_24_23), .in1(tmp00_25_23), .out(tmp01_12_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002934(.in0(tmp00_26_23), .in1(tmp00_27_23), .out(tmp01_13_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002935(.in0(tmp00_28_23), .in1(tmp00_29_23), .out(tmp01_14_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002936(.in0(tmp00_30_23), .in1(tmp00_31_23), .out(tmp01_15_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002937(.in0(tmp00_32_23), .in1(tmp00_33_23), .out(tmp01_16_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002938(.in0(tmp00_34_23), .in1(tmp00_35_23), .out(tmp01_17_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002939(.in0(tmp00_36_23), .in1(tmp00_37_23), .out(tmp01_18_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002940(.in0(tmp00_38_23), .in1(tmp00_39_23), .out(tmp01_19_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002941(.in0(tmp00_40_23), .in1(tmp00_41_23), .out(tmp01_20_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002942(.in0(tmp00_42_23), .in1(tmp00_43_23), .out(tmp01_21_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002943(.in0(tmp00_44_23), .in1(tmp00_45_23), .out(tmp01_22_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002944(.in0(tmp00_46_23), .in1(tmp00_47_23), .out(tmp01_23_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002945(.in0(tmp00_48_23), .in1(tmp00_49_23), .out(tmp01_24_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002946(.in0(tmp00_50_23), .in1(tmp00_51_23), .out(tmp01_25_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002947(.in0(tmp00_52_23), .in1(tmp00_53_23), .out(tmp01_26_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002948(.in0(tmp00_54_23), .in1(tmp00_55_23), .out(tmp01_27_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002949(.in0(tmp00_56_23), .in1(tmp00_57_23), .out(tmp01_28_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002950(.in0(tmp00_58_23), .in1(tmp00_59_23), .out(tmp01_29_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002951(.in0(tmp00_60_23), .in1(tmp00_61_23), .out(tmp01_30_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002952(.in0(tmp00_62_23), .in1(tmp00_63_23), .out(tmp01_31_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002953(.in0(tmp00_64_23), .in1(tmp00_65_23), .out(tmp01_32_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002954(.in0(tmp00_66_23), .in1(tmp00_67_23), .out(tmp01_33_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002955(.in0(tmp00_68_23), .in1(tmp00_69_23), .out(tmp01_34_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002956(.in0(tmp00_70_23), .in1(tmp00_71_23), .out(tmp01_35_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002957(.in0(tmp00_72_23), .in1(tmp00_73_23), .out(tmp01_36_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002958(.in0(tmp00_74_23), .in1(tmp00_75_23), .out(tmp01_37_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002959(.in0(tmp00_76_23), .in1(tmp00_77_23), .out(tmp01_38_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002960(.in0(tmp00_78_23), .in1(tmp00_79_23), .out(tmp01_39_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002961(.in0(tmp00_80_23), .in1(tmp00_81_23), .out(tmp01_40_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002962(.in0(tmp00_82_23), .in1(tmp00_83_23), .out(tmp01_41_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002963(.in0(tmp00_84_23), .in1(tmp00_85_23), .out(tmp01_42_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002964(.in0(tmp00_86_23), .in1(tmp00_87_23), .out(tmp01_43_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002965(.in0(tmp00_88_23), .in1(tmp00_89_23), .out(tmp01_44_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002966(.in0(tmp00_90_23), .in1(tmp00_91_23), .out(tmp01_45_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002967(.in0(tmp00_92_23), .in1(tmp00_93_23), .out(tmp01_46_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002968(.in0(tmp00_94_23), .in1(tmp00_95_23), .out(tmp01_47_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002969(.in0(tmp00_96_23), .in1(tmp00_97_23), .out(tmp01_48_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002970(.in0(tmp00_98_23), .in1(tmp00_99_23), .out(tmp01_49_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002971(.in0(tmp00_100_23), .in1(tmp00_101_23), .out(tmp01_50_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002972(.in0(tmp00_102_23), .in1(tmp00_103_23), .out(tmp01_51_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002973(.in0(tmp00_104_23), .in1(tmp00_105_23), .out(tmp01_52_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002974(.in0(tmp00_106_23), .in1(tmp00_107_23), .out(tmp01_53_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002975(.in0(tmp00_108_23), .in1(tmp00_109_23), .out(tmp01_54_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002976(.in0(tmp00_110_23), .in1(tmp00_111_23), .out(tmp01_55_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002977(.in0(tmp00_112_23), .in1(tmp00_113_23), .out(tmp01_56_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002978(.in0(tmp00_114_23), .in1(tmp00_115_23), .out(tmp01_57_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002979(.in0(tmp00_116_23), .in1(tmp00_117_23), .out(tmp01_58_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002980(.in0(tmp00_118_23), .in1(tmp00_119_23), .out(tmp01_59_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002981(.in0(tmp00_120_23), .in1(tmp00_121_23), .out(tmp01_60_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002982(.in0(tmp00_122_23), .in1(tmp00_123_23), .out(tmp01_61_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002983(.in0(tmp00_124_23), .in1(tmp00_125_23), .out(tmp01_62_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add002984(.in0(tmp00_126_23), .in1(tmp00_127_23), .out(tmp01_63_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002985(.in0(tmp01_0_23), .in1(tmp01_1_23), .out(tmp02_0_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002986(.in0(tmp01_2_23), .in1(tmp01_3_23), .out(tmp02_1_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002987(.in0(tmp01_4_23), .in1(tmp01_5_23), .out(tmp02_2_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002988(.in0(tmp01_6_23), .in1(tmp01_7_23), .out(tmp02_3_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002989(.in0(tmp01_8_23), .in1(tmp01_9_23), .out(tmp02_4_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002990(.in0(tmp01_10_23), .in1(tmp01_11_23), .out(tmp02_5_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002991(.in0(tmp01_12_23), .in1(tmp01_13_23), .out(tmp02_6_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002992(.in0(tmp01_14_23), .in1(tmp01_15_23), .out(tmp02_7_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002993(.in0(tmp01_16_23), .in1(tmp01_17_23), .out(tmp02_8_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002994(.in0(tmp01_18_23), .in1(tmp01_19_23), .out(tmp02_9_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002995(.in0(tmp01_20_23), .in1(tmp01_21_23), .out(tmp02_10_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002996(.in0(tmp01_22_23), .in1(tmp01_23_23), .out(tmp02_11_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002997(.in0(tmp01_24_23), .in1(tmp01_25_23), .out(tmp02_12_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002998(.in0(tmp01_26_23), .in1(tmp01_27_23), .out(tmp02_13_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add002999(.in0(tmp01_28_23), .in1(tmp01_29_23), .out(tmp02_14_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003000(.in0(tmp01_30_23), .in1(tmp01_31_23), .out(tmp02_15_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003001(.in0(tmp01_32_23), .in1(tmp01_33_23), .out(tmp02_16_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003002(.in0(tmp01_34_23), .in1(tmp01_35_23), .out(tmp02_17_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003003(.in0(tmp01_36_23), .in1(tmp01_37_23), .out(tmp02_18_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003004(.in0(tmp01_38_23), .in1(tmp01_39_23), .out(tmp02_19_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003005(.in0(tmp01_40_23), .in1(tmp01_41_23), .out(tmp02_20_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003006(.in0(tmp01_42_23), .in1(tmp01_43_23), .out(tmp02_21_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003007(.in0(tmp01_44_23), .in1(tmp01_45_23), .out(tmp02_22_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003008(.in0(tmp01_46_23), .in1(tmp01_47_23), .out(tmp02_23_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003009(.in0(tmp01_48_23), .in1(tmp01_49_23), .out(tmp02_24_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003010(.in0(tmp01_50_23), .in1(tmp01_51_23), .out(tmp02_25_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003011(.in0(tmp01_52_23), .in1(tmp01_53_23), .out(tmp02_26_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003012(.in0(tmp01_54_23), .in1(tmp01_55_23), .out(tmp02_27_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003013(.in0(tmp01_56_23), .in1(tmp01_57_23), .out(tmp02_28_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003014(.in0(tmp01_58_23), .in1(tmp01_59_23), .out(tmp02_29_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003015(.in0(tmp01_60_23), .in1(tmp01_61_23), .out(tmp02_30_23));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003016(.in0(tmp01_62_23), .in1(tmp01_63_23), .out(tmp02_31_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003017(.in0(tmp02_0_23), .in1(tmp02_1_23), .out(tmp03_0_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003018(.in0(tmp02_2_23), .in1(tmp02_3_23), .out(tmp03_1_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003019(.in0(tmp02_4_23), .in1(tmp02_5_23), .out(tmp03_2_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003020(.in0(tmp02_6_23), .in1(tmp02_7_23), .out(tmp03_3_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003021(.in0(tmp02_8_23), .in1(tmp02_9_23), .out(tmp03_4_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003022(.in0(tmp02_10_23), .in1(tmp02_11_23), .out(tmp03_5_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003023(.in0(tmp02_12_23), .in1(tmp02_13_23), .out(tmp03_6_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003024(.in0(tmp02_14_23), .in1(tmp02_15_23), .out(tmp03_7_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003025(.in0(tmp02_16_23), .in1(tmp02_17_23), .out(tmp03_8_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003026(.in0(tmp02_18_23), .in1(tmp02_19_23), .out(tmp03_9_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003027(.in0(tmp02_20_23), .in1(tmp02_21_23), .out(tmp03_10_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003028(.in0(tmp02_22_23), .in1(tmp02_23_23), .out(tmp03_11_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003029(.in0(tmp02_24_23), .in1(tmp02_25_23), .out(tmp03_12_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003030(.in0(tmp02_26_23), .in1(tmp02_27_23), .out(tmp03_13_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003031(.in0(tmp02_28_23), .in1(tmp02_29_23), .out(tmp03_14_23));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003032(.in0(tmp02_30_23), .in1(tmp02_31_23), .out(tmp03_15_23));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003033(.in0(tmp03_0_23), .in1(tmp03_1_23), .out(tmp04_0_23));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003034(.in0(tmp03_2_23), .in1(tmp03_3_23), .out(tmp04_1_23));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003035(.in0(tmp03_4_23), .in1(tmp03_5_23), .out(tmp04_2_23));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003036(.in0(tmp03_6_23), .in1(tmp03_7_23), .out(tmp04_3_23));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003037(.in0(tmp03_8_23), .in1(tmp03_9_23), .out(tmp04_4_23));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003038(.in0(tmp03_10_23), .in1(tmp03_11_23), .out(tmp04_5_23));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003039(.in0(tmp03_12_23), .in1(tmp03_13_23), .out(tmp04_6_23));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003040(.in0(tmp03_14_23), .in1(tmp03_15_23), .out(tmp04_7_23));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003041(.in0(tmp04_0_23), .in1(tmp04_1_23), .out(tmp05_0_23));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003042(.in0(tmp04_2_23), .in1(tmp04_3_23), .out(tmp05_1_23));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003043(.in0(tmp04_4_23), .in1(tmp04_5_23), .out(tmp05_2_23));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003044(.in0(tmp04_6_23), .in1(tmp04_7_23), .out(tmp05_3_23));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003045(.in0(tmp05_0_23), .in1(tmp05_1_23), .out(tmp06_0_23));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003046(.in0(tmp05_2_23), .in1(tmp05_3_23), .out(tmp06_1_23));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add003047(.in0(tmp06_0_23), .in1(tmp06_1_23), .out(tmp07_0_23));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003048(.in0(tmp00_0_24), .in1(tmp00_1_24), .out(tmp01_0_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003049(.in0(tmp00_2_24), .in1(tmp00_3_24), .out(tmp01_1_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003050(.in0(tmp00_4_24), .in1(tmp00_5_24), .out(tmp01_2_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003051(.in0(tmp00_6_24), .in1(tmp00_7_24), .out(tmp01_3_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003052(.in0(tmp00_8_24), .in1(tmp00_9_24), .out(tmp01_4_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003053(.in0(tmp00_10_24), .in1(tmp00_11_24), .out(tmp01_5_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003054(.in0(tmp00_12_24), .in1(tmp00_13_24), .out(tmp01_6_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003055(.in0(tmp00_14_24), .in1(tmp00_15_24), .out(tmp01_7_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003056(.in0(tmp00_16_24), .in1(tmp00_17_24), .out(tmp01_8_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003057(.in0(tmp00_18_24), .in1(tmp00_19_24), .out(tmp01_9_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003058(.in0(tmp00_20_24), .in1(tmp00_21_24), .out(tmp01_10_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003059(.in0(tmp00_22_24), .in1(tmp00_23_24), .out(tmp01_11_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003060(.in0(tmp00_24_24), .in1(tmp00_25_24), .out(tmp01_12_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003061(.in0(tmp00_26_24), .in1(tmp00_27_24), .out(tmp01_13_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003062(.in0(tmp00_28_24), .in1(tmp00_29_24), .out(tmp01_14_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003063(.in0(tmp00_30_24), .in1(tmp00_31_24), .out(tmp01_15_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003064(.in0(tmp00_32_24), .in1(tmp00_33_24), .out(tmp01_16_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003065(.in0(tmp00_34_24), .in1(tmp00_35_24), .out(tmp01_17_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003066(.in0(tmp00_36_24), .in1(tmp00_37_24), .out(tmp01_18_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003067(.in0(tmp00_38_24), .in1(tmp00_39_24), .out(tmp01_19_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003068(.in0(tmp00_40_24), .in1(tmp00_41_24), .out(tmp01_20_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003069(.in0(tmp00_42_24), .in1(tmp00_43_24), .out(tmp01_21_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003070(.in0(tmp00_44_24), .in1(tmp00_45_24), .out(tmp01_22_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003071(.in0(tmp00_46_24), .in1(tmp00_47_24), .out(tmp01_23_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003072(.in0(tmp00_48_24), .in1(tmp00_49_24), .out(tmp01_24_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003073(.in0(tmp00_50_24), .in1(tmp00_51_24), .out(tmp01_25_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003074(.in0(tmp00_52_24), .in1(tmp00_53_24), .out(tmp01_26_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003075(.in0(tmp00_54_24), .in1(tmp00_55_24), .out(tmp01_27_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003076(.in0(tmp00_56_24), .in1(tmp00_57_24), .out(tmp01_28_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003077(.in0(tmp00_58_24), .in1(tmp00_59_24), .out(tmp01_29_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003078(.in0(tmp00_60_24), .in1(tmp00_61_24), .out(tmp01_30_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003079(.in0(tmp00_62_24), .in1(tmp00_63_24), .out(tmp01_31_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003080(.in0(tmp00_64_24), .in1(tmp00_65_24), .out(tmp01_32_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003081(.in0(tmp00_66_24), .in1(tmp00_67_24), .out(tmp01_33_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003082(.in0(tmp00_68_24), .in1(tmp00_69_24), .out(tmp01_34_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003083(.in0(tmp00_70_24), .in1(tmp00_71_24), .out(tmp01_35_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003084(.in0(tmp00_72_24), .in1(tmp00_73_24), .out(tmp01_36_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003085(.in0(tmp00_74_24), .in1(tmp00_75_24), .out(tmp01_37_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003086(.in0(tmp00_76_24), .in1(tmp00_77_24), .out(tmp01_38_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003087(.in0(tmp00_78_24), .in1(tmp00_79_24), .out(tmp01_39_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003088(.in0(tmp00_80_24), .in1(tmp00_81_24), .out(tmp01_40_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003089(.in0(tmp00_82_24), .in1(tmp00_83_24), .out(tmp01_41_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003090(.in0(tmp00_84_24), .in1(tmp00_85_24), .out(tmp01_42_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003091(.in0(tmp00_86_24), .in1(tmp00_87_24), .out(tmp01_43_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003092(.in0(tmp00_88_24), .in1(tmp00_89_24), .out(tmp01_44_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003093(.in0(tmp00_90_24), .in1(tmp00_91_24), .out(tmp01_45_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003094(.in0(tmp00_92_24), .in1(tmp00_93_24), .out(tmp01_46_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003095(.in0(tmp00_94_24), .in1(tmp00_95_24), .out(tmp01_47_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003096(.in0(tmp00_96_24), .in1(tmp00_97_24), .out(tmp01_48_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003097(.in0(tmp00_98_24), .in1(tmp00_99_24), .out(tmp01_49_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003098(.in0(tmp00_100_24), .in1(tmp00_101_24), .out(tmp01_50_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003099(.in0(tmp00_102_24), .in1(tmp00_103_24), .out(tmp01_51_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003100(.in0(tmp00_104_24), .in1(tmp00_105_24), .out(tmp01_52_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003101(.in0(tmp00_106_24), .in1(tmp00_107_24), .out(tmp01_53_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003102(.in0(tmp00_108_24), .in1(tmp00_109_24), .out(tmp01_54_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003103(.in0(tmp00_110_24), .in1(tmp00_111_24), .out(tmp01_55_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003104(.in0(tmp00_112_24), .in1(tmp00_113_24), .out(tmp01_56_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003105(.in0(tmp00_114_24), .in1(tmp00_115_24), .out(tmp01_57_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003106(.in0(tmp00_116_24), .in1(tmp00_117_24), .out(tmp01_58_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003107(.in0(tmp00_118_24), .in1(tmp00_119_24), .out(tmp01_59_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003108(.in0(tmp00_120_24), .in1(tmp00_121_24), .out(tmp01_60_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003109(.in0(tmp00_122_24), .in1(tmp00_123_24), .out(tmp01_61_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003110(.in0(tmp00_124_24), .in1(tmp00_125_24), .out(tmp01_62_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003111(.in0(tmp00_126_24), .in1(tmp00_127_24), .out(tmp01_63_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003112(.in0(tmp01_0_24), .in1(tmp01_1_24), .out(tmp02_0_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003113(.in0(tmp01_2_24), .in1(tmp01_3_24), .out(tmp02_1_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003114(.in0(tmp01_4_24), .in1(tmp01_5_24), .out(tmp02_2_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003115(.in0(tmp01_6_24), .in1(tmp01_7_24), .out(tmp02_3_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003116(.in0(tmp01_8_24), .in1(tmp01_9_24), .out(tmp02_4_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003117(.in0(tmp01_10_24), .in1(tmp01_11_24), .out(tmp02_5_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003118(.in0(tmp01_12_24), .in1(tmp01_13_24), .out(tmp02_6_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003119(.in0(tmp01_14_24), .in1(tmp01_15_24), .out(tmp02_7_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003120(.in0(tmp01_16_24), .in1(tmp01_17_24), .out(tmp02_8_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003121(.in0(tmp01_18_24), .in1(tmp01_19_24), .out(tmp02_9_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003122(.in0(tmp01_20_24), .in1(tmp01_21_24), .out(tmp02_10_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003123(.in0(tmp01_22_24), .in1(tmp01_23_24), .out(tmp02_11_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003124(.in0(tmp01_24_24), .in1(tmp01_25_24), .out(tmp02_12_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003125(.in0(tmp01_26_24), .in1(tmp01_27_24), .out(tmp02_13_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003126(.in0(tmp01_28_24), .in1(tmp01_29_24), .out(tmp02_14_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003127(.in0(tmp01_30_24), .in1(tmp01_31_24), .out(tmp02_15_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003128(.in0(tmp01_32_24), .in1(tmp01_33_24), .out(tmp02_16_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003129(.in0(tmp01_34_24), .in1(tmp01_35_24), .out(tmp02_17_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003130(.in0(tmp01_36_24), .in1(tmp01_37_24), .out(tmp02_18_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003131(.in0(tmp01_38_24), .in1(tmp01_39_24), .out(tmp02_19_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003132(.in0(tmp01_40_24), .in1(tmp01_41_24), .out(tmp02_20_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003133(.in0(tmp01_42_24), .in1(tmp01_43_24), .out(tmp02_21_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003134(.in0(tmp01_44_24), .in1(tmp01_45_24), .out(tmp02_22_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003135(.in0(tmp01_46_24), .in1(tmp01_47_24), .out(tmp02_23_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003136(.in0(tmp01_48_24), .in1(tmp01_49_24), .out(tmp02_24_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003137(.in0(tmp01_50_24), .in1(tmp01_51_24), .out(tmp02_25_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003138(.in0(tmp01_52_24), .in1(tmp01_53_24), .out(tmp02_26_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003139(.in0(tmp01_54_24), .in1(tmp01_55_24), .out(tmp02_27_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003140(.in0(tmp01_56_24), .in1(tmp01_57_24), .out(tmp02_28_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003141(.in0(tmp01_58_24), .in1(tmp01_59_24), .out(tmp02_29_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003142(.in0(tmp01_60_24), .in1(tmp01_61_24), .out(tmp02_30_24));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003143(.in0(tmp01_62_24), .in1(tmp01_63_24), .out(tmp02_31_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003144(.in0(tmp02_0_24), .in1(tmp02_1_24), .out(tmp03_0_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003145(.in0(tmp02_2_24), .in1(tmp02_3_24), .out(tmp03_1_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003146(.in0(tmp02_4_24), .in1(tmp02_5_24), .out(tmp03_2_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003147(.in0(tmp02_6_24), .in1(tmp02_7_24), .out(tmp03_3_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003148(.in0(tmp02_8_24), .in1(tmp02_9_24), .out(tmp03_4_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003149(.in0(tmp02_10_24), .in1(tmp02_11_24), .out(tmp03_5_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003150(.in0(tmp02_12_24), .in1(tmp02_13_24), .out(tmp03_6_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003151(.in0(tmp02_14_24), .in1(tmp02_15_24), .out(tmp03_7_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003152(.in0(tmp02_16_24), .in1(tmp02_17_24), .out(tmp03_8_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003153(.in0(tmp02_18_24), .in1(tmp02_19_24), .out(tmp03_9_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003154(.in0(tmp02_20_24), .in1(tmp02_21_24), .out(tmp03_10_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003155(.in0(tmp02_22_24), .in1(tmp02_23_24), .out(tmp03_11_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003156(.in0(tmp02_24_24), .in1(tmp02_25_24), .out(tmp03_12_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003157(.in0(tmp02_26_24), .in1(tmp02_27_24), .out(tmp03_13_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003158(.in0(tmp02_28_24), .in1(tmp02_29_24), .out(tmp03_14_24));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003159(.in0(tmp02_30_24), .in1(tmp02_31_24), .out(tmp03_15_24));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003160(.in0(tmp03_0_24), .in1(tmp03_1_24), .out(tmp04_0_24));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003161(.in0(tmp03_2_24), .in1(tmp03_3_24), .out(tmp04_1_24));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003162(.in0(tmp03_4_24), .in1(tmp03_5_24), .out(tmp04_2_24));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003163(.in0(tmp03_6_24), .in1(tmp03_7_24), .out(tmp04_3_24));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003164(.in0(tmp03_8_24), .in1(tmp03_9_24), .out(tmp04_4_24));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003165(.in0(tmp03_10_24), .in1(tmp03_11_24), .out(tmp04_5_24));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003166(.in0(tmp03_12_24), .in1(tmp03_13_24), .out(tmp04_6_24));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003167(.in0(tmp03_14_24), .in1(tmp03_15_24), .out(tmp04_7_24));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003168(.in0(tmp04_0_24), .in1(tmp04_1_24), .out(tmp05_0_24));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003169(.in0(tmp04_2_24), .in1(tmp04_3_24), .out(tmp05_1_24));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003170(.in0(tmp04_4_24), .in1(tmp04_5_24), .out(tmp05_2_24));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003171(.in0(tmp04_6_24), .in1(tmp04_7_24), .out(tmp05_3_24));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003172(.in0(tmp05_0_24), .in1(tmp05_1_24), .out(tmp06_0_24));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003173(.in0(tmp05_2_24), .in1(tmp05_3_24), .out(tmp06_1_24));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add003174(.in0(tmp06_0_24), .in1(tmp06_1_24), .out(tmp07_0_24));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003175(.in0(tmp00_0_25), .in1(tmp00_1_25), .out(tmp01_0_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003176(.in0(tmp00_2_25), .in1(tmp00_3_25), .out(tmp01_1_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003177(.in0(tmp00_4_25), .in1(tmp00_5_25), .out(tmp01_2_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003178(.in0(tmp00_6_25), .in1(tmp00_7_25), .out(tmp01_3_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003179(.in0(tmp00_8_25), .in1(tmp00_9_25), .out(tmp01_4_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003180(.in0(tmp00_10_25), .in1(tmp00_11_25), .out(tmp01_5_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003181(.in0(tmp00_12_25), .in1(tmp00_13_25), .out(tmp01_6_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003182(.in0(tmp00_14_25), .in1(tmp00_15_25), .out(tmp01_7_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003183(.in0(tmp00_16_25), .in1(tmp00_17_25), .out(tmp01_8_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003184(.in0(tmp00_18_25), .in1(tmp00_19_25), .out(tmp01_9_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003185(.in0(tmp00_20_25), .in1(tmp00_21_25), .out(tmp01_10_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003186(.in0(tmp00_22_25), .in1(tmp00_23_25), .out(tmp01_11_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003187(.in0(tmp00_24_25), .in1(tmp00_25_25), .out(tmp01_12_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003188(.in0(tmp00_26_25), .in1(tmp00_27_25), .out(tmp01_13_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003189(.in0(tmp00_28_25), .in1(tmp00_29_25), .out(tmp01_14_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003190(.in0(tmp00_30_25), .in1(tmp00_31_25), .out(tmp01_15_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003191(.in0(tmp00_32_25), .in1(tmp00_33_25), .out(tmp01_16_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003192(.in0(tmp00_34_25), .in1(tmp00_35_25), .out(tmp01_17_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003193(.in0(tmp00_36_25), .in1(tmp00_37_25), .out(tmp01_18_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003194(.in0(tmp00_38_25), .in1(tmp00_39_25), .out(tmp01_19_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003195(.in0(tmp00_40_25), .in1(tmp00_41_25), .out(tmp01_20_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003196(.in0(tmp00_42_25), .in1(tmp00_43_25), .out(tmp01_21_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003197(.in0(tmp00_44_25), .in1(tmp00_45_25), .out(tmp01_22_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003198(.in0(tmp00_46_25), .in1(tmp00_47_25), .out(tmp01_23_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003199(.in0(tmp00_48_25), .in1(tmp00_49_25), .out(tmp01_24_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003200(.in0(tmp00_50_25), .in1(tmp00_51_25), .out(tmp01_25_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003201(.in0(tmp00_52_25), .in1(tmp00_53_25), .out(tmp01_26_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003202(.in0(tmp00_54_25), .in1(tmp00_55_25), .out(tmp01_27_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003203(.in0(tmp00_56_25), .in1(tmp00_57_25), .out(tmp01_28_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003204(.in0(tmp00_58_25), .in1(tmp00_59_25), .out(tmp01_29_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003205(.in0(tmp00_60_25), .in1(tmp00_61_25), .out(tmp01_30_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003206(.in0(tmp00_62_25), .in1(tmp00_63_25), .out(tmp01_31_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003207(.in0(tmp00_64_25), .in1(tmp00_65_25), .out(tmp01_32_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003208(.in0(tmp00_66_25), .in1(tmp00_67_25), .out(tmp01_33_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003209(.in0(tmp00_68_25), .in1(tmp00_69_25), .out(tmp01_34_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003210(.in0(tmp00_70_25), .in1(tmp00_71_25), .out(tmp01_35_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003211(.in0(tmp00_72_25), .in1(tmp00_73_25), .out(tmp01_36_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003212(.in0(tmp00_74_25), .in1(tmp00_75_25), .out(tmp01_37_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003213(.in0(tmp00_76_25), .in1(tmp00_77_25), .out(tmp01_38_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003214(.in0(tmp00_78_25), .in1(tmp00_79_25), .out(tmp01_39_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003215(.in0(tmp00_80_25), .in1(tmp00_81_25), .out(tmp01_40_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003216(.in0(tmp00_82_25), .in1(tmp00_83_25), .out(tmp01_41_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003217(.in0(tmp00_84_25), .in1(tmp00_85_25), .out(tmp01_42_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003218(.in0(tmp00_86_25), .in1(tmp00_87_25), .out(tmp01_43_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003219(.in0(tmp00_88_25), .in1(tmp00_89_25), .out(tmp01_44_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003220(.in0(tmp00_90_25), .in1(tmp00_91_25), .out(tmp01_45_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003221(.in0(tmp00_92_25), .in1(tmp00_93_25), .out(tmp01_46_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003222(.in0(tmp00_94_25), .in1(tmp00_95_25), .out(tmp01_47_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003223(.in0(tmp00_96_25), .in1(tmp00_97_25), .out(tmp01_48_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003224(.in0(tmp00_98_25), .in1(tmp00_99_25), .out(tmp01_49_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003225(.in0(tmp00_100_25), .in1(tmp00_101_25), .out(tmp01_50_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003226(.in0(tmp00_102_25), .in1(tmp00_103_25), .out(tmp01_51_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003227(.in0(tmp00_104_25), .in1(tmp00_105_25), .out(tmp01_52_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003228(.in0(tmp00_106_25), .in1(tmp00_107_25), .out(tmp01_53_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003229(.in0(tmp00_108_25), .in1(tmp00_109_25), .out(tmp01_54_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003230(.in0(tmp00_110_25), .in1(tmp00_111_25), .out(tmp01_55_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003231(.in0(tmp00_112_25), .in1(tmp00_113_25), .out(tmp01_56_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003232(.in0(tmp00_114_25), .in1(tmp00_115_25), .out(tmp01_57_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003233(.in0(tmp00_116_25), .in1(tmp00_117_25), .out(tmp01_58_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003234(.in0(tmp00_118_25), .in1(tmp00_119_25), .out(tmp01_59_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003235(.in0(tmp00_120_25), .in1(tmp00_121_25), .out(tmp01_60_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003236(.in0(tmp00_122_25), .in1(tmp00_123_25), .out(tmp01_61_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003237(.in0(tmp00_124_25), .in1(tmp00_125_25), .out(tmp01_62_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003238(.in0(tmp00_126_25), .in1(tmp00_127_25), .out(tmp01_63_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003239(.in0(tmp01_0_25), .in1(tmp01_1_25), .out(tmp02_0_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003240(.in0(tmp01_2_25), .in1(tmp01_3_25), .out(tmp02_1_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003241(.in0(tmp01_4_25), .in1(tmp01_5_25), .out(tmp02_2_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003242(.in0(tmp01_6_25), .in1(tmp01_7_25), .out(tmp02_3_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003243(.in0(tmp01_8_25), .in1(tmp01_9_25), .out(tmp02_4_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003244(.in0(tmp01_10_25), .in1(tmp01_11_25), .out(tmp02_5_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003245(.in0(tmp01_12_25), .in1(tmp01_13_25), .out(tmp02_6_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003246(.in0(tmp01_14_25), .in1(tmp01_15_25), .out(tmp02_7_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003247(.in0(tmp01_16_25), .in1(tmp01_17_25), .out(tmp02_8_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003248(.in0(tmp01_18_25), .in1(tmp01_19_25), .out(tmp02_9_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003249(.in0(tmp01_20_25), .in1(tmp01_21_25), .out(tmp02_10_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003250(.in0(tmp01_22_25), .in1(tmp01_23_25), .out(tmp02_11_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003251(.in0(tmp01_24_25), .in1(tmp01_25_25), .out(tmp02_12_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003252(.in0(tmp01_26_25), .in1(tmp01_27_25), .out(tmp02_13_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003253(.in0(tmp01_28_25), .in1(tmp01_29_25), .out(tmp02_14_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003254(.in0(tmp01_30_25), .in1(tmp01_31_25), .out(tmp02_15_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003255(.in0(tmp01_32_25), .in1(tmp01_33_25), .out(tmp02_16_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003256(.in0(tmp01_34_25), .in1(tmp01_35_25), .out(tmp02_17_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003257(.in0(tmp01_36_25), .in1(tmp01_37_25), .out(tmp02_18_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003258(.in0(tmp01_38_25), .in1(tmp01_39_25), .out(tmp02_19_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003259(.in0(tmp01_40_25), .in1(tmp01_41_25), .out(tmp02_20_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003260(.in0(tmp01_42_25), .in1(tmp01_43_25), .out(tmp02_21_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003261(.in0(tmp01_44_25), .in1(tmp01_45_25), .out(tmp02_22_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003262(.in0(tmp01_46_25), .in1(tmp01_47_25), .out(tmp02_23_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003263(.in0(tmp01_48_25), .in1(tmp01_49_25), .out(tmp02_24_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003264(.in0(tmp01_50_25), .in1(tmp01_51_25), .out(tmp02_25_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003265(.in0(tmp01_52_25), .in1(tmp01_53_25), .out(tmp02_26_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003266(.in0(tmp01_54_25), .in1(tmp01_55_25), .out(tmp02_27_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003267(.in0(tmp01_56_25), .in1(tmp01_57_25), .out(tmp02_28_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003268(.in0(tmp01_58_25), .in1(tmp01_59_25), .out(tmp02_29_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003269(.in0(tmp01_60_25), .in1(tmp01_61_25), .out(tmp02_30_25));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003270(.in0(tmp01_62_25), .in1(tmp01_63_25), .out(tmp02_31_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003271(.in0(tmp02_0_25), .in1(tmp02_1_25), .out(tmp03_0_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003272(.in0(tmp02_2_25), .in1(tmp02_3_25), .out(tmp03_1_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003273(.in0(tmp02_4_25), .in1(tmp02_5_25), .out(tmp03_2_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003274(.in0(tmp02_6_25), .in1(tmp02_7_25), .out(tmp03_3_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003275(.in0(tmp02_8_25), .in1(tmp02_9_25), .out(tmp03_4_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003276(.in0(tmp02_10_25), .in1(tmp02_11_25), .out(tmp03_5_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003277(.in0(tmp02_12_25), .in1(tmp02_13_25), .out(tmp03_6_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003278(.in0(tmp02_14_25), .in1(tmp02_15_25), .out(tmp03_7_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003279(.in0(tmp02_16_25), .in1(tmp02_17_25), .out(tmp03_8_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003280(.in0(tmp02_18_25), .in1(tmp02_19_25), .out(tmp03_9_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003281(.in0(tmp02_20_25), .in1(tmp02_21_25), .out(tmp03_10_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003282(.in0(tmp02_22_25), .in1(tmp02_23_25), .out(tmp03_11_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003283(.in0(tmp02_24_25), .in1(tmp02_25_25), .out(tmp03_12_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003284(.in0(tmp02_26_25), .in1(tmp02_27_25), .out(tmp03_13_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003285(.in0(tmp02_28_25), .in1(tmp02_29_25), .out(tmp03_14_25));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003286(.in0(tmp02_30_25), .in1(tmp02_31_25), .out(tmp03_15_25));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003287(.in0(tmp03_0_25), .in1(tmp03_1_25), .out(tmp04_0_25));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003288(.in0(tmp03_2_25), .in1(tmp03_3_25), .out(tmp04_1_25));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003289(.in0(tmp03_4_25), .in1(tmp03_5_25), .out(tmp04_2_25));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003290(.in0(tmp03_6_25), .in1(tmp03_7_25), .out(tmp04_3_25));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003291(.in0(tmp03_8_25), .in1(tmp03_9_25), .out(tmp04_4_25));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003292(.in0(tmp03_10_25), .in1(tmp03_11_25), .out(tmp04_5_25));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003293(.in0(tmp03_12_25), .in1(tmp03_13_25), .out(tmp04_6_25));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003294(.in0(tmp03_14_25), .in1(tmp03_15_25), .out(tmp04_7_25));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003295(.in0(tmp04_0_25), .in1(tmp04_1_25), .out(tmp05_0_25));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003296(.in0(tmp04_2_25), .in1(tmp04_3_25), .out(tmp05_1_25));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003297(.in0(tmp04_4_25), .in1(tmp04_5_25), .out(tmp05_2_25));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003298(.in0(tmp04_6_25), .in1(tmp04_7_25), .out(tmp05_3_25));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003299(.in0(tmp05_0_25), .in1(tmp05_1_25), .out(tmp06_0_25));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003300(.in0(tmp05_2_25), .in1(tmp05_3_25), .out(tmp06_1_25));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add003301(.in0(tmp06_0_25), .in1(tmp06_1_25), .out(tmp07_0_25));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003302(.in0(tmp00_0_26), .in1(tmp00_1_26), .out(tmp01_0_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003303(.in0(tmp00_2_26), .in1(tmp00_3_26), .out(tmp01_1_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003304(.in0(tmp00_4_26), .in1(tmp00_5_26), .out(tmp01_2_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003305(.in0(tmp00_6_26), .in1(tmp00_7_26), .out(tmp01_3_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003306(.in0(tmp00_8_26), .in1(tmp00_9_26), .out(tmp01_4_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003307(.in0(tmp00_10_26), .in1(tmp00_11_26), .out(tmp01_5_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003308(.in0(tmp00_12_26), .in1(tmp00_13_26), .out(tmp01_6_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003309(.in0(tmp00_14_26), .in1(tmp00_15_26), .out(tmp01_7_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003310(.in0(tmp00_16_26), .in1(tmp00_17_26), .out(tmp01_8_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003311(.in0(tmp00_18_26), .in1(tmp00_19_26), .out(tmp01_9_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003312(.in0(tmp00_20_26), .in1(tmp00_21_26), .out(tmp01_10_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003313(.in0(tmp00_22_26), .in1(tmp00_23_26), .out(tmp01_11_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003314(.in0(tmp00_24_26), .in1(tmp00_25_26), .out(tmp01_12_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003315(.in0(tmp00_26_26), .in1(tmp00_27_26), .out(tmp01_13_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003316(.in0(tmp00_28_26), .in1(tmp00_29_26), .out(tmp01_14_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003317(.in0(tmp00_30_26), .in1(tmp00_31_26), .out(tmp01_15_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003318(.in0(tmp00_32_26), .in1(tmp00_33_26), .out(tmp01_16_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003319(.in0(tmp00_34_26), .in1(tmp00_35_26), .out(tmp01_17_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003320(.in0(tmp00_36_26), .in1(tmp00_37_26), .out(tmp01_18_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003321(.in0(tmp00_38_26), .in1(tmp00_39_26), .out(tmp01_19_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003322(.in0(tmp00_40_26), .in1(tmp00_41_26), .out(tmp01_20_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003323(.in0(tmp00_42_26), .in1(tmp00_43_26), .out(tmp01_21_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003324(.in0(tmp00_44_26), .in1(tmp00_45_26), .out(tmp01_22_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003325(.in0(tmp00_46_26), .in1(tmp00_47_26), .out(tmp01_23_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003326(.in0(tmp00_48_26), .in1(tmp00_49_26), .out(tmp01_24_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003327(.in0(tmp00_50_26), .in1(tmp00_51_26), .out(tmp01_25_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003328(.in0(tmp00_52_26), .in1(tmp00_53_26), .out(tmp01_26_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003329(.in0(tmp00_54_26), .in1(tmp00_55_26), .out(tmp01_27_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003330(.in0(tmp00_56_26), .in1(tmp00_57_26), .out(tmp01_28_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003331(.in0(tmp00_58_26), .in1(tmp00_59_26), .out(tmp01_29_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003332(.in0(tmp00_60_26), .in1(tmp00_61_26), .out(tmp01_30_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003333(.in0(tmp00_62_26), .in1(tmp00_63_26), .out(tmp01_31_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003334(.in0(tmp00_64_26), .in1(tmp00_65_26), .out(tmp01_32_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003335(.in0(tmp00_66_26), .in1(tmp00_67_26), .out(tmp01_33_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003336(.in0(tmp00_68_26), .in1(tmp00_69_26), .out(tmp01_34_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003337(.in0(tmp00_70_26), .in1(tmp00_71_26), .out(tmp01_35_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003338(.in0(tmp00_72_26), .in1(tmp00_73_26), .out(tmp01_36_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003339(.in0(tmp00_74_26), .in1(tmp00_75_26), .out(tmp01_37_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003340(.in0(tmp00_76_26), .in1(tmp00_77_26), .out(tmp01_38_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003341(.in0(tmp00_78_26), .in1(tmp00_79_26), .out(tmp01_39_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003342(.in0(tmp00_80_26), .in1(tmp00_81_26), .out(tmp01_40_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003343(.in0(tmp00_82_26), .in1(tmp00_83_26), .out(tmp01_41_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003344(.in0(tmp00_84_26), .in1(tmp00_85_26), .out(tmp01_42_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003345(.in0(tmp00_86_26), .in1(tmp00_87_26), .out(tmp01_43_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003346(.in0(tmp00_88_26), .in1(tmp00_89_26), .out(tmp01_44_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003347(.in0(tmp00_90_26), .in1(tmp00_91_26), .out(tmp01_45_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003348(.in0(tmp00_92_26), .in1(tmp00_93_26), .out(tmp01_46_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003349(.in0(tmp00_94_26), .in1(tmp00_95_26), .out(tmp01_47_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003350(.in0(tmp00_96_26), .in1(tmp00_97_26), .out(tmp01_48_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003351(.in0(tmp00_98_26), .in1(tmp00_99_26), .out(tmp01_49_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003352(.in0(tmp00_100_26), .in1(tmp00_101_26), .out(tmp01_50_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003353(.in0(tmp00_102_26), .in1(tmp00_103_26), .out(tmp01_51_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003354(.in0(tmp00_104_26), .in1(tmp00_105_26), .out(tmp01_52_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003355(.in0(tmp00_106_26), .in1(tmp00_107_26), .out(tmp01_53_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003356(.in0(tmp00_108_26), .in1(tmp00_109_26), .out(tmp01_54_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003357(.in0(tmp00_110_26), .in1(tmp00_111_26), .out(tmp01_55_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003358(.in0(tmp00_112_26), .in1(tmp00_113_26), .out(tmp01_56_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003359(.in0(tmp00_114_26), .in1(tmp00_115_26), .out(tmp01_57_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003360(.in0(tmp00_116_26), .in1(tmp00_117_26), .out(tmp01_58_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003361(.in0(tmp00_118_26), .in1(tmp00_119_26), .out(tmp01_59_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003362(.in0(tmp00_120_26), .in1(tmp00_121_26), .out(tmp01_60_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003363(.in0(tmp00_122_26), .in1(tmp00_123_26), .out(tmp01_61_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003364(.in0(tmp00_124_26), .in1(tmp00_125_26), .out(tmp01_62_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003365(.in0(tmp00_126_26), .in1(tmp00_127_26), .out(tmp01_63_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003366(.in0(tmp01_0_26), .in1(tmp01_1_26), .out(tmp02_0_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003367(.in0(tmp01_2_26), .in1(tmp01_3_26), .out(tmp02_1_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003368(.in0(tmp01_4_26), .in1(tmp01_5_26), .out(tmp02_2_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003369(.in0(tmp01_6_26), .in1(tmp01_7_26), .out(tmp02_3_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003370(.in0(tmp01_8_26), .in1(tmp01_9_26), .out(tmp02_4_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003371(.in0(tmp01_10_26), .in1(tmp01_11_26), .out(tmp02_5_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003372(.in0(tmp01_12_26), .in1(tmp01_13_26), .out(tmp02_6_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003373(.in0(tmp01_14_26), .in1(tmp01_15_26), .out(tmp02_7_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003374(.in0(tmp01_16_26), .in1(tmp01_17_26), .out(tmp02_8_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003375(.in0(tmp01_18_26), .in1(tmp01_19_26), .out(tmp02_9_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003376(.in0(tmp01_20_26), .in1(tmp01_21_26), .out(tmp02_10_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003377(.in0(tmp01_22_26), .in1(tmp01_23_26), .out(tmp02_11_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003378(.in0(tmp01_24_26), .in1(tmp01_25_26), .out(tmp02_12_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003379(.in0(tmp01_26_26), .in1(tmp01_27_26), .out(tmp02_13_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003380(.in0(tmp01_28_26), .in1(tmp01_29_26), .out(tmp02_14_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003381(.in0(tmp01_30_26), .in1(tmp01_31_26), .out(tmp02_15_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003382(.in0(tmp01_32_26), .in1(tmp01_33_26), .out(tmp02_16_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003383(.in0(tmp01_34_26), .in1(tmp01_35_26), .out(tmp02_17_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003384(.in0(tmp01_36_26), .in1(tmp01_37_26), .out(tmp02_18_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003385(.in0(tmp01_38_26), .in1(tmp01_39_26), .out(tmp02_19_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003386(.in0(tmp01_40_26), .in1(tmp01_41_26), .out(tmp02_20_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003387(.in0(tmp01_42_26), .in1(tmp01_43_26), .out(tmp02_21_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003388(.in0(tmp01_44_26), .in1(tmp01_45_26), .out(tmp02_22_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003389(.in0(tmp01_46_26), .in1(tmp01_47_26), .out(tmp02_23_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003390(.in0(tmp01_48_26), .in1(tmp01_49_26), .out(tmp02_24_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003391(.in0(tmp01_50_26), .in1(tmp01_51_26), .out(tmp02_25_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003392(.in0(tmp01_52_26), .in1(tmp01_53_26), .out(tmp02_26_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003393(.in0(tmp01_54_26), .in1(tmp01_55_26), .out(tmp02_27_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003394(.in0(tmp01_56_26), .in1(tmp01_57_26), .out(tmp02_28_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003395(.in0(tmp01_58_26), .in1(tmp01_59_26), .out(tmp02_29_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003396(.in0(tmp01_60_26), .in1(tmp01_61_26), .out(tmp02_30_26));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003397(.in0(tmp01_62_26), .in1(tmp01_63_26), .out(tmp02_31_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003398(.in0(tmp02_0_26), .in1(tmp02_1_26), .out(tmp03_0_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003399(.in0(tmp02_2_26), .in1(tmp02_3_26), .out(tmp03_1_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003400(.in0(tmp02_4_26), .in1(tmp02_5_26), .out(tmp03_2_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003401(.in0(tmp02_6_26), .in1(tmp02_7_26), .out(tmp03_3_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003402(.in0(tmp02_8_26), .in1(tmp02_9_26), .out(tmp03_4_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003403(.in0(tmp02_10_26), .in1(tmp02_11_26), .out(tmp03_5_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003404(.in0(tmp02_12_26), .in1(tmp02_13_26), .out(tmp03_6_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003405(.in0(tmp02_14_26), .in1(tmp02_15_26), .out(tmp03_7_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003406(.in0(tmp02_16_26), .in1(tmp02_17_26), .out(tmp03_8_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003407(.in0(tmp02_18_26), .in1(tmp02_19_26), .out(tmp03_9_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003408(.in0(tmp02_20_26), .in1(tmp02_21_26), .out(tmp03_10_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003409(.in0(tmp02_22_26), .in1(tmp02_23_26), .out(tmp03_11_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003410(.in0(tmp02_24_26), .in1(tmp02_25_26), .out(tmp03_12_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003411(.in0(tmp02_26_26), .in1(tmp02_27_26), .out(tmp03_13_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003412(.in0(tmp02_28_26), .in1(tmp02_29_26), .out(tmp03_14_26));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003413(.in0(tmp02_30_26), .in1(tmp02_31_26), .out(tmp03_15_26));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003414(.in0(tmp03_0_26), .in1(tmp03_1_26), .out(tmp04_0_26));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003415(.in0(tmp03_2_26), .in1(tmp03_3_26), .out(tmp04_1_26));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003416(.in0(tmp03_4_26), .in1(tmp03_5_26), .out(tmp04_2_26));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003417(.in0(tmp03_6_26), .in1(tmp03_7_26), .out(tmp04_3_26));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003418(.in0(tmp03_8_26), .in1(tmp03_9_26), .out(tmp04_4_26));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003419(.in0(tmp03_10_26), .in1(tmp03_11_26), .out(tmp04_5_26));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003420(.in0(tmp03_12_26), .in1(tmp03_13_26), .out(tmp04_6_26));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003421(.in0(tmp03_14_26), .in1(tmp03_15_26), .out(tmp04_7_26));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003422(.in0(tmp04_0_26), .in1(tmp04_1_26), .out(tmp05_0_26));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003423(.in0(tmp04_2_26), .in1(tmp04_3_26), .out(tmp05_1_26));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003424(.in0(tmp04_4_26), .in1(tmp04_5_26), .out(tmp05_2_26));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003425(.in0(tmp04_6_26), .in1(tmp04_7_26), .out(tmp05_3_26));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003426(.in0(tmp05_0_26), .in1(tmp05_1_26), .out(tmp06_0_26));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003427(.in0(tmp05_2_26), .in1(tmp05_3_26), .out(tmp06_1_26));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add003428(.in0(tmp06_0_26), .in1(tmp06_1_26), .out(tmp07_0_26));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003429(.in0(tmp00_0_27), .in1(tmp00_1_27), .out(tmp01_0_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003430(.in0(tmp00_2_27), .in1(tmp00_3_27), .out(tmp01_1_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003431(.in0(tmp00_4_27), .in1(tmp00_5_27), .out(tmp01_2_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003432(.in0(tmp00_6_27), .in1(tmp00_7_27), .out(tmp01_3_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003433(.in0(tmp00_8_27), .in1(tmp00_9_27), .out(tmp01_4_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003434(.in0(tmp00_10_27), .in1(tmp00_11_27), .out(tmp01_5_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003435(.in0(tmp00_12_27), .in1(tmp00_13_27), .out(tmp01_6_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003436(.in0(tmp00_14_27), .in1(tmp00_15_27), .out(tmp01_7_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003437(.in0(tmp00_16_27), .in1(tmp00_17_27), .out(tmp01_8_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003438(.in0(tmp00_18_27), .in1(tmp00_19_27), .out(tmp01_9_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003439(.in0(tmp00_20_27), .in1(tmp00_21_27), .out(tmp01_10_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003440(.in0(tmp00_22_27), .in1(tmp00_23_27), .out(tmp01_11_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003441(.in0(tmp00_24_27), .in1(tmp00_25_27), .out(tmp01_12_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003442(.in0(tmp00_26_27), .in1(tmp00_27_27), .out(tmp01_13_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003443(.in0(tmp00_28_27), .in1(tmp00_29_27), .out(tmp01_14_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003444(.in0(tmp00_30_27), .in1(tmp00_31_27), .out(tmp01_15_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003445(.in0(tmp00_32_27), .in1(tmp00_33_27), .out(tmp01_16_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003446(.in0(tmp00_34_27), .in1(tmp00_35_27), .out(tmp01_17_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003447(.in0(tmp00_36_27), .in1(tmp00_37_27), .out(tmp01_18_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003448(.in0(tmp00_38_27), .in1(tmp00_39_27), .out(tmp01_19_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003449(.in0(tmp00_40_27), .in1(tmp00_41_27), .out(tmp01_20_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003450(.in0(tmp00_42_27), .in1(tmp00_43_27), .out(tmp01_21_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003451(.in0(tmp00_44_27), .in1(tmp00_45_27), .out(tmp01_22_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003452(.in0(tmp00_46_27), .in1(tmp00_47_27), .out(tmp01_23_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003453(.in0(tmp00_48_27), .in1(tmp00_49_27), .out(tmp01_24_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003454(.in0(tmp00_50_27), .in1(tmp00_51_27), .out(tmp01_25_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003455(.in0(tmp00_52_27), .in1(tmp00_53_27), .out(tmp01_26_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003456(.in0(tmp00_54_27), .in1(tmp00_55_27), .out(tmp01_27_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003457(.in0(tmp00_56_27), .in1(tmp00_57_27), .out(tmp01_28_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003458(.in0(tmp00_58_27), .in1(tmp00_59_27), .out(tmp01_29_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003459(.in0(tmp00_60_27), .in1(tmp00_61_27), .out(tmp01_30_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003460(.in0(tmp00_62_27), .in1(tmp00_63_27), .out(tmp01_31_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003461(.in0(tmp00_64_27), .in1(tmp00_65_27), .out(tmp01_32_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003462(.in0(tmp00_66_27), .in1(tmp00_67_27), .out(tmp01_33_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003463(.in0(tmp00_68_27), .in1(tmp00_69_27), .out(tmp01_34_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003464(.in0(tmp00_70_27), .in1(tmp00_71_27), .out(tmp01_35_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003465(.in0(tmp00_72_27), .in1(tmp00_73_27), .out(tmp01_36_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003466(.in0(tmp00_74_27), .in1(tmp00_75_27), .out(tmp01_37_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003467(.in0(tmp00_76_27), .in1(tmp00_77_27), .out(tmp01_38_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003468(.in0(tmp00_78_27), .in1(tmp00_79_27), .out(tmp01_39_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003469(.in0(tmp00_80_27), .in1(tmp00_81_27), .out(tmp01_40_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003470(.in0(tmp00_82_27), .in1(tmp00_83_27), .out(tmp01_41_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003471(.in0(tmp00_84_27), .in1(tmp00_85_27), .out(tmp01_42_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003472(.in0(tmp00_86_27), .in1(tmp00_87_27), .out(tmp01_43_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003473(.in0(tmp00_88_27), .in1(tmp00_89_27), .out(tmp01_44_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003474(.in0(tmp00_90_27), .in1(tmp00_91_27), .out(tmp01_45_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003475(.in0(tmp00_92_27), .in1(tmp00_93_27), .out(tmp01_46_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003476(.in0(tmp00_94_27), .in1(tmp00_95_27), .out(tmp01_47_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003477(.in0(tmp00_96_27), .in1(tmp00_97_27), .out(tmp01_48_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003478(.in0(tmp00_98_27), .in1(tmp00_99_27), .out(tmp01_49_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003479(.in0(tmp00_100_27), .in1(tmp00_101_27), .out(tmp01_50_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003480(.in0(tmp00_102_27), .in1(tmp00_103_27), .out(tmp01_51_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003481(.in0(tmp00_104_27), .in1(tmp00_105_27), .out(tmp01_52_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003482(.in0(tmp00_106_27), .in1(tmp00_107_27), .out(tmp01_53_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003483(.in0(tmp00_108_27), .in1(tmp00_109_27), .out(tmp01_54_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003484(.in0(tmp00_110_27), .in1(tmp00_111_27), .out(tmp01_55_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003485(.in0(tmp00_112_27), .in1(tmp00_113_27), .out(tmp01_56_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003486(.in0(tmp00_114_27), .in1(tmp00_115_27), .out(tmp01_57_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003487(.in0(tmp00_116_27), .in1(tmp00_117_27), .out(tmp01_58_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003488(.in0(tmp00_118_27), .in1(tmp00_119_27), .out(tmp01_59_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003489(.in0(tmp00_120_27), .in1(tmp00_121_27), .out(tmp01_60_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003490(.in0(tmp00_122_27), .in1(tmp00_123_27), .out(tmp01_61_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003491(.in0(tmp00_124_27), .in1(tmp00_125_27), .out(tmp01_62_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003492(.in0(tmp00_126_27), .in1(tmp00_127_27), .out(tmp01_63_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003493(.in0(tmp01_0_27), .in1(tmp01_1_27), .out(tmp02_0_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003494(.in0(tmp01_2_27), .in1(tmp01_3_27), .out(tmp02_1_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003495(.in0(tmp01_4_27), .in1(tmp01_5_27), .out(tmp02_2_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003496(.in0(tmp01_6_27), .in1(tmp01_7_27), .out(tmp02_3_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003497(.in0(tmp01_8_27), .in1(tmp01_9_27), .out(tmp02_4_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003498(.in0(tmp01_10_27), .in1(tmp01_11_27), .out(tmp02_5_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003499(.in0(tmp01_12_27), .in1(tmp01_13_27), .out(tmp02_6_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003500(.in0(tmp01_14_27), .in1(tmp01_15_27), .out(tmp02_7_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003501(.in0(tmp01_16_27), .in1(tmp01_17_27), .out(tmp02_8_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003502(.in0(tmp01_18_27), .in1(tmp01_19_27), .out(tmp02_9_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003503(.in0(tmp01_20_27), .in1(tmp01_21_27), .out(tmp02_10_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003504(.in0(tmp01_22_27), .in1(tmp01_23_27), .out(tmp02_11_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003505(.in0(tmp01_24_27), .in1(tmp01_25_27), .out(tmp02_12_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003506(.in0(tmp01_26_27), .in1(tmp01_27_27), .out(tmp02_13_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003507(.in0(tmp01_28_27), .in1(tmp01_29_27), .out(tmp02_14_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003508(.in0(tmp01_30_27), .in1(tmp01_31_27), .out(tmp02_15_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003509(.in0(tmp01_32_27), .in1(tmp01_33_27), .out(tmp02_16_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003510(.in0(tmp01_34_27), .in1(tmp01_35_27), .out(tmp02_17_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003511(.in0(tmp01_36_27), .in1(tmp01_37_27), .out(tmp02_18_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003512(.in0(tmp01_38_27), .in1(tmp01_39_27), .out(tmp02_19_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003513(.in0(tmp01_40_27), .in1(tmp01_41_27), .out(tmp02_20_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003514(.in0(tmp01_42_27), .in1(tmp01_43_27), .out(tmp02_21_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003515(.in0(tmp01_44_27), .in1(tmp01_45_27), .out(tmp02_22_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003516(.in0(tmp01_46_27), .in1(tmp01_47_27), .out(tmp02_23_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003517(.in0(tmp01_48_27), .in1(tmp01_49_27), .out(tmp02_24_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003518(.in0(tmp01_50_27), .in1(tmp01_51_27), .out(tmp02_25_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003519(.in0(tmp01_52_27), .in1(tmp01_53_27), .out(tmp02_26_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003520(.in0(tmp01_54_27), .in1(tmp01_55_27), .out(tmp02_27_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003521(.in0(tmp01_56_27), .in1(tmp01_57_27), .out(tmp02_28_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003522(.in0(tmp01_58_27), .in1(tmp01_59_27), .out(tmp02_29_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003523(.in0(tmp01_60_27), .in1(tmp01_61_27), .out(tmp02_30_27));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003524(.in0(tmp01_62_27), .in1(tmp01_63_27), .out(tmp02_31_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003525(.in0(tmp02_0_27), .in1(tmp02_1_27), .out(tmp03_0_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003526(.in0(tmp02_2_27), .in1(tmp02_3_27), .out(tmp03_1_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003527(.in0(tmp02_4_27), .in1(tmp02_5_27), .out(tmp03_2_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003528(.in0(tmp02_6_27), .in1(tmp02_7_27), .out(tmp03_3_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003529(.in0(tmp02_8_27), .in1(tmp02_9_27), .out(tmp03_4_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003530(.in0(tmp02_10_27), .in1(tmp02_11_27), .out(tmp03_5_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003531(.in0(tmp02_12_27), .in1(tmp02_13_27), .out(tmp03_6_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003532(.in0(tmp02_14_27), .in1(tmp02_15_27), .out(tmp03_7_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003533(.in0(tmp02_16_27), .in1(tmp02_17_27), .out(tmp03_8_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003534(.in0(tmp02_18_27), .in1(tmp02_19_27), .out(tmp03_9_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003535(.in0(tmp02_20_27), .in1(tmp02_21_27), .out(tmp03_10_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003536(.in0(tmp02_22_27), .in1(tmp02_23_27), .out(tmp03_11_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003537(.in0(tmp02_24_27), .in1(tmp02_25_27), .out(tmp03_12_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003538(.in0(tmp02_26_27), .in1(tmp02_27_27), .out(tmp03_13_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003539(.in0(tmp02_28_27), .in1(tmp02_29_27), .out(tmp03_14_27));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003540(.in0(tmp02_30_27), .in1(tmp02_31_27), .out(tmp03_15_27));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003541(.in0(tmp03_0_27), .in1(tmp03_1_27), .out(tmp04_0_27));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003542(.in0(tmp03_2_27), .in1(tmp03_3_27), .out(tmp04_1_27));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003543(.in0(tmp03_4_27), .in1(tmp03_5_27), .out(tmp04_2_27));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003544(.in0(tmp03_6_27), .in1(tmp03_7_27), .out(tmp04_3_27));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003545(.in0(tmp03_8_27), .in1(tmp03_9_27), .out(tmp04_4_27));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003546(.in0(tmp03_10_27), .in1(tmp03_11_27), .out(tmp04_5_27));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003547(.in0(tmp03_12_27), .in1(tmp03_13_27), .out(tmp04_6_27));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003548(.in0(tmp03_14_27), .in1(tmp03_15_27), .out(tmp04_7_27));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003549(.in0(tmp04_0_27), .in1(tmp04_1_27), .out(tmp05_0_27));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003550(.in0(tmp04_2_27), .in1(tmp04_3_27), .out(tmp05_1_27));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003551(.in0(tmp04_4_27), .in1(tmp04_5_27), .out(tmp05_2_27));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003552(.in0(tmp04_6_27), .in1(tmp04_7_27), .out(tmp05_3_27));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003553(.in0(tmp05_0_27), .in1(tmp05_1_27), .out(tmp06_0_27));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003554(.in0(tmp05_2_27), .in1(tmp05_3_27), .out(tmp06_1_27));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add003555(.in0(tmp06_0_27), .in1(tmp06_1_27), .out(tmp07_0_27));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003556(.in0(tmp00_0_28), .in1(tmp00_1_28), .out(tmp01_0_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003557(.in0(tmp00_2_28), .in1(tmp00_3_28), .out(tmp01_1_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003558(.in0(tmp00_4_28), .in1(tmp00_5_28), .out(tmp01_2_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003559(.in0(tmp00_6_28), .in1(tmp00_7_28), .out(tmp01_3_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003560(.in0(tmp00_8_28), .in1(tmp00_9_28), .out(tmp01_4_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003561(.in0(tmp00_10_28), .in1(tmp00_11_28), .out(tmp01_5_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003562(.in0(tmp00_12_28), .in1(tmp00_13_28), .out(tmp01_6_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003563(.in0(tmp00_14_28), .in1(tmp00_15_28), .out(tmp01_7_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003564(.in0(tmp00_16_28), .in1(tmp00_17_28), .out(tmp01_8_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003565(.in0(tmp00_18_28), .in1(tmp00_19_28), .out(tmp01_9_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003566(.in0(tmp00_20_28), .in1(tmp00_21_28), .out(tmp01_10_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003567(.in0(tmp00_22_28), .in1(tmp00_23_28), .out(tmp01_11_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003568(.in0(tmp00_24_28), .in1(tmp00_25_28), .out(tmp01_12_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003569(.in0(tmp00_26_28), .in1(tmp00_27_28), .out(tmp01_13_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003570(.in0(tmp00_28_28), .in1(tmp00_29_28), .out(tmp01_14_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003571(.in0(tmp00_30_28), .in1(tmp00_31_28), .out(tmp01_15_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003572(.in0(tmp00_32_28), .in1(tmp00_33_28), .out(tmp01_16_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003573(.in0(tmp00_34_28), .in1(tmp00_35_28), .out(tmp01_17_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003574(.in0(tmp00_36_28), .in1(tmp00_37_28), .out(tmp01_18_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003575(.in0(tmp00_38_28), .in1(tmp00_39_28), .out(tmp01_19_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003576(.in0(tmp00_40_28), .in1(tmp00_41_28), .out(tmp01_20_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003577(.in0(tmp00_42_28), .in1(tmp00_43_28), .out(tmp01_21_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003578(.in0(tmp00_44_28), .in1(tmp00_45_28), .out(tmp01_22_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003579(.in0(tmp00_46_28), .in1(tmp00_47_28), .out(tmp01_23_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003580(.in0(tmp00_48_28), .in1(tmp00_49_28), .out(tmp01_24_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003581(.in0(tmp00_50_28), .in1(tmp00_51_28), .out(tmp01_25_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003582(.in0(tmp00_52_28), .in1(tmp00_53_28), .out(tmp01_26_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003583(.in0(tmp00_54_28), .in1(tmp00_55_28), .out(tmp01_27_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003584(.in0(tmp00_56_28), .in1(tmp00_57_28), .out(tmp01_28_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003585(.in0(tmp00_58_28), .in1(tmp00_59_28), .out(tmp01_29_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003586(.in0(tmp00_60_28), .in1(tmp00_61_28), .out(tmp01_30_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003587(.in0(tmp00_62_28), .in1(tmp00_63_28), .out(tmp01_31_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003588(.in0(tmp00_64_28), .in1(tmp00_65_28), .out(tmp01_32_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003589(.in0(tmp00_66_28), .in1(tmp00_67_28), .out(tmp01_33_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003590(.in0(tmp00_68_28), .in1(tmp00_69_28), .out(tmp01_34_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003591(.in0(tmp00_70_28), .in1(tmp00_71_28), .out(tmp01_35_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003592(.in0(tmp00_72_28), .in1(tmp00_73_28), .out(tmp01_36_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003593(.in0(tmp00_74_28), .in1(tmp00_75_28), .out(tmp01_37_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003594(.in0(tmp00_76_28), .in1(tmp00_77_28), .out(tmp01_38_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003595(.in0(tmp00_78_28), .in1(tmp00_79_28), .out(tmp01_39_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003596(.in0(tmp00_80_28), .in1(tmp00_81_28), .out(tmp01_40_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003597(.in0(tmp00_82_28), .in1(tmp00_83_28), .out(tmp01_41_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003598(.in0(tmp00_84_28), .in1(tmp00_85_28), .out(tmp01_42_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003599(.in0(tmp00_86_28), .in1(tmp00_87_28), .out(tmp01_43_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003600(.in0(tmp00_88_28), .in1(tmp00_89_28), .out(tmp01_44_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003601(.in0(tmp00_90_28), .in1(tmp00_91_28), .out(tmp01_45_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003602(.in0(tmp00_92_28), .in1(tmp00_93_28), .out(tmp01_46_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003603(.in0(tmp00_94_28), .in1(tmp00_95_28), .out(tmp01_47_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003604(.in0(tmp00_96_28), .in1(tmp00_97_28), .out(tmp01_48_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003605(.in0(tmp00_98_28), .in1(tmp00_99_28), .out(tmp01_49_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003606(.in0(tmp00_100_28), .in1(tmp00_101_28), .out(tmp01_50_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003607(.in0(tmp00_102_28), .in1(tmp00_103_28), .out(tmp01_51_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003608(.in0(tmp00_104_28), .in1(tmp00_105_28), .out(tmp01_52_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003609(.in0(tmp00_106_28), .in1(tmp00_107_28), .out(tmp01_53_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003610(.in0(tmp00_108_28), .in1(tmp00_109_28), .out(tmp01_54_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003611(.in0(tmp00_110_28), .in1(tmp00_111_28), .out(tmp01_55_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003612(.in0(tmp00_112_28), .in1(tmp00_113_28), .out(tmp01_56_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003613(.in0(tmp00_114_28), .in1(tmp00_115_28), .out(tmp01_57_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003614(.in0(tmp00_116_28), .in1(tmp00_117_28), .out(tmp01_58_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003615(.in0(tmp00_118_28), .in1(tmp00_119_28), .out(tmp01_59_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003616(.in0(tmp00_120_28), .in1(tmp00_121_28), .out(tmp01_60_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003617(.in0(tmp00_122_28), .in1(tmp00_123_28), .out(tmp01_61_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003618(.in0(tmp00_124_28), .in1(tmp00_125_28), .out(tmp01_62_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003619(.in0(tmp00_126_28), .in1(tmp00_127_28), .out(tmp01_63_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003620(.in0(tmp01_0_28), .in1(tmp01_1_28), .out(tmp02_0_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003621(.in0(tmp01_2_28), .in1(tmp01_3_28), .out(tmp02_1_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003622(.in0(tmp01_4_28), .in1(tmp01_5_28), .out(tmp02_2_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003623(.in0(tmp01_6_28), .in1(tmp01_7_28), .out(tmp02_3_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003624(.in0(tmp01_8_28), .in1(tmp01_9_28), .out(tmp02_4_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003625(.in0(tmp01_10_28), .in1(tmp01_11_28), .out(tmp02_5_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003626(.in0(tmp01_12_28), .in1(tmp01_13_28), .out(tmp02_6_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003627(.in0(tmp01_14_28), .in1(tmp01_15_28), .out(tmp02_7_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003628(.in0(tmp01_16_28), .in1(tmp01_17_28), .out(tmp02_8_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003629(.in0(tmp01_18_28), .in1(tmp01_19_28), .out(tmp02_9_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003630(.in0(tmp01_20_28), .in1(tmp01_21_28), .out(tmp02_10_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003631(.in0(tmp01_22_28), .in1(tmp01_23_28), .out(tmp02_11_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003632(.in0(tmp01_24_28), .in1(tmp01_25_28), .out(tmp02_12_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003633(.in0(tmp01_26_28), .in1(tmp01_27_28), .out(tmp02_13_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003634(.in0(tmp01_28_28), .in1(tmp01_29_28), .out(tmp02_14_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003635(.in0(tmp01_30_28), .in1(tmp01_31_28), .out(tmp02_15_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003636(.in0(tmp01_32_28), .in1(tmp01_33_28), .out(tmp02_16_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003637(.in0(tmp01_34_28), .in1(tmp01_35_28), .out(tmp02_17_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003638(.in0(tmp01_36_28), .in1(tmp01_37_28), .out(tmp02_18_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003639(.in0(tmp01_38_28), .in1(tmp01_39_28), .out(tmp02_19_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003640(.in0(tmp01_40_28), .in1(tmp01_41_28), .out(tmp02_20_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003641(.in0(tmp01_42_28), .in1(tmp01_43_28), .out(tmp02_21_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003642(.in0(tmp01_44_28), .in1(tmp01_45_28), .out(tmp02_22_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003643(.in0(tmp01_46_28), .in1(tmp01_47_28), .out(tmp02_23_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003644(.in0(tmp01_48_28), .in1(tmp01_49_28), .out(tmp02_24_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003645(.in0(tmp01_50_28), .in1(tmp01_51_28), .out(tmp02_25_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003646(.in0(tmp01_52_28), .in1(tmp01_53_28), .out(tmp02_26_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003647(.in0(tmp01_54_28), .in1(tmp01_55_28), .out(tmp02_27_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003648(.in0(tmp01_56_28), .in1(tmp01_57_28), .out(tmp02_28_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003649(.in0(tmp01_58_28), .in1(tmp01_59_28), .out(tmp02_29_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003650(.in0(tmp01_60_28), .in1(tmp01_61_28), .out(tmp02_30_28));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003651(.in0(tmp01_62_28), .in1(tmp01_63_28), .out(tmp02_31_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003652(.in0(tmp02_0_28), .in1(tmp02_1_28), .out(tmp03_0_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003653(.in0(tmp02_2_28), .in1(tmp02_3_28), .out(tmp03_1_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003654(.in0(tmp02_4_28), .in1(tmp02_5_28), .out(tmp03_2_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003655(.in0(tmp02_6_28), .in1(tmp02_7_28), .out(tmp03_3_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003656(.in0(tmp02_8_28), .in1(tmp02_9_28), .out(tmp03_4_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003657(.in0(tmp02_10_28), .in1(tmp02_11_28), .out(tmp03_5_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003658(.in0(tmp02_12_28), .in1(tmp02_13_28), .out(tmp03_6_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003659(.in0(tmp02_14_28), .in1(tmp02_15_28), .out(tmp03_7_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003660(.in0(tmp02_16_28), .in1(tmp02_17_28), .out(tmp03_8_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003661(.in0(tmp02_18_28), .in1(tmp02_19_28), .out(tmp03_9_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003662(.in0(tmp02_20_28), .in1(tmp02_21_28), .out(tmp03_10_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003663(.in0(tmp02_22_28), .in1(tmp02_23_28), .out(tmp03_11_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003664(.in0(tmp02_24_28), .in1(tmp02_25_28), .out(tmp03_12_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003665(.in0(tmp02_26_28), .in1(tmp02_27_28), .out(tmp03_13_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003666(.in0(tmp02_28_28), .in1(tmp02_29_28), .out(tmp03_14_28));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003667(.in0(tmp02_30_28), .in1(tmp02_31_28), .out(tmp03_15_28));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003668(.in0(tmp03_0_28), .in1(tmp03_1_28), .out(tmp04_0_28));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003669(.in0(tmp03_2_28), .in1(tmp03_3_28), .out(tmp04_1_28));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003670(.in0(tmp03_4_28), .in1(tmp03_5_28), .out(tmp04_2_28));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003671(.in0(tmp03_6_28), .in1(tmp03_7_28), .out(tmp04_3_28));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003672(.in0(tmp03_8_28), .in1(tmp03_9_28), .out(tmp04_4_28));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003673(.in0(tmp03_10_28), .in1(tmp03_11_28), .out(tmp04_5_28));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003674(.in0(tmp03_12_28), .in1(tmp03_13_28), .out(tmp04_6_28));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003675(.in0(tmp03_14_28), .in1(tmp03_15_28), .out(tmp04_7_28));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003676(.in0(tmp04_0_28), .in1(tmp04_1_28), .out(tmp05_0_28));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003677(.in0(tmp04_2_28), .in1(tmp04_3_28), .out(tmp05_1_28));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003678(.in0(tmp04_4_28), .in1(tmp04_5_28), .out(tmp05_2_28));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003679(.in0(tmp04_6_28), .in1(tmp04_7_28), .out(tmp05_3_28));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003680(.in0(tmp05_0_28), .in1(tmp05_1_28), .out(tmp06_0_28));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003681(.in0(tmp05_2_28), .in1(tmp05_3_28), .out(tmp06_1_28));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add003682(.in0(tmp06_0_28), .in1(tmp06_1_28), .out(tmp07_0_28));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003683(.in0(tmp00_0_29), .in1(tmp00_1_29), .out(tmp01_0_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003684(.in0(tmp00_2_29), .in1(tmp00_3_29), .out(tmp01_1_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003685(.in0(tmp00_4_29), .in1(tmp00_5_29), .out(tmp01_2_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003686(.in0(tmp00_6_29), .in1(tmp00_7_29), .out(tmp01_3_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003687(.in0(tmp00_8_29), .in1(tmp00_9_29), .out(tmp01_4_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003688(.in0(tmp00_10_29), .in1(tmp00_11_29), .out(tmp01_5_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003689(.in0(tmp00_12_29), .in1(tmp00_13_29), .out(tmp01_6_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003690(.in0(tmp00_14_29), .in1(tmp00_15_29), .out(tmp01_7_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003691(.in0(tmp00_16_29), .in1(tmp00_17_29), .out(tmp01_8_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003692(.in0(tmp00_18_29), .in1(tmp00_19_29), .out(tmp01_9_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003693(.in0(tmp00_20_29), .in1(tmp00_21_29), .out(tmp01_10_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003694(.in0(tmp00_22_29), .in1(tmp00_23_29), .out(tmp01_11_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003695(.in0(tmp00_24_29), .in1(tmp00_25_29), .out(tmp01_12_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003696(.in0(tmp00_26_29), .in1(tmp00_27_29), .out(tmp01_13_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003697(.in0(tmp00_28_29), .in1(tmp00_29_29), .out(tmp01_14_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003698(.in0(tmp00_30_29), .in1(tmp00_31_29), .out(tmp01_15_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003699(.in0(tmp00_32_29), .in1(tmp00_33_29), .out(tmp01_16_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003700(.in0(tmp00_34_29), .in1(tmp00_35_29), .out(tmp01_17_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003701(.in0(tmp00_36_29), .in1(tmp00_37_29), .out(tmp01_18_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003702(.in0(tmp00_38_29), .in1(tmp00_39_29), .out(tmp01_19_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003703(.in0(tmp00_40_29), .in1(tmp00_41_29), .out(tmp01_20_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003704(.in0(tmp00_42_29), .in1(tmp00_43_29), .out(tmp01_21_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003705(.in0(tmp00_44_29), .in1(tmp00_45_29), .out(tmp01_22_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003706(.in0(tmp00_46_29), .in1(tmp00_47_29), .out(tmp01_23_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003707(.in0(tmp00_48_29), .in1(tmp00_49_29), .out(tmp01_24_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003708(.in0(tmp00_50_29), .in1(tmp00_51_29), .out(tmp01_25_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003709(.in0(tmp00_52_29), .in1(tmp00_53_29), .out(tmp01_26_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003710(.in0(tmp00_54_29), .in1(tmp00_55_29), .out(tmp01_27_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003711(.in0(tmp00_56_29), .in1(tmp00_57_29), .out(tmp01_28_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003712(.in0(tmp00_58_29), .in1(tmp00_59_29), .out(tmp01_29_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003713(.in0(tmp00_60_29), .in1(tmp00_61_29), .out(tmp01_30_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003714(.in0(tmp00_62_29), .in1(tmp00_63_29), .out(tmp01_31_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003715(.in0(tmp00_64_29), .in1(tmp00_65_29), .out(tmp01_32_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003716(.in0(tmp00_66_29), .in1(tmp00_67_29), .out(tmp01_33_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003717(.in0(tmp00_68_29), .in1(tmp00_69_29), .out(tmp01_34_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003718(.in0(tmp00_70_29), .in1(tmp00_71_29), .out(tmp01_35_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003719(.in0(tmp00_72_29), .in1(tmp00_73_29), .out(tmp01_36_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003720(.in0(tmp00_74_29), .in1(tmp00_75_29), .out(tmp01_37_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003721(.in0(tmp00_76_29), .in1(tmp00_77_29), .out(tmp01_38_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003722(.in0(tmp00_78_29), .in1(tmp00_79_29), .out(tmp01_39_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003723(.in0(tmp00_80_29), .in1(tmp00_81_29), .out(tmp01_40_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003724(.in0(tmp00_82_29), .in1(tmp00_83_29), .out(tmp01_41_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003725(.in0(tmp00_84_29), .in1(tmp00_85_29), .out(tmp01_42_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003726(.in0(tmp00_86_29), .in1(tmp00_87_29), .out(tmp01_43_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003727(.in0(tmp00_88_29), .in1(tmp00_89_29), .out(tmp01_44_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003728(.in0(tmp00_90_29), .in1(tmp00_91_29), .out(tmp01_45_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003729(.in0(tmp00_92_29), .in1(tmp00_93_29), .out(tmp01_46_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003730(.in0(tmp00_94_29), .in1(tmp00_95_29), .out(tmp01_47_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003731(.in0(tmp00_96_29), .in1(tmp00_97_29), .out(tmp01_48_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003732(.in0(tmp00_98_29), .in1(tmp00_99_29), .out(tmp01_49_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003733(.in0(tmp00_100_29), .in1(tmp00_101_29), .out(tmp01_50_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003734(.in0(tmp00_102_29), .in1(tmp00_103_29), .out(tmp01_51_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003735(.in0(tmp00_104_29), .in1(tmp00_105_29), .out(tmp01_52_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003736(.in0(tmp00_106_29), .in1(tmp00_107_29), .out(tmp01_53_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003737(.in0(tmp00_108_29), .in1(tmp00_109_29), .out(tmp01_54_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003738(.in0(tmp00_110_29), .in1(tmp00_111_29), .out(tmp01_55_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003739(.in0(tmp00_112_29), .in1(tmp00_113_29), .out(tmp01_56_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003740(.in0(tmp00_114_29), .in1(tmp00_115_29), .out(tmp01_57_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003741(.in0(tmp00_116_29), .in1(tmp00_117_29), .out(tmp01_58_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003742(.in0(tmp00_118_29), .in1(tmp00_119_29), .out(tmp01_59_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003743(.in0(tmp00_120_29), .in1(tmp00_121_29), .out(tmp01_60_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003744(.in0(tmp00_122_29), .in1(tmp00_123_29), .out(tmp01_61_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003745(.in0(tmp00_124_29), .in1(tmp00_125_29), .out(tmp01_62_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003746(.in0(tmp00_126_29), .in1(tmp00_127_29), .out(tmp01_63_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003747(.in0(tmp01_0_29), .in1(tmp01_1_29), .out(tmp02_0_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003748(.in0(tmp01_2_29), .in1(tmp01_3_29), .out(tmp02_1_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003749(.in0(tmp01_4_29), .in1(tmp01_5_29), .out(tmp02_2_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003750(.in0(tmp01_6_29), .in1(tmp01_7_29), .out(tmp02_3_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003751(.in0(tmp01_8_29), .in1(tmp01_9_29), .out(tmp02_4_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003752(.in0(tmp01_10_29), .in1(tmp01_11_29), .out(tmp02_5_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003753(.in0(tmp01_12_29), .in1(tmp01_13_29), .out(tmp02_6_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003754(.in0(tmp01_14_29), .in1(tmp01_15_29), .out(tmp02_7_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003755(.in0(tmp01_16_29), .in1(tmp01_17_29), .out(tmp02_8_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003756(.in0(tmp01_18_29), .in1(tmp01_19_29), .out(tmp02_9_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003757(.in0(tmp01_20_29), .in1(tmp01_21_29), .out(tmp02_10_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003758(.in0(tmp01_22_29), .in1(tmp01_23_29), .out(tmp02_11_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003759(.in0(tmp01_24_29), .in1(tmp01_25_29), .out(tmp02_12_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003760(.in0(tmp01_26_29), .in1(tmp01_27_29), .out(tmp02_13_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003761(.in0(tmp01_28_29), .in1(tmp01_29_29), .out(tmp02_14_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003762(.in0(tmp01_30_29), .in1(tmp01_31_29), .out(tmp02_15_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003763(.in0(tmp01_32_29), .in1(tmp01_33_29), .out(tmp02_16_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003764(.in0(tmp01_34_29), .in1(tmp01_35_29), .out(tmp02_17_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003765(.in0(tmp01_36_29), .in1(tmp01_37_29), .out(tmp02_18_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003766(.in0(tmp01_38_29), .in1(tmp01_39_29), .out(tmp02_19_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003767(.in0(tmp01_40_29), .in1(tmp01_41_29), .out(tmp02_20_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003768(.in0(tmp01_42_29), .in1(tmp01_43_29), .out(tmp02_21_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003769(.in0(tmp01_44_29), .in1(tmp01_45_29), .out(tmp02_22_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003770(.in0(tmp01_46_29), .in1(tmp01_47_29), .out(tmp02_23_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003771(.in0(tmp01_48_29), .in1(tmp01_49_29), .out(tmp02_24_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003772(.in0(tmp01_50_29), .in1(tmp01_51_29), .out(tmp02_25_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003773(.in0(tmp01_52_29), .in1(tmp01_53_29), .out(tmp02_26_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003774(.in0(tmp01_54_29), .in1(tmp01_55_29), .out(tmp02_27_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003775(.in0(tmp01_56_29), .in1(tmp01_57_29), .out(tmp02_28_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003776(.in0(tmp01_58_29), .in1(tmp01_59_29), .out(tmp02_29_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003777(.in0(tmp01_60_29), .in1(tmp01_61_29), .out(tmp02_30_29));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003778(.in0(tmp01_62_29), .in1(tmp01_63_29), .out(tmp02_31_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003779(.in0(tmp02_0_29), .in1(tmp02_1_29), .out(tmp03_0_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003780(.in0(tmp02_2_29), .in1(tmp02_3_29), .out(tmp03_1_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003781(.in0(tmp02_4_29), .in1(tmp02_5_29), .out(tmp03_2_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003782(.in0(tmp02_6_29), .in1(tmp02_7_29), .out(tmp03_3_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003783(.in0(tmp02_8_29), .in1(tmp02_9_29), .out(tmp03_4_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003784(.in0(tmp02_10_29), .in1(tmp02_11_29), .out(tmp03_5_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003785(.in0(tmp02_12_29), .in1(tmp02_13_29), .out(tmp03_6_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003786(.in0(tmp02_14_29), .in1(tmp02_15_29), .out(tmp03_7_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003787(.in0(tmp02_16_29), .in1(tmp02_17_29), .out(tmp03_8_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003788(.in0(tmp02_18_29), .in1(tmp02_19_29), .out(tmp03_9_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003789(.in0(tmp02_20_29), .in1(tmp02_21_29), .out(tmp03_10_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003790(.in0(tmp02_22_29), .in1(tmp02_23_29), .out(tmp03_11_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003791(.in0(tmp02_24_29), .in1(tmp02_25_29), .out(tmp03_12_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003792(.in0(tmp02_26_29), .in1(tmp02_27_29), .out(tmp03_13_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003793(.in0(tmp02_28_29), .in1(tmp02_29_29), .out(tmp03_14_29));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003794(.in0(tmp02_30_29), .in1(tmp02_31_29), .out(tmp03_15_29));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003795(.in0(tmp03_0_29), .in1(tmp03_1_29), .out(tmp04_0_29));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003796(.in0(tmp03_2_29), .in1(tmp03_3_29), .out(tmp04_1_29));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003797(.in0(tmp03_4_29), .in1(tmp03_5_29), .out(tmp04_2_29));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003798(.in0(tmp03_6_29), .in1(tmp03_7_29), .out(tmp04_3_29));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003799(.in0(tmp03_8_29), .in1(tmp03_9_29), .out(tmp04_4_29));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003800(.in0(tmp03_10_29), .in1(tmp03_11_29), .out(tmp04_5_29));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003801(.in0(tmp03_12_29), .in1(tmp03_13_29), .out(tmp04_6_29));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003802(.in0(tmp03_14_29), .in1(tmp03_15_29), .out(tmp04_7_29));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003803(.in0(tmp04_0_29), .in1(tmp04_1_29), .out(tmp05_0_29));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003804(.in0(tmp04_2_29), .in1(tmp04_3_29), .out(tmp05_1_29));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003805(.in0(tmp04_4_29), .in1(tmp04_5_29), .out(tmp05_2_29));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003806(.in0(tmp04_6_29), .in1(tmp04_7_29), .out(tmp05_3_29));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003807(.in0(tmp05_0_29), .in1(tmp05_1_29), .out(tmp06_0_29));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003808(.in0(tmp05_2_29), .in1(tmp05_3_29), .out(tmp06_1_29));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add003809(.in0(tmp06_0_29), .in1(tmp06_1_29), .out(tmp07_0_29));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003810(.in0(tmp00_0_30), .in1(tmp00_1_30), .out(tmp01_0_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003811(.in0(tmp00_2_30), .in1(tmp00_3_30), .out(tmp01_1_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003812(.in0(tmp00_4_30), .in1(tmp00_5_30), .out(tmp01_2_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003813(.in0(tmp00_6_30), .in1(tmp00_7_30), .out(tmp01_3_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003814(.in0(tmp00_8_30), .in1(tmp00_9_30), .out(tmp01_4_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003815(.in0(tmp00_10_30), .in1(tmp00_11_30), .out(tmp01_5_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003816(.in0(tmp00_12_30), .in1(tmp00_13_30), .out(tmp01_6_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003817(.in0(tmp00_14_30), .in1(tmp00_15_30), .out(tmp01_7_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003818(.in0(tmp00_16_30), .in1(tmp00_17_30), .out(tmp01_8_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003819(.in0(tmp00_18_30), .in1(tmp00_19_30), .out(tmp01_9_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003820(.in0(tmp00_20_30), .in1(tmp00_21_30), .out(tmp01_10_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003821(.in0(tmp00_22_30), .in1(tmp00_23_30), .out(tmp01_11_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003822(.in0(tmp00_24_30), .in1(tmp00_25_30), .out(tmp01_12_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003823(.in0(tmp00_26_30), .in1(tmp00_27_30), .out(tmp01_13_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003824(.in0(tmp00_28_30), .in1(tmp00_29_30), .out(tmp01_14_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003825(.in0(tmp00_30_30), .in1(tmp00_31_30), .out(tmp01_15_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003826(.in0(tmp00_32_30), .in1(tmp00_33_30), .out(tmp01_16_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003827(.in0(tmp00_34_30), .in1(tmp00_35_30), .out(tmp01_17_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003828(.in0(tmp00_36_30), .in1(tmp00_37_30), .out(tmp01_18_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003829(.in0(tmp00_38_30), .in1(tmp00_39_30), .out(tmp01_19_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003830(.in0(tmp00_40_30), .in1(tmp00_41_30), .out(tmp01_20_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003831(.in0(tmp00_42_30), .in1(tmp00_43_30), .out(tmp01_21_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003832(.in0(tmp00_44_30), .in1(tmp00_45_30), .out(tmp01_22_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003833(.in0(tmp00_46_30), .in1(tmp00_47_30), .out(tmp01_23_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003834(.in0(tmp00_48_30), .in1(tmp00_49_30), .out(tmp01_24_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003835(.in0(tmp00_50_30), .in1(tmp00_51_30), .out(tmp01_25_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003836(.in0(tmp00_52_30), .in1(tmp00_53_30), .out(tmp01_26_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003837(.in0(tmp00_54_30), .in1(tmp00_55_30), .out(tmp01_27_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003838(.in0(tmp00_56_30), .in1(tmp00_57_30), .out(tmp01_28_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003839(.in0(tmp00_58_30), .in1(tmp00_59_30), .out(tmp01_29_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003840(.in0(tmp00_60_30), .in1(tmp00_61_30), .out(tmp01_30_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003841(.in0(tmp00_62_30), .in1(tmp00_63_30), .out(tmp01_31_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003842(.in0(tmp00_64_30), .in1(tmp00_65_30), .out(tmp01_32_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003843(.in0(tmp00_66_30), .in1(tmp00_67_30), .out(tmp01_33_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003844(.in0(tmp00_68_30), .in1(tmp00_69_30), .out(tmp01_34_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003845(.in0(tmp00_70_30), .in1(tmp00_71_30), .out(tmp01_35_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003846(.in0(tmp00_72_30), .in1(tmp00_73_30), .out(tmp01_36_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003847(.in0(tmp00_74_30), .in1(tmp00_75_30), .out(tmp01_37_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003848(.in0(tmp00_76_30), .in1(tmp00_77_30), .out(tmp01_38_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003849(.in0(tmp00_78_30), .in1(tmp00_79_30), .out(tmp01_39_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003850(.in0(tmp00_80_30), .in1(tmp00_81_30), .out(tmp01_40_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003851(.in0(tmp00_82_30), .in1(tmp00_83_30), .out(tmp01_41_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003852(.in0(tmp00_84_30), .in1(tmp00_85_30), .out(tmp01_42_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003853(.in0(tmp00_86_30), .in1(tmp00_87_30), .out(tmp01_43_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003854(.in0(tmp00_88_30), .in1(tmp00_89_30), .out(tmp01_44_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003855(.in0(tmp00_90_30), .in1(tmp00_91_30), .out(tmp01_45_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003856(.in0(tmp00_92_30), .in1(tmp00_93_30), .out(tmp01_46_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003857(.in0(tmp00_94_30), .in1(tmp00_95_30), .out(tmp01_47_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003858(.in0(tmp00_96_30), .in1(tmp00_97_30), .out(tmp01_48_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003859(.in0(tmp00_98_30), .in1(tmp00_99_30), .out(tmp01_49_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003860(.in0(tmp00_100_30), .in1(tmp00_101_30), .out(tmp01_50_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003861(.in0(tmp00_102_30), .in1(tmp00_103_30), .out(tmp01_51_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003862(.in0(tmp00_104_30), .in1(tmp00_105_30), .out(tmp01_52_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003863(.in0(tmp00_106_30), .in1(tmp00_107_30), .out(tmp01_53_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003864(.in0(tmp00_108_30), .in1(tmp00_109_30), .out(tmp01_54_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003865(.in0(tmp00_110_30), .in1(tmp00_111_30), .out(tmp01_55_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003866(.in0(tmp00_112_30), .in1(tmp00_113_30), .out(tmp01_56_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003867(.in0(tmp00_114_30), .in1(tmp00_115_30), .out(tmp01_57_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003868(.in0(tmp00_116_30), .in1(tmp00_117_30), .out(tmp01_58_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003869(.in0(tmp00_118_30), .in1(tmp00_119_30), .out(tmp01_59_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003870(.in0(tmp00_120_30), .in1(tmp00_121_30), .out(tmp01_60_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003871(.in0(tmp00_122_30), .in1(tmp00_123_30), .out(tmp01_61_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003872(.in0(tmp00_124_30), .in1(tmp00_125_30), .out(tmp01_62_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003873(.in0(tmp00_126_30), .in1(tmp00_127_30), .out(tmp01_63_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003874(.in0(tmp01_0_30), .in1(tmp01_1_30), .out(tmp02_0_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003875(.in0(tmp01_2_30), .in1(tmp01_3_30), .out(tmp02_1_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003876(.in0(tmp01_4_30), .in1(tmp01_5_30), .out(tmp02_2_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003877(.in0(tmp01_6_30), .in1(tmp01_7_30), .out(tmp02_3_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003878(.in0(tmp01_8_30), .in1(tmp01_9_30), .out(tmp02_4_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003879(.in0(tmp01_10_30), .in1(tmp01_11_30), .out(tmp02_5_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003880(.in0(tmp01_12_30), .in1(tmp01_13_30), .out(tmp02_6_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003881(.in0(tmp01_14_30), .in1(tmp01_15_30), .out(tmp02_7_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003882(.in0(tmp01_16_30), .in1(tmp01_17_30), .out(tmp02_8_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003883(.in0(tmp01_18_30), .in1(tmp01_19_30), .out(tmp02_9_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003884(.in0(tmp01_20_30), .in1(tmp01_21_30), .out(tmp02_10_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003885(.in0(tmp01_22_30), .in1(tmp01_23_30), .out(tmp02_11_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003886(.in0(tmp01_24_30), .in1(tmp01_25_30), .out(tmp02_12_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003887(.in0(tmp01_26_30), .in1(tmp01_27_30), .out(tmp02_13_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003888(.in0(tmp01_28_30), .in1(tmp01_29_30), .out(tmp02_14_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003889(.in0(tmp01_30_30), .in1(tmp01_31_30), .out(tmp02_15_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003890(.in0(tmp01_32_30), .in1(tmp01_33_30), .out(tmp02_16_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003891(.in0(tmp01_34_30), .in1(tmp01_35_30), .out(tmp02_17_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003892(.in0(tmp01_36_30), .in1(tmp01_37_30), .out(tmp02_18_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003893(.in0(tmp01_38_30), .in1(tmp01_39_30), .out(tmp02_19_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003894(.in0(tmp01_40_30), .in1(tmp01_41_30), .out(tmp02_20_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003895(.in0(tmp01_42_30), .in1(tmp01_43_30), .out(tmp02_21_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003896(.in0(tmp01_44_30), .in1(tmp01_45_30), .out(tmp02_22_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003897(.in0(tmp01_46_30), .in1(tmp01_47_30), .out(tmp02_23_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003898(.in0(tmp01_48_30), .in1(tmp01_49_30), .out(tmp02_24_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003899(.in0(tmp01_50_30), .in1(tmp01_51_30), .out(tmp02_25_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003900(.in0(tmp01_52_30), .in1(tmp01_53_30), .out(tmp02_26_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003901(.in0(tmp01_54_30), .in1(tmp01_55_30), .out(tmp02_27_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003902(.in0(tmp01_56_30), .in1(tmp01_57_30), .out(tmp02_28_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003903(.in0(tmp01_58_30), .in1(tmp01_59_30), .out(tmp02_29_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003904(.in0(tmp01_60_30), .in1(tmp01_61_30), .out(tmp02_30_30));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add003905(.in0(tmp01_62_30), .in1(tmp01_63_30), .out(tmp02_31_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003906(.in0(tmp02_0_30), .in1(tmp02_1_30), .out(tmp03_0_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003907(.in0(tmp02_2_30), .in1(tmp02_3_30), .out(tmp03_1_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003908(.in0(tmp02_4_30), .in1(tmp02_5_30), .out(tmp03_2_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003909(.in0(tmp02_6_30), .in1(tmp02_7_30), .out(tmp03_3_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003910(.in0(tmp02_8_30), .in1(tmp02_9_30), .out(tmp03_4_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003911(.in0(tmp02_10_30), .in1(tmp02_11_30), .out(tmp03_5_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003912(.in0(tmp02_12_30), .in1(tmp02_13_30), .out(tmp03_6_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003913(.in0(tmp02_14_30), .in1(tmp02_15_30), .out(tmp03_7_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003914(.in0(tmp02_16_30), .in1(tmp02_17_30), .out(tmp03_8_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003915(.in0(tmp02_18_30), .in1(tmp02_19_30), .out(tmp03_9_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003916(.in0(tmp02_20_30), .in1(tmp02_21_30), .out(tmp03_10_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003917(.in0(tmp02_22_30), .in1(tmp02_23_30), .out(tmp03_11_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003918(.in0(tmp02_24_30), .in1(tmp02_25_30), .out(tmp03_12_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003919(.in0(tmp02_26_30), .in1(tmp02_27_30), .out(tmp03_13_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003920(.in0(tmp02_28_30), .in1(tmp02_29_30), .out(tmp03_14_30));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add003921(.in0(tmp02_30_30), .in1(tmp02_31_30), .out(tmp03_15_30));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003922(.in0(tmp03_0_30), .in1(tmp03_1_30), .out(tmp04_0_30));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003923(.in0(tmp03_2_30), .in1(tmp03_3_30), .out(tmp04_1_30));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003924(.in0(tmp03_4_30), .in1(tmp03_5_30), .out(tmp04_2_30));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003925(.in0(tmp03_6_30), .in1(tmp03_7_30), .out(tmp04_3_30));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003926(.in0(tmp03_8_30), .in1(tmp03_9_30), .out(tmp04_4_30));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003927(.in0(tmp03_10_30), .in1(tmp03_11_30), .out(tmp04_5_30));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003928(.in0(tmp03_12_30), .in1(tmp03_13_30), .out(tmp04_6_30));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add003929(.in0(tmp03_14_30), .in1(tmp03_15_30), .out(tmp04_7_30));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003930(.in0(tmp04_0_30), .in1(tmp04_1_30), .out(tmp05_0_30));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003931(.in0(tmp04_2_30), .in1(tmp04_3_30), .out(tmp05_1_30));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003932(.in0(tmp04_4_30), .in1(tmp04_5_30), .out(tmp05_2_30));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add003933(.in0(tmp04_6_30), .in1(tmp04_7_30), .out(tmp05_3_30));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003934(.in0(tmp05_0_30), .in1(tmp05_1_30), .out(tmp06_0_30));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add003935(.in0(tmp05_2_30), .in1(tmp05_3_30), .out(tmp06_1_30));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add003936(.in0(tmp06_0_30), .in1(tmp06_1_30), .out(tmp07_0_30));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003937(.in0(tmp00_0_31), .in1(tmp00_1_31), .out(tmp01_0_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003938(.in0(tmp00_2_31), .in1(tmp00_3_31), .out(tmp01_1_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003939(.in0(tmp00_4_31), .in1(tmp00_5_31), .out(tmp01_2_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003940(.in0(tmp00_6_31), .in1(tmp00_7_31), .out(tmp01_3_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003941(.in0(tmp00_8_31), .in1(tmp00_9_31), .out(tmp01_4_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003942(.in0(tmp00_10_31), .in1(tmp00_11_31), .out(tmp01_5_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003943(.in0(tmp00_12_31), .in1(tmp00_13_31), .out(tmp01_6_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003944(.in0(tmp00_14_31), .in1(tmp00_15_31), .out(tmp01_7_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003945(.in0(tmp00_16_31), .in1(tmp00_17_31), .out(tmp01_8_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003946(.in0(tmp00_18_31), .in1(tmp00_19_31), .out(tmp01_9_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003947(.in0(tmp00_20_31), .in1(tmp00_21_31), .out(tmp01_10_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003948(.in0(tmp00_22_31), .in1(tmp00_23_31), .out(tmp01_11_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003949(.in0(tmp00_24_31), .in1(tmp00_25_31), .out(tmp01_12_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003950(.in0(tmp00_26_31), .in1(tmp00_27_31), .out(tmp01_13_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003951(.in0(tmp00_28_31), .in1(tmp00_29_31), .out(tmp01_14_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003952(.in0(tmp00_30_31), .in1(tmp00_31_31), .out(tmp01_15_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003953(.in0(tmp00_32_31), .in1(tmp00_33_31), .out(tmp01_16_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003954(.in0(tmp00_34_31), .in1(tmp00_35_31), .out(tmp01_17_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003955(.in0(tmp00_36_31), .in1(tmp00_37_31), .out(tmp01_18_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003956(.in0(tmp00_38_31), .in1(tmp00_39_31), .out(tmp01_19_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003957(.in0(tmp00_40_31), .in1(tmp00_41_31), .out(tmp01_20_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003958(.in0(tmp00_42_31), .in1(tmp00_43_31), .out(tmp01_21_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003959(.in0(tmp00_44_31), .in1(tmp00_45_31), .out(tmp01_22_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003960(.in0(tmp00_46_31), .in1(tmp00_47_31), .out(tmp01_23_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003961(.in0(tmp00_48_31), .in1(tmp00_49_31), .out(tmp01_24_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003962(.in0(tmp00_50_31), .in1(tmp00_51_31), .out(tmp01_25_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003963(.in0(tmp00_52_31), .in1(tmp00_53_31), .out(tmp01_26_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003964(.in0(tmp00_54_31), .in1(tmp00_55_31), .out(tmp01_27_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003965(.in0(tmp00_56_31), .in1(tmp00_57_31), .out(tmp01_28_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003966(.in0(tmp00_58_31), .in1(tmp00_59_31), .out(tmp01_29_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003967(.in0(tmp00_60_31), .in1(tmp00_61_31), .out(tmp01_30_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003968(.in0(tmp00_62_31), .in1(tmp00_63_31), .out(tmp01_31_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003969(.in0(tmp00_64_31), .in1(tmp00_65_31), .out(tmp01_32_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003970(.in0(tmp00_66_31), .in1(tmp00_67_31), .out(tmp01_33_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003971(.in0(tmp00_68_31), .in1(tmp00_69_31), .out(tmp01_34_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003972(.in0(tmp00_70_31), .in1(tmp00_71_31), .out(tmp01_35_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003973(.in0(tmp00_72_31), .in1(tmp00_73_31), .out(tmp01_36_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003974(.in0(tmp00_74_31), .in1(tmp00_75_31), .out(tmp01_37_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003975(.in0(tmp00_76_31), .in1(tmp00_77_31), .out(tmp01_38_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003976(.in0(tmp00_78_31), .in1(tmp00_79_31), .out(tmp01_39_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003977(.in0(tmp00_80_31), .in1(tmp00_81_31), .out(tmp01_40_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003978(.in0(tmp00_82_31), .in1(tmp00_83_31), .out(tmp01_41_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003979(.in0(tmp00_84_31), .in1(tmp00_85_31), .out(tmp01_42_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003980(.in0(tmp00_86_31), .in1(tmp00_87_31), .out(tmp01_43_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003981(.in0(tmp00_88_31), .in1(tmp00_89_31), .out(tmp01_44_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003982(.in0(tmp00_90_31), .in1(tmp00_91_31), .out(tmp01_45_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003983(.in0(tmp00_92_31), .in1(tmp00_93_31), .out(tmp01_46_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003984(.in0(tmp00_94_31), .in1(tmp00_95_31), .out(tmp01_47_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003985(.in0(tmp00_96_31), .in1(tmp00_97_31), .out(tmp01_48_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003986(.in0(tmp00_98_31), .in1(tmp00_99_31), .out(tmp01_49_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003987(.in0(tmp00_100_31), .in1(tmp00_101_31), .out(tmp01_50_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003988(.in0(tmp00_102_31), .in1(tmp00_103_31), .out(tmp01_51_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003989(.in0(tmp00_104_31), .in1(tmp00_105_31), .out(tmp01_52_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003990(.in0(tmp00_106_31), .in1(tmp00_107_31), .out(tmp01_53_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003991(.in0(tmp00_108_31), .in1(tmp00_109_31), .out(tmp01_54_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003992(.in0(tmp00_110_31), .in1(tmp00_111_31), .out(tmp01_55_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003993(.in0(tmp00_112_31), .in1(tmp00_113_31), .out(tmp01_56_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003994(.in0(tmp00_114_31), .in1(tmp00_115_31), .out(tmp01_57_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003995(.in0(tmp00_116_31), .in1(tmp00_117_31), .out(tmp01_58_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003996(.in0(tmp00_118_31), .in1(tmp00_119_31), .out(tmp01_59_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003997(.in0(tmp00_120_31), .in1(tmp00_121_31), .out(tmp01_60_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003998(.in0(tmp00_122_31), .in1(tmp00_123_31), .out(tmp01_61_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add003999(.in0(tmp00_124_31), .in1(tmp00_125_31), .out(tmp01_62_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004000(.in0(tmp00_126_31), .in1(tmp00_127_31), .out(tmp01_63_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004001(.in0(tmp01_0_31), .in1(tmp01_1_31), .out(tmp02_0_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004002(.in0(tmp01_2_31), .in1(tmp01_3_31), .out(tmp02_1_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004003(.in0(tmp01_4_31), .in1(tmp01_5_31), .out(tmp02_2_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004004(.in0(tmp01_6_31), .in1(tmp01_7_31), .out(tmp02_3_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004005(.in0(tmp01_8_31), .in1(tmp01_9_31), .out(tmp02_4_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004006(.in0(tmp01_10_31), .in1(tmp01_11_31), .out(tmp02_5_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004007(.in0(tmp01_12_31), .in1(tmp01_13_31), .out(tmp02_6_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004008(.in0(tmp01_14_31), .in1(tmp01_15_31), .out(tmp02_7_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004009(.in0(tmp01_16_31), .in1(tmp01_17_31), .out(tmp02_8_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004010(.in0(tmp01_18_31), .in1(tmp01_19_31), .out(tmp02_9_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004011(.in0(tmp01_20_31), .in1(tmp01_21_31), .out(tmp02_10_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004012(.in0(tmp01_22_31), .in1(tmp01_23_31), .out(tmp02_11_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004013(.in0(tmp01_24_31), .in1(tmp01_25_31), .out(tmp02_12_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004014(.in0(tmp01_26_31), .in1(tmp01_27_31), .out(tmp02_13_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004015(.in0(tmp01_28_31), .in1(tmp01_29_31), .out(tmp02_14_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004016(.in0(tmp01_30_31), .in1(tmp01_31_31), .out(tmp02_15_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004017(.in0(tmp01_32_31), .in1(tmp01_33_31), .out(tmp02_16_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004018(.in0(tmp01_34_31), .in1(tmp01_35_31), .out(tmp02_17_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004019(.in0(tmp01_36_31), .in1(tmp01_37_31), .out(tmp02_18_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004020(.in0(tmp01_38_31), .in1(tmp01_39_31), .out(tmp02_19_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004021(.in0(tmp01_40_31), .in1(tmp01_41_31), .out(tmp02_20_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004022(.in0(tmp01_42_31), .in1(tmp01_43_31), .out(tmp02_21_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004023(.in0(tmp01_44_31), .in1(tmp01_45_31), .out(tmp02_22_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004024(.in0(tmp01_46_31), .in1(tmp01_47_31), .out(tmp02_23_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004025(.in0(tmp01_48_31), .in1(tmp01_49_31), .out(tmp02_24_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004026(.in0(tmp01_50_31), .in1(tmp01_51_31), .out(tmp02_25_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004027(.in0(tmp01_52_31), .in1(tmp01_53_31), .out(tmp02_26_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004028(.in0(tmp01_54_31), .in1(tmp01_55_31), .out(tmp02_27_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004029(.in0(tmp01_56_31), .in1(tmp01_57_31), .out(tmp02_28_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004030(.in0(tmp01_58_31), .in1(tmp01_59_31), .out(tmp02_29_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004031(.in0(tmp01_60_31), .in1(tmp01_61_31), .out(tmp02_30_31));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004032(.in0(tmp01_62_31), .in1(tmp01_63_31), .out(tmp02_31_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004033(.in0(tmp02_0_31), .in1(tmp02_1_31), .out(tmp03_0_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004034(.in0(tmp02_2_31), .in1(tmp02_3_31), .out(tmp03_1_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004035(.in0(tmp02_4_31), .in1(tmp02_5_31), .out(tmp03_2_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004036(.in0(tmp02_6_31), .in1(tmp02_7_31), .out(tmp03_3_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004037(.in0(tmp02_8_31), .in1(tmp02_9_31), .out(tmp03_4_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004038(.in0(tmp02_10_31), .in1(tmp02_11_31), .out(tmp03_5_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004039(.in0(tmp02_12_31), .in1(tmp02_13_31), .out(tmp03_6_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004040(.in0(tmp02_14_31), .in1(tmp02_15_31), .out(tmp03_7_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004041(.in0(tmp02_16_31), .in1(tmp02_17_31), .out(tmp03_8_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004042(.in0(tmp02_18_31), .in1(tmp02_19_31), .out(tmp03_9_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004043(.in0(tmp02_20_31), .in1(tmp02_21_31), .out(tmp03_10_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004044(.in0(tmp02_22_31), .in1(tmp02_23_31), .out(tmp03_11_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004045(.in0(tmp02_24_31), .in1(tmp02_25_31), .out(tmp03_12_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004046(.in0(tmp02_26_31), .in1(tmp02_27_31), .out(tmp03_13_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004047(.in0(tmp02_28_31), .in1(tmp02_29_31), .out(tmp03_14_31));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004048(.in0(tmp02_30_31), .in1(tmp02_31_31), .out(tmp03_15_31));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004049(.in0(tmp03_0_31), .in1(tmp03_1_31), .out(tmp04_0_31));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004050(.in0(tmp03_2_31), .in1(tmp03_3_31), .out(tmp04_1_31));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004051(.in0(tmp03_4_31), .in1(tmp03_5_31), .out(tmp04_2_31));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004052(.in0(tmp03_6_31), .in1(tmp03_7_31), .out(tmp04_3_31));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004053(.in0(tmp03_8_31), .in1(tmp03_9_31), .out(tmp04_4_31));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004054(.in0(tmp03_10_31), .in1(tmp03_11_31), .out(tmp04_5_31));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004055(.in0(tmp03_12_31), .in1(tmp03_13_31), .out(tmp04_6_31));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004056(.in0(tmp03_14_31), .in1(tmp03_15_31), .out(tmp04_7_31));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004057(.in0(tmp04_0_31), .in1(tmp04_1_31), .out(tmp05_0_31));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004058(.in0(tmp04_2_31), .in1(tmp04_3_31), .out(tmp05_1_31));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004059(.in0(tmp04_4_31), .in1(tmp04_5_31), .out(tmp05_2_31));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004060(.in0(tmp04_6_31), .in1(tmp04_7_31), .out(tmp05_3_31));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004061(.in0(tmp05_0_31), .in1(tmp05_1_31), .out(tmp06_0_31));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004062(.in0(tmp05_2_31), .in1(tmp05_3_31), .out(tmp06_1_31));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add004063(.in0(tmp06_0_31), .in1(tmp06_1_31), .out(tmp07_0_31));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004064(.in0(tmp00_0_32), .in1(tmp00_1_32), .out(tmp01_0_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004065(.in0(tmp00_2_32), .in1(tmp00_3_32), .out(tmp01_1_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004066(.in0(tmp00_4_32), .in1(tmp00_5_32), .out(tmp01_2_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004067(.in0(tmp00_6_32), .in1(tmp00_7_32), .out(tmp01_3_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004068(.in0(tmp00_8_32), .in1(tmp00_9_32), .out(tmp01_4_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004069(.in0(tmp00_10_32), .in1(tmp00_11_32), .out(tmp01_5_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004070(.in0(tmp00_12_32), .in1(tmp00_13_32), .out(tmp01_6_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004071(.in0(tmp00_14_32), .in1(tmp00_15_32), .out(tmp01_7_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004072(.in0(tmp00_16_32), .in1(tmp00_17_32), .out(tmp01_8_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004073(.in0(tmp00_18_32), .in1(tmp00_19_32), .out(tmp01_9_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004074(.in0(tmp00_20_32), .in1(tmp00_21_32), .out(tmp01_10_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004075(.in0(tmp00_22_32), .in1(tmp00_23_32), .out(tmp01_11_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004076(.in0(tmp00_24_32), .in1(tmp00_25_32), .out(tmp01_12_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004077(.in0(tmp00_26_32), .in1(tmp00_27_32), .out(tmp01_13_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004078(.in0(tmp00_28_32), .in1(tmp00_29_32), .out(tmp01_14_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004079(.in0(tmp00_30_32), .in1(tmp00_31_32), .out(tmp01_15_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004080(.in0(tmp00_32_32), .in1(tmp00_33_32), .out(tmp01_16_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004081(.in0(tmp00_34_32), .in1(tmp00_35_32), .out(tmp01_17_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004082(.in0(tmp00_36_32), .in1(tmp00_37_32), .out(tmp01_18_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004083(.in0(tmp00_38_32), .in1(tmp00_39_32), .out(tmp01_19_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004084(.in0(tmp00_40_32), .in1(tmp00_41_32), .out(tmp01_20_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004085(.in0(tmp00_42_32), .in1(tmp00_43_32), .out(tmp01_21_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004086(.in0(tmp00_44_32), .in1(tmp00_45_32), .out(tmp01_22_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004087(.in0(tmp00_46_32), .in1(tmp00_47_32), .out(tmp01_23_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004088(.in0(tmp00_48_32), .in1(tmp00_49_32), .out(tmp01_24_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004089(.in0(tmp00_50_32), .in1(tmp00_51_32), .out(tmp01_25_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004090(.in0(tmp00_52_32), .in1(tmp00_53_32), .out(tmp01_26_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004091(.in0(tmp00_54_32), .in1(tmp00_55_32), .out(tmp01_27_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004092(.in0(tmp00_56_32), .in1(tmp00_57_32), .out(tmp01_28_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004093(.in0(tmp00_58_32), .in1(tmp00_59_32), .out(tmp01_29_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004094(.in0(tmp00_60_32), .in1(tmp00_61_32), .out(tmp01_30_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004095(.in0(tmp00_62_32), .in1(tmp00_63_32), .out(tmp01_31_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004096(.in0(tmp00_64_32), .in1(tmp00_65_32), .out(tmp01_32_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004097(.in0(tmp00_66_32), .in1(tmp00_67_32), .out(tmp01_33_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004098(.in0(tmp00_68_32), .in1(tmp00_69_32), .out(tmp01_34_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004099(.in0(tmp00_70_32), .in1(tmp00_71_32), .out(tmp01_35_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004100(.in0(tmp00_72_32), .in1(tmp00_73_32), .out(tmp01_36_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004101(.in0(tmp00_74_32), .in1(tmp00_75_32), .out(tmp01_37_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004102(.in0(tmp00_76_32), .in1(tmp00_77_32), .out(tmp01_38_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004103(.in0(tmp00_78_32), .in1(tmp00_79_32), .out(tmp01_39_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004104(.in0(tmp00_80_32), .in1(tmp00_81_32), .out(tmp01_40_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004105(.in0(tmp00_82_32), .in1(tmp00_83_32), .out(tmp01_41_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004106(.in0(tmp00_84_32), .in1(tmp00_85_32), .out(tmp01_42_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004107(.in0(tmp00_86_32), .in1(tmp00_87_32), .out(tmp01_43_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004108(.in0(tmp00_88_32), .in1(tmp00_89_32), .out(tmp01_44_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004109(.in0(tmp00_90_32), .in1(tmp00_91_32), .out(tmp01_45_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004110(.in0(tmp00_92_32), .in1(tmp00_93_32), .out(tmp01_46_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004111(.in0(tmp00_94_32), .in1(tmp00_95_32), .out(tmp01_47_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004112(.in0(tmp00_96_32), .in1(tmp00_97_32), .out(tmp01_48_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004113(.in0(tmp00_98_32), .in1(tmp00_99_32), .out(tmp01_49_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004114(.in0(tmp00_100_32), .in1(tmp00_101_32), .out(tmp01_50_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004115(.in0(tmp00_102_32), .in1(tmp00_103_32), .out(tmp01_51_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004116(.in0(tmp00_104_32), .in1(tmp00_105_32), .out(tmp01_52_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004117(.in0(tmp00_106_32), .in1(tmp00_107_32), .out(tmp01_53_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004118(.in0(tmp00_108_32), .in1(tmp00_109_32), .out(tmp01_54_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004119(.in0(tmp00_110_32), .in1(tmp00_111_32), .out(tmp01_55_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004120(.in0(tmp00_112_32), .in1(tmp00_113_32), .out(tmp01_56_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004121(.in0(tmp00_114_32), .in1(tmp00_115_32), .out(tmp01_57_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004122(.in0(tmp00_116_32), .in1(tmp00_117_32), .out(tmp01_58_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004123(.in0(tmp00_118_32), .in1(tmp00_119_32), .out(tmp01_59_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004124(.in0(tmp00_120_32), .in1(tmp00_121_32), .out(tmp01_60_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004125(.in0(tmp00_122_32), .in1(tmp00_123_32), .out(tmp01_61_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004126(.in0(tmp00_124_32), .in1(tmp00_125_32), .out(tmp01_62_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004127(.in0(tmp00_126_32), .in1(tmp00_127_32), .out(tmp01_63_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004128(.in0(tmp01_0_32), .in1(tmp01_1_32), .out(tmp02_0_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004129(.in0(tmp01_2_32), .in1(tmp01_3_32), .out(tmp02_1_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004130(.in0(tmp01_4_32), .in1(tmp01_5_32), .out(tmp02_2_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004131(.in0(tmp01_6_32), .in1(tmp01_7_32), .out(tmp02_3_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004132(.in0(tmp01_8_32), .in1(tmp01_9_32), .out(tmp02_4_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004133(.in0(tmp01_10_32), .in1(tmp01_11_32), .out(tmp02_5_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004134(.in0(tmp01_12_32), .in1(tmp01_13_32), .out(tmp02_6_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004135(.in0(tmp01_14_32), .in1(tmp01_15_32), .out(tmp02_7_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004136(.in0(tmp01_16_32), .in1(tmp01_17_32), .out(tmp02_8_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004137(.in0(tmp01_18_32), .in1(tmp01_19_32), .out(tmp02_9_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004138(.in0(tmp01_20_32), .in1(tmp01_21_32), .out(tmp02_10_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004139(.in0(tmp01_22_32), .in1(tmp01_23_32), .out(tmp02_11_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004140(.in0(tmp01_24_32), .in1(tmp01_25_32), .out(tmp02_12_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004141(.in0(tmp01_26_32), .in1(tmp01_27_32), .out(tmp02_13_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004142(.in0(tmp01_28_32), .in1(tmp01_29_32), .out(tmp02_14_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004143(.in0(tmp01_30_32), .in1(tmp01_31_32), .out(tmp02_15_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004144(.in0(tmp01_32_32), .in1(tmp01_33_32), .out(tmp02_16_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004145(.in0(tmp01_34_32), .in1(tmp01_35_32), .out(tmp02_17_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004146(.in0(tmp01_36_32), .in1(tmp01_37_32), .out(tmp02_18_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004147(.in0(tmp01_38_32), .in1(tmp01_39_32), .out(tmp02_19_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004148(.in0(tmp01_40_32), .in1(tmp01_41_32), .out(tmp02_20_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004149(.in0(tmp01_42_32), .in1(tmp01_43_32), .out(tmp02_21_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004150(.in0(tmp01_44_32), .in1(tmp01_45_32), .out(tmp02_22_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004151(.in0(tmp01_46_32), .in1(tmp01_47_32), .out(tmp02_23_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004152(.in0(tmp01_48_32), .in1(tmp01_49_32), .out(tmp02_24_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004153(.in0(tmp01_50_32), .in1(tmp01_51_32), .out(tmp02_25_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004154(.in0(tmp01_52_32), .in1(tmp01_53_32), .out(tmp02_26_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004155(.in0(tmp01_54_32), .in1(tmp01_55_32), .out(tmp02_27_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004156(.in0(tmp01_56_32), .in1(tmp01_57_32), .out(tmp02_28_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004157(.in0(tmp01_58_32), .in1(tmp01_59_32), .out(tmp02_29_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004158(.in0(tmp01_60_32), .in1(tmp01_61_32), .out(tmp02_30_32));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004159(.in0(tmp01_62_32), .in1(tmp01_63_32), .out(tmp02_31_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004160(.in0(tmp02_0_32), .in1(tmp02_1_32), .out(tmp03_0_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004161(.in0(tmp02_2_32), .in1(tmp02_3_32), .out(tmp03_1_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004162(.in0(tmp02_4_32), .in1(tmp02_5_32), .out(tmp03_2_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004163(.in0(tmp02_6_32), .in1(tmp02_7_32), .out(tmp03_3_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004164(.in0(tmp02_8_32), .in1(tmp02_9_32), .out(tmp03_4_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004165(.in0(tmp02_10_32), .in1(tmp02_11_32), .out(tmp03_5_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004166(.in0(tmp02_12_32), .in1(tmp02_13_32), .out(tmp03_6_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004167(.in0(tmp02_14_32), .in1(tmp02_15_32), .out(tmp03_7_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004168(.in0(tmp02_16_32), .in1(tmp02_17_32), .out(tmp03_8_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004169(.in0(tmp02_18_32), .in1(tmp02_19_32), .out(tmp03_9_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004170(.in0(tmp02_20_32), .in1(tmp02_21_32), .out(tmp03_10_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004171(.in0(tmp02_22_32), .in1(tmp02_23_32), .out(tmp03_11_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004172(.in0(tmp02_24_32), .in1(tmp02_25_32), .out(tmp03_12_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004173(.in0(tmp02_26_32), .in1(tmp02_27_32), .out(tmp03_13_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004174(.in0(tmp02_28_32), .in1(tmp02_29_32), .out(tmp03_14_32));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004175(.in0(tmp02_30_32), .in1(tmp02_31_32), .out(tmp03_15_32));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004176(.in0(tmp03_0_32), .in1(tmp03_1_32), .out(tmp04_0_32));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004177(.in0(tmp03_2_32), .in1(tmp03_3_32), .out(tmp04_1_32));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004178(.in0(tmp03_4_32), .in1(tmp03_5_32), .out(tmp04_2_32));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004179(.in0(tmp03_6_32), .in1(tmp03_7_32), .out(tmp04_3_32));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004180(.in0(tmp03_8_32), .in1(tmp03_9_32), .out(tmp04_4_32));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004181(.in0(tmp03_10_32), .in1(tmp03_11_32), .out(tmp04_5_32));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004182(.in0(tmp03_12_32), .in1(tmp03_13_32), .out(tmp04_6_32));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004183(.in0(tmp03_14_32), .in1(tmp03_15_32), .out(tmp04_7_32));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004184(.in0(tmp04_0_32), .in1(tmp04_1_32), .out(tmp05_0_32));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004185(.in0(tmp04_2_32), .in1(tmp04_3_32), .out(tmp05_1_32));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004186(.in0(tmp04_4_32), .in1(tmp04_5_32), .out(tmp05_2_32));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004187(.in0(tmp04_6_32), .in1(tmp04_7_32), .out(tmp05_3_32));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004188(.in0(tmp05_0_32), .in1(tmp05_1_32), .out(tmp06_0_32));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004189(.in0(tmp05_2_32), .in1(tmp05_3_32), .out(tmp06_1_32));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add004190(.in0(tmp06_0_32), .in1(tmp06_1_32), .out(tmp07_0_32));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004191(.in0(tmp00_0_33), .in1(tmp00_1_33), .out(tmp01_0_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004192(.in0(tmp00_2_33), .in1(tmp00_3_33), .out(tmp01_1_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004193(.in0(tmp00_4_33), .in1(tmp00_5_33), .out(tmp01_2_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004194(.in0(tmp00_6_33), .in1(tmp00_7_33), .out(tmp01_3_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004195(.in0(tmp00_8_33), .in1(tmp00_9_33), .out(tmp01_4_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004196(.in0(tmp00_10_33), .in1(tmp00_11_33), .out(tmp01_5_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004197(.in0(tmp00_12_33), .in1(tmp00_13_33), .out(tmp01_6_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004198(.in0(tmp00_14_33), .in1(tmp00_15_33), .out(tmp01_7_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004199(.in0(tmp00_16_33), .in1(tmp00_17_33), .out(tmp01_8_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004200(.in0(tmp00_18_33), .in1(tmp00_19_33), .out(tmp01_9_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004201(.in0(tmp00_20_33), .in1(tmp00_21_33), .out(tmp01_10_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004202(.in0(tmp00_22_33), .in1(tmp00_23_33), .out(tmp01_11_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004203(.in0(tmp00_24_33), .in1(tmp00_25_33), .out(tmp01_12_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004204(.in0(tmp00_26_33), .in1(tmp00_27_33), .out(tmp01_13_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004205(.in0(tmp00_28_33), .in1(tmp00_29_33), .out(tmp01_14_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004206(.in0(tmp00_30_33), .in1(tmp00_31_33), .out(tmp01_15_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004207(.in0(tmp00_32_33), .in1(tmp00_33_33), .out(tmp01_16_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004208(.in0(tmp00_34_33), .in1(tmp00_35_33), .out(tmp01_17_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004209(.in0(tmp00_36_33), .in1(tmp00_37_33), .out(tmp01_18_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004210(.in0(tmp00_38_33), .in1(tmp00_39_33), .out(tmp01_19_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004211(.in0(tmp00_40_33), .in1(tmp00_41_33), .out(tmp01_20_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004212(.in0(tmp00_42_33), .in1(tmp00_43_33), .out(tmp01_21_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004213(.in0(tmp00_44_33), .in1(tmp00_45_33), .out(tmp01_22_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004214(.in0(tmp00_46_33), .in1(tmp00_47_33), .out(tmp01_23_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004215(.in0(tmp00_48_33), .in1(tmp00_49_33), .out(tmp01_24_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004216(.in0(tmp00_50_33), .in1(tmp00_51_33), .out(tmp01_25_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004217(.in0(tmp00_52_33), .in1(tmp00_53_33), .out(tmp01_26_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004218(.in0(tmp00_54_33), .in1(tmp00_55_33), .out(tmp01_27_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004219(.in0(tmp00_56_33), .in1(tmp00_57_33), .out(tmp01_28_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004220(.in0(tmp00_58_33), .in1(tmp00_59_33), .out(tmp01_29_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004221(.in0(tmp00_60_33), .in1(tmp00_61_33), .out(tmp01_30_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004222(.in0(tmp00_62_33), .in1(tmp00_63_33), .out(tmp01_31_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004223(.in0(tmp00_64_33), .in1(tmp00_65_33), .out(tmp01_32_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004224(.in0(tmp00_66_33), .in1(tmp00_67_33), .out(tmp01_33_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004225(.in0(tmp00_68_33), .in1(tmp00_69_33), .out(tmp01_34_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004226(.in0(tmp00_70_33), .in1(tmp00_71_33), .out(tmp01_35_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004227(.in0(tmp00_72_33), .in1(tmp00_73_33), .out(tmp01_36_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004228(.in0(tmp00_74_33), .in1(tmp00_75_33), .out(tmp01_37_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004229(.in0(tmp00_76_33), .in1(tmp00_77_33), .out(tmp01_38_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004230(.in0(tmp00_78_33), .in1(tmp00_79_33), .out(tmp01_39_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004231(.in0(tmp00_80_33), .in1(tmp00_81_33), .out(tmp01_40_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004232(.in0(tmp00_82_33), .in1(tmp00_83_33), .out(tmp01_41_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004233(.in0(tmp00_84_33), .in1(tmp00_85_33), .out(tmp01_42_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004234(.in0(tmp00_86_33), .in1(tmp00_87_33), .out(tmp01_43_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004235(.in0(tmp00_88_33), .in1(tmp00_89_33), .out(tmp01_44_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004236(.in0(tmp00_90_33), .in1(tmp00_91_33), .out(tmp01_45_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004237(.in0(tmp00_92_33), .in1(tmp00_93_33), .out(tmp01_46_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004238(.in0(tmp00_94_33), .in1(tmp00_95_33), .out(tmp01_47_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004239(.in0(tmp00_96_33), .in1(tmp00_97_33), .out(tmp01_48_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004240(.in0(tmp00_98_33), .in1(tmp00_99_33), .out(tmp01_49_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004241(.in0(tmp00_100_33), .in1(tmp00_101_33), .out(tmp01_50_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004242(.in0(tmp00_102_33), .in1(tmp00_103_33), .out(tmp01_51_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004243(.in0(tmp00_104_33), .in1(tmp00_105_33), .out(tmp01_52_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004244(.in0(tmp00_106_33), .in1(tmp00_107_33), .out(tmp01_53_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004245(.in0(tmp00_108_33), .in1(tmp00_109_33), .out(tmp01_54_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004246(.in0(tmp00_110_33), .in1(tmp00_111_33), .out(tmp01_55_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004247(.in0(tmp00_112_33), .in1(tmp00_113_33), .out(tmp01_56_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004248(.in0(tmp00_114_33), .in1(tmp00_115_33), .out(tmp01_57_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004249(.in0(tmp00_116_33), .in1(tmp00_117_33), .out(tmp01_58_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004250(.in0(tmp00_118_33), .in1(tmp00_119_33), .out(tmp01_59_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004251(.in0(tmp00_120_33), .in1(tmp00_121_33), .out(tmp01_60_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004252(.in0(tmp00_122_33), .in1(tmp00_123_33), .out(tmp01_61_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004253(.in0(tmp00_124_33), .in1(tmp00_125_33), .out(tmp01_62_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004254(.in0(tmp00_126_33), .in1(tmp00_127_33), .out(tmp01_63_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004255(.in0(tmp01_0_33), .in1(tmp01_1_33), .out(tmp02_0_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004256(.in0(tmp01_2_33), .in1(tmp01_3_33), .out(tmp02_1_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004257(.in0(tmp01_4_33), .in1(tmp01_5_33), .out(tmp02_2_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004258(.in0(tmp01_6_33), .in1(tmp01_7_33), .out(tmp02_3_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004259(.in0(tmp01_8_33), .in1(tmp01_9_33), .out(tmp02_4_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004260(.in0(tmp01_10_33), .in1(tmp01_11_33), .out(tmp02_5_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004261(.in0(tmp01_12_33), .in1(tmp01_13_33), .out(tmp02_6_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004262(.in0(tmp01_14_33), .in1(tmp01_15_33), .out(tmp02_7_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004263(.in0(tmp01_16_33), .in1(tmp01_17_33), .out(tmp02_8_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004264(.in0(tmp01_18_33), .in1(tmp01_19_33), .out(tmp02_9_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004265(.in0(tmp01_20_33), .in1(tmp01_21_33), .out(tmp02_10_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004266(.in0(tmp01_22_33), .in1(tmp01_23_33), .out(tmp02_11_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004267(.in0(tmp01_24_33), .in1(tmp01_25_33), .out(tmp02_12_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004268(.in0(tmp01_26_33), .in1(tmp01_27_33), .out(tmp02_13_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004269(.in0(tmp01_28_33), .in1(tmp01_29_33), .out(tmp02_14_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004270(.in0(tmp01_30_33), .in1(tmp01_31_33), .out(tmp02_15_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004271(.in0(tmp01_32_33), .in1(tmp01_33_33), .out(tmp02_16_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004272(.in0(tmp01_34_33), .in1(tmp01_35_33), .out(tmp02_17_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004273(.in0(tmp01_36_33), .in1(tmp01_37_33), .out(tmp02_18_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004274(.in0(tmp01_38_33), .in1(tmp01_39_33), .out(tmp02_19_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004275(.in0(tmp01_40_33), .in1(tmp01_41_33), .out(tmp02_20_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004276(.in0(tmp01_42_33), .in1(tmp01_43_33), .out(tmp02_21_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004277(.in0(tmp01_44_33), .in1(tmp01_45_33), .out(tmp02_22_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004278(.in0(tmp01_46_33), .in1(tmp01_47_33), .out(tmp02_23_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004279(.in0(tmp01_48_33), .in1(tmp01_49_33), .out(tmp02_24_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004280(.in0(tmp01_50_33), .in1(tmp01_51_33), .out(tmp02_25_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004281(.in0(tmp01_52_33), .in1(tmp01_53_33), .out(tmp02_26_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004282(.in0(tmp01_54_33), .in1(tmp01_55_33), .out(tmp02_27_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004283(.in0(tmp01_56_33), .in1(tmp01_57_33), .out(tmp02_28_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004284(.in0(tmp01_58_33), .in1(tmp01_59_33), .out(tmp02_29_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004285(.in0(tmp01_60_33), .in1(tmp01_61_33), .out(tmp02_30_33));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004286(.in0(tmp01_62_33), .in1(tmp01_63_33), .out(tmp02_31_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004287(.in0(tmp02_0_33), .in1(tmp02_1_33), .out(tmp03_0_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004288(.in0(tmp02_2_33), .in1(tmp02_3_33), .out(tmp03_1_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004289(.in0(tmp02_4_33), .in1(tmp02_5_33), .out(tmp03_2_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004290(.in0(tmp02_6_33), .in1(tmp02_7_33), .out(tmp03_3_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004291(.in0(tmp02_8_33), .in1(tmp02_9_33), .out(tmp03_4_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004292(.in0(tmp02_10_33), .in1(tmp02_11_33), .out(tmp03_5_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004293(.in0(tmp02_12_33), .in1(tmp02_13_33), .out(tmp03_6_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004294(.in0(tmp02_14_33), .in1(tmp02_15_33), .out(tmp03_7_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004295(.in0(tmp02_16_33), .in1(tmp02_17_33), .out(tmp03_8_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004296(.in0(tmp02_18_33), .in1(tmp02_19_33), .out(tmp03_9_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004297(.in0(tmp02_20_33), .in1(tmp02_21_33), .out(tmp03_10_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004298(.in0(tmp02_22_33), .in1(tmp02_23_33), .out(tmp03_11_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004299(.in0(tmp02_24_33), .in1(tmp02_25_33), .out(tmp03_12_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004300(.in0(tmp02_26_33), .in1(tmp02_27_33), .out(tmp03_13_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004301(.in0(tmp02_28_33), .in1(tmp02_29_33), .out(tmp03_14_33));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004302(.in0(tmp02_30_33), .in1(tmp02_31_33), .out(tmp03_15_33));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004303(.in0(tmp03_0_33), .in1(tmp03_1_33), .out(tmp04_0_33));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004304(.in0(tmp03_2_33), .in1(tmp03_3_33), .out(tmp04_1_33));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004305(.in0(tmp03_4_33), .in1(tmp03_5_33), .out(tmp04_2_33));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004306(.in0(tmp03_6_33), .in1(tmp03_7_33), .out(tmp04_3_33));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004307(.in0(tmp03_8_33), .in1(tmp03_9_33), .out(tmp04_4_33));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004308(.in0(tmp03_10_33), .in1(tmp03_11_33), .out(tmp04_5_33));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004309(.in0(tmp03_12_33), .in1(tmp03_13_33), .out(tmp04_6_33));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004310(.in0(tmp03_14_33), .in1(tmp03_15_33), .out(tmp04_7_33));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004311(.in0(tmp04_0_33), .in1(tmp04_1_33), .out(tmp05_0_33));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004312(.in0(tmp04_2_33), .in1(tmp04_3_33), .out(tmp05_1_33));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004313(.in0(tmp04_4_33), .in1(tmp04_5_33), .out(tmp05_2_33));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004314(.in0(tmp04_6_33), .in1(tmp04_7_33), .out(tmp05_3_33));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004315(.in0(tmp05_0_33), .in1(tmp05_1_33), .out(tmp06_0_33));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004316(.in0(tmp05_2_33), .in1(tmp05_3_33), .out(tmp06_1_33));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add004317(.in0(tmp06_0_33), .in1(tmp06_1_33), .out(tmp07_0_33));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004318(.in0(tmp00_0_34), .in1(tmp00_1_34), .out(tmp01_0_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004319(.in0(tmp00_2_34), .in1(tmp00_3_34), .out(tmp01_1_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004320(.in0(tmp00_4_34), .in1(tmp00_5_34), .out(tmp01_2_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004321(.in0(tmp00_6_34), .in1(tmp00_7_34), .out(tmp01_3_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004322(.in0(tmp00_8_34), .in1(tmp00_9_34), .out(tmp01_4_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004323(.in0(tmp00_10_34), .in1(tmp00_11_34), .out(tmp01_5_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004324(.in0(tmp00_12_34), .in1(tmp00_13_34), .out(tmp01_6_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004325(.in0(tmp00_14_34), .in1(tmp00_15_34), .out(tmp01_7_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004326(.in0(tmp00_16_34), .in1(tmp00_17_34), .out(tmp01_8_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004327(.in0(tmp00_18_34), .in1(tmp00_19_34), .out(tmp01_9_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004328(.in0(tmp00_20_34), .in1(tmp00_21_34), .out(tmp01_10_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004329(.in0(tmp00_22_34), .in1(tmp00_23_34), .out(tmp01_11_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004330(.in0(tmp00_24_34), .in1(tmp00_25_34), .out(tmp01_12_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004331(.in0(tmp00_26_34), .in1(tmp00_27_34), .out(tmp01_13_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004332(.in0(tmp00_28_34), .in1(tmp00_29_34), .out(tmp01_14_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004333(.in0(tmp00_30_34), .in1(tmp00_31_34), .out(tmp01_15_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004334(.in0(tmp00_32_34), .in1(tmp00_33_34), .out(tmp01_16_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004335(.in0(tmp00_34_34), .in1(tmp00_35_34), .out(tmp01_17_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004336(.in0(tmp00_36_34), .in1(tmp00_37_34), .out(tmp01_18_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004337(.in0(tmp00_38_34), .in1(tmp00_39_34), .out(tmp01_19_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004338(.in0(tmp00_40_34), .in1(tmp00_41_34), .out(tmp01_20_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004339(.in0(tmp00_42_34), .in1(tmp00_43_34), .out(tmp01_21_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004340(.in0(tmp00_44_34), .in1(tmp00_45_34), .out(tmp01_22_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004341(.in0(tmp00_46_34), .in1(tmp00_47_34), .out(tmp01_23_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004342(.in0(tmp00_48_34), .in1(tmp00_49_34), .out(tmp01_24_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004343(.in0(tmp00_50_34), .in1(tmp00_51_34), .out(tmp01_25_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004344(.in0(tmp00_52_34), .in1(tmp00_53_34), .out(tmp01_26_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004345(.in0(tmp00_54_34), .in1(tmp00_55_34), .out(tmp01_27_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004346(.in0(tmp00_56_34), .in1(tmp00_57_34), .out(tmp01_28_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004347(.in0(tmp00_58_34), .in1(tmp00_59_34), .out(tmp01_29_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004348(.in0(tmp00_60_34), .in1(tmp00_61_34), .out(tmp01_30_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004349(.in0(tmp00_62_34), .in1(tmp00_63_34), .out(tmp01_31_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004350(.in0(tmp00_64_34), .in1(tmp00_65_34), .out(tmp01_32_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004351(.in0(tmp00_66_34), .in1(tmp00_67_34), .out(tmp01_33_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004352(.in0(tmp00_68_34), .in1(tmp00_69_34), .out(tmp01_34_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004353(.in0(tmp00_70_34), .in1(tmp00_71_34), .out(tmp01_35_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004354(.in0(tmp00_72_34), .in1(tmp00_73_34), .out(tmp01_36_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004355(.in0(tmp00_74_34), .in1(tmp00_75_34), .out(tmp01_37_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004356(.in0(tmp00_76_34), .in1(tmp00_77_34), .out(tmp01_38_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004357(.in0(tmp00_78_34), .in1(tmp00_79_34), .out(tmp01_39_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004358(.in0(tmp00_80_34), .in1(tmp00_81_34), .out(tmp01_40_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004359(.in0(tmp00_82_34), .in1(tmp00_83_34), .out(tmp01_41_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004360(.in0(tmp00_84_34), .in1(tmp00_85_34), .out(tmp01_42_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004361(.in0(tmp00_86_34), .in1(tmp00_87_34), .out(tmp01_43_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004362(.in0(tmp00_88_34), .in1(tmp00_89_34), .out(tmp01_44_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004363(.in0(tmp00_90_34), .in1(tmp00_91_34), .out(tmp01_45_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004364(.in0(tmp00_92_34), .in1(tmp00_93_34), .out(tmp01_46_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004365(.in0(tmp00_94_34), .in1(tmp00_95_34), .out(tmp01_47_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004366(.in0(tmp00_96_34), .in1(tmp00_97_34), .out(tmp01_48_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004367(.in0(tmp00_98_34), .in1(tmp00_99_34), .out(tmp01_49_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004368(.in0(tmp00_100_34), .in1(tmp00_101_34), .out(tmp01_50_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004369(.in0(tmp00_102_34), .in1(tmp00_103_34), .out(tmp01_51_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004370(.in0(tmp00_104_34), .in1(tmp00_105_34), .out(tmp01_52_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004371(.in0(tmp00_106_34), .in1(tmp00_107_34), .out(tmp01_53_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004372(.in0(tmp00_108_34), .in1(tmp00_109_34), .out(tmp01_54_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004373(.in0(tmp00_110_34), .in1(tmp00_111_34), .out(tmp01_55_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004374(.in0(tmp00_112_34), .in1(tmp00_113_34), .out(tmp01_56_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004375(.in0(tmp00_114_34), .in1(tmp00_115_34), .out(tmp01_57_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004376(.in0(tmp00_116_34), .in1(tmp00_117_34), .out(tmp01_58_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004377(.in0(tmp00_118_34), .in1(tmp00_119_34), .out(tmp01_59_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004378(.in0(tmp00_120_34), .in1(tmp00_121_34), .out(tmp01_60_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004379(.in0(tmp00_122_34), .in1(tmp00_123_34), .out(tmp01_61_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004380(.in0(tmp00_124_34), .in1(tmp00_125_34), .out(tmp01_62_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004381(.in0(tmp00_126_34), .in1(tmp00_127_34), .out(tmp01_63_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004382(.in0(tmp01_0_34), .in1(tmp01_1_34), .out(tmp02_0_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004383(.in0(tmp01_2_34), .in1(tmp01_3_34), .out(tmp02_1_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004384(.in0(tmp01_4_34), .in1(tmp01_5_34), .out(tmp02_2_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004385(.in0(tmp01_6_34), .in1(tmp01_7_34), .out(tmp02_3_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004386(.in0(tmp01_8_34), .in1(tmp01_9_34), .out(tmp02_4_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004387(.in0(tmp01_10_34), .in1(tmp01_11_34), .out(tmp02_5_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004388(.in0(tmp01_12_34), .in1(tmp01_13_34), .out(tmp02_6_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004389(.in0(tmp01_14_34), .in1(tmp01_15_34), .out(tmp02_7_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004390(.in0(tmp01_16_34), .in1(tmp01_17_34), .out(tmp02_8_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004391(.in0(tmp01_18_34), .in1(tmp01_19_34), .out(tmp02_9_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004392(.in0(tmp01_20_34), .in1(tmp01_21_34), .out(tmp02_10_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004393(.in0(tmp01_22_34), .in1(tmp01_23_34), .out(tmp02_11_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004394(.in0(tmp01_24_34), .in1(tmp01_25_34), .out(tmp02_12_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004395(.in0(tmp01_26_34), .in1(tmp01_27_34), .out(tmp02_13_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004396(.in0(tmp01_28_34), .in1(tmp01_29_34), .out(tmp02_14_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004397(.in0(tmp01_30_34), .in1(tmp01_31_34), .out(tmp02_15_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004398(.in0(tmp01_32_34), .in1(tmp01_33_34), .out(tmp02_16_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004399(.in0(tmp01_34_34), .in1(tmp01_35_34), .out(tmp02_17_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004400(.in0(tmp01_36_34), .in1(tmp01_37_34), .out(tmp02_18_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004401(.in0(tmp01_38_34), .in1(tmp01_39_34), .out(tmp02_19_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004402(.in0(tmp01_40_34), .in1(tmp01_41_34), .out(tmp02_20_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004403(.in0(tmp01_42_34), .in1(tmp01_43_34), .out(tmp02_21_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004404(.in0(tmp01_44_34), .in1(tmp01_45_34), .out(tmp02_22_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004405(.in0(tmp01_46_34), .in1(tmp01_47_34), .out(tmp02_23_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004406(.in0(tmp01_48_34), .in1(tmp01_49_34), .out(tmp02_24_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004407(.in0(tmp01_50_34), .in1(tmp01_51_34), .out(tmp02_25_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004408(.in0(tmp01_52_34), .in1(tmp01_53_34), .out(tmp02_26_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004409(.in0(tmp01_54_34), .in1(tmp01_55_34), .out(tmp02_27_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004410(.in0(tmp01_56_34), .in1(tmp01_57_34), .out(tmp02_28_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004411(.in0(tmp01_58_34), .in1(tmp01_59_34), .out(tmp02_29_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004412(.in0(tmp01_60_34), .in1(tmp01_61_34), .out(tmp02_30_34));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004413(.in0(tmp01_62_34), .in1(tmp01_63_34), .out(tmp02_31_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004414(.in0(tmp02_0_34), .in1(tmp02_1_34), .out(tmp03_0_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004415(.in0(tmp02_2_34), .in1(tmp02_3_34), .out(tmp03_1_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004416(.in0(tmp02_4_34), .in1(tmp02_5_34), .out(tmp03_2_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004417(.in0(tmp02_6_34), .in1(tmp02_7_34), .out(tmp03_3_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004418(.in0(tmp02_8_34), .in1(tmp02_9_34), .out(tmp03_4_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004419(.in0(tmp02_10_34), .in1(tmp02_11_34), .out(tmp03_5_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004420(.in0(tmp02_12_34), .in1(tmp02_13_34), .out(tmp03_6_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004421(.in0(tmp02_14_34), .in1(tmp02_15_34), .out(tmp03_7_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004422(.in0(tmp02_16_34), .in1(tmp02_17_34), .out(tmp03_8_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004423(.in0(tmp02_18_34), .in1(tmp02_19_34), .out(tmp03_9_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004424(.in0(tmp02_20_34), .in1(tmp02_21_34), .out(tmp03_10_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004425(.in0(tmp02_22_34), .in1(tmp02_23_34), .out(tmp03_11_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004426(.in0(tmp02_24_34), .in1(tmp02_25_34), .out(tmp03_12_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004427(.in0(tmp02_26_34), .in1(tmp02_27_34), .out(tmp03_13_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004428(.in0(tmp02_28_34), .in1(tmp02_29_34), .out(tmp03_14_34));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004429(.in0(tmp02_30_34), .in1(tmp02_31_34), .out(tmp03_15_34));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004430(.in0(tmp03_0_34), .in1(tmp03_1_34), .out(tmp04_0_34));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004431(.in0(tmp03_2_34), .in1(tmp03_3_34), .out(tmp04_1_34));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004432(.in0(tmp03_4_34), .in1(tmp03_5_34), .out(tmp04_2_34));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004433(.in0(tmp03_6_34), .in1(tmp03_7_34), .out(tmp04_3_34));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004434(.in0(tmp03_8_34), .in1(tmp03_9_34), .out(tmp04_4_34));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004435(.in0(tmp03_10_34), .in1(tmp03_11_34), .out(tmp04_5_34));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004436(.in0(tmp03_12_34), .in1(tmp03_13_34), .out(tmp04_6_34));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004437(.in0(tmp03_14_34), .in1(tmp03_15_34), .out(tmp04_7_34));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004438(.in0(tmp04_0_34), .in1(tmp04_1_34), .out(tmp05_0_34));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004439(.in0(tmp04_2_34), .in1(tmp04_3_34), .out(tmp05_1_34));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004440(.in0(tmp04_4_34), .in1(tmp04_5_34), .out(tmp05_2_34));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004441(.in0(tmp04_6_34), .in1(tmp04_7_34), .out(tmp05_3_34));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004442(.in0(tmp05_0_34), .in1(tmp05_1_34), .out(tmp06_0_34));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004443(.in0(tmp05_2_34), .in1(tmp05_3_34), .out(tmp06_1_34));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add004444(.in0(tmp06_0_34), .in1(tmp06_1_34), .out(tmp07_0_34));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004445(.in0(tmp00_0_35), .in1(tmp00_1_35), .out(tmp01_0_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004446(.in0(tmp00_2_35), .in1(tmp00_3_35), .out(tmp01_1_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004447(.in0(tmp00_4_35), .in1(tmp00_5_35), .out(tmp01_2_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004448(.in0(tmp00_6_35), .in1(tmp00_7_35), .out(tmp01_3_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004449(.in0(tmp00_8_35), .in1(tmp00_9_35), .out(tmp01_4_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004450(.in0(tmp00_10_35), .in1(tmp00_11_35), .out(tmp01_5_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004451(.in0(tmp00_12_35), .in1(tmp00_13_35), .out(tmp01_6_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004452(.in0(tmp00_14_35), .in1(tmp00_15_35), .out(tmp01_7_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004453(.in0(tmp00_16_35), .in1(tmp00_17_35), .out(tmp01_8_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004454(.in0(tmp00_18_35), .in1(tmp00_19_35), .out(tmp01_9_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004455(.in0(tmp00_20_35), .in1(tmp00_21_35), .out(tmp01_10_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004456(.in0(tmp00_22_35), .in1(tmp00_23_35), .out(tmp01_11_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004457(.in0(tmp00_24_35), .in1(tmp00_25_35), .out(tmp01_12_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004458(.in0(tmp00_26_35), .in1(tmp00_27_35), .out(tmp01_13_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004459(.in0(tmp00_28_35), .in1(tmp00_29_35), .out(tmp01_14_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004460(.in0(tmp00_30_35), .in1(tmp00_31_35), .out(tmp01_15_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004461(.in0(tmp00_32_35), .in1(tmp00_33_35), .out(tmp01_16_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004462(.in0(tmp00_34_35), .in1(tmp00_35_35), .out(tmp01_17_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004463(.in0(tmp00_36_35), .in1(tmp00_37_35), .out(tmp01_18_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004464(.in0(tmp00_38_35), .in1(tmp00_39_35), .out(tmp01_19_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004465(.in0(tmp00_40_35), .in1(tmp00_41_35), .out(tmp01_20_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004466(.in0(tmp00_42_35), .in1(tmp00_43_35), .out(tmp01_21_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004467(.in0(tmp00_44_35), .in1(tmp00_45_35), .out(tmp01_22_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004468(.in0(tmp00_46_35), .in1(tmp00_47_35), .out(tmp01_23_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004469(.in0(tmp00_48_35), .in1(tmp00_49_35), .out(tmp01_24_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004470(.in0(tmp00_50_35), .in1(tmp00_51_35), .out(tmp01_25_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004471(.in0(tmp00_52_35), .in1(tmp00_53_35), .out(tmp01_26_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004472(.in0(tmp00_54_35), .in1(tmp00_55_35), .out(tmp01_27_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004473(.in0(tmp00_56_35), .in1(tmp00_57_35), .out(tmp01_28_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004474(.in0(tmp00_58_35), .in1(tmp00_59_35), .out(tmp01_29_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004475(.in0(tmp00_60_35), .in1(tmp00_61_35), .out(tmp01_30_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004476(.in0(tmp00_62_35), .in1(tmp00_63_35), .out(tmp01_31_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004477(.in0(tmp00_64_35), .in1(tmp00_65_35), .out(tmp01_32_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004478(.in0(tmp00_66_35), .in1(tmp00_67_35), .out(tmp01_33_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004479(.in0(tmp00_68_35), .in1(tmp00_69_35), .out(tmp01_34_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004480(.in0(tmp00_70_35), .in1(tmp00_71_35), .out(tmp01_35_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004481(.in0(tmp00_72_35), .in1(tmp00_73_35), .out(tmp01_36_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004482(.in0(tmp00_74_35), .in1(tmp00_75_35), .out(tmp01_37_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004483(.in0(tmp00_76_35), .in1(tmp00_77_35), .out(tmp01_38_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004484(.in0(tmp00_78_35), .in1(tmp00_79_35), .out(tmp01_39_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004485(.in0(tmp00_80_35), .in1(tmp00_81_35), .out(tmp01_40_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004486(.in0(tmp00_82_35), .in1(tmp00_83_35), .out(tmp01_41_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004487(.in0(tmp00_84_35), .in1(tmp00_85_35), .out(tmp01_42_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004488(.in0(tmp00_86_35), .in1(tmp00_87_35), .out(tmp01_43_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004489(.in0(tmp00_88_35), .in1(tmp00_89_35), .out(tmp01_44_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004490(.in0(tmp00_90_35), .in1(tmp00_91_35), .out(tmp01_45_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004491(.in0(tmp00_92_35), .in1(tmp00_93_35), .out(tmp01_46_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004492(.in0(tmp00_94_35), .in1(tmp00_95_35), .out(tmp01_47_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004493(.in0(tmp00_96_35), .in1(tmp00_97_35), .out(tmp01_48_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004494(.in0(tmp00_98_35), .in1(tmp00_99_35), .out(tmp01_49_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004495(.in0(tmp00_100_35), .in1(tmp00_101_35), .out(tmp01_50_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004496(.in0(tmp00_102_35), .in1(tmp00_103_35), .out(tmp01_51_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004497(.in0(tmp00_104_35), .in1(tmp00_105_35), .out(tmp01_52_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004498(.in0(tmp00_106_35), .in1(tmp00_107_35), .out(tmp01_53_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004499(.in0(tmp00_108_35), .in1(tmp00_109_35), .out(tmp01_54_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004500(.in0(tmp00_110_35), .in1(tmp00_111_35), .out(tmp01_55_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004501(.in0(tmp00_112_35), .in1(tmp00_113_35), .out(tmp01_56_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004502(.in0(tmp00_114_35), .in1(tmp00_115_35), .out(tmp01_57_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004503(.in0(tmp00_116_35), .in1(tmp00_117_35), .out(tmp01_58_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004504(.in0(tmp00_118_35), .in1(tmp00_119_35), .out(tmp01_59_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004505(.in0(tmp00_120_35), .in1(tmp00_121_35), .out(tmp01_60_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004506(.in0(tmp00_122_35), .in1(tmp00_123_35), .out(tmp01_61_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004507(.in0(tmp00_124_35), .in1(tmp00_125_35), .out(tmp01_62_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004508(.in0(tmp00_126_35), .in1(tmp00_127_35), .out(tmp01_63_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004509(.in0(tmp01_0_35), .in1(tmp01_1_35), .out(tmp02_0_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004510(.in0(tmp01_2_35), .in1(tmp01_3_35), .out(tmp02_1_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004511(.in0(tmp01_4_35), .in1(tmp01_5_35), .out(tmp02_2_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004512(.in0(tmp01_6_35), .in1(tmp01_7_35), .out(tmp02_3_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004513(.in0(tmp01_8_35), .in1(tmp01_9_35), .out(tmp02_4_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004514(.in0(tmp01_10_35), .in1(tmp01_11_35), .out(tmp02_5_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004515(.in0(tmp01_12_35), .in1(tmp01_13_35), .out(tmp02_6_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004516(.in0(tmp01_14_35), .in1(tmp01_15_35), .out(tmp02_7_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004517(.in0(tmp01_16_35), .in1(tmp01_17_35), .out(tmp02_8_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004518(.in0(tmp01_18_35), .in1(tmp01_19_35), .out(tmp02_9_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004519(.in0(tmp01_20_35), .in1(tmp01_21_35), .out(tmp02_10_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004520(.in0(tmp01_22_35), .in1(tmp01_23_35), .out(tmp02_11_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004521(.in0(tmp01_24_35), .in1(tmp01_25_35), .out(tmp02_12_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004522(.in0(tmp01_26_35), .in1(tmp01_27_35), .out(tmp02_13_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004523(.in0(tmp01_28_35), .in1(tmp01_29_35), .out(tmp02_14_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004524(.in0(tmp01_30_35), .in1(tmp01_31_35), .out(tmp02_15_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004525(.in0(tmp01_32_35), .in1(tmp01_33_35), .out(tmp02_16_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004526(.in0(tmp01_34_35), .in1(tmp01_35_35), .out(tmp02_17_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004527(.in0(tmp01_36_35), .in1(tmp01_37_35), .out(tmp02_18_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004528(.in0(tmp01_38_35), .in1(tmp01_39_35), .out(tmp02_19_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004529(.in0(tmp01_40_35), .in1(tmp01_41_35), .out(tmp02_20_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004530(.in0(tmp01_42_35), .in1(tmp01_43_35), .out(tmp02_21_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004531(.in0(tmp01_44_35), .in1(tmp01_45_35), .out(tmp02_22_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004532(.in0(tmp01_46_35), .in1(tmp01_47_35), .out(tmp02_23_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004533(.in0(tmp01_48_35), .in1(tmp01_49_35), .out(tmp02_24_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004534(.in0(tmp01_50_35), .in1(tmp01_51_35), .out(tmp02_25_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004535(.in0(tmp01_52_35), .in1(tmp01_53_35), .out(tmp02_26_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004536(.in0(tmp01_54_35), .in1(tmp01_55_35), .out(tmp02_27_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004537(.in0(tmp01_56_35), .in1(tmp01_57_35), .out(tmp02_28_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004538(.in0(tmp01_58_35), .in1(tmp01_59_35), .out(tmp02_29_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004539(.in0(tmp01_60_35), .in1(tmp01_61_35), .out(tmp02_30_35));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004540(.in0(tmp01_62_35), .in1(tmp01_63_35), .out(tmp02_31_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004541(.in0(tmp02_0_35), .in1(tmp02_1_35), .out(tmp03_0_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004542(.in0(tmp02_2_35), .in1(tmp02_3_35), .out(tmp03_1_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004543(.in0(tmp02_4_35), .in1(tmp02_5_35), .out(tmp03_2_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004544(.in0(tmp02_6_35), .in1(tmp02_7_35), .out(tmp03_3_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004545(.in0(tmp02_8_35), .in1(tmp02_9_35), .out(tmp03_4_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004546(.in0(tmp02_10_35), .in1(tmp02_11_35), .out(tmp03_5_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004547(.in0(tmp02_12_35), .in1(tmp02_13_35), .out(tmp03_6_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004548(.in0(tmp02_14_35), .in1(tmp02_15_35), .out(tmp03_7_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004549(.in0(tmp02_16_35), .in1(tmp02_17_35), .out(tmp03_8_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004550(.in0(tmp02_18_35), .in1(tmp02_19_35), .out(tmp03_9_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004551(.in0(tmp02_20_35), .in1(tmp02_21_35), .out(tmp03_10_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004552(.in0(tmp02_22_35), .in1(tmp02_23_35), .out(tmp03_11_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004553(.in0(tmp02_24_35), .in1(tmp02_25_35), .out(tmp03_12_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004554(.in0(tmp02_26_35), .in1(tmp02_27_35), .out(tmp03_13_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004555(.in0(tmp02_28_35), .in1(tmp02_29_35), .out(tmp03_14_35));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004556(.in0(tmp02_30_35), .in1(tmp02_31_35), .out(tmp03_15_35));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004557(.in0(tmp03_0_35), .in1(tmp03_1_35), .out(tmp04_0_35));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004558(.in0(tmp03_2_35), .in1(tmp03_3_35), .out(tmp04_1_35));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004559(.in0(tmp03_4_35), .in1(tmp03_5_35), .out(tmp04_2_35));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004560(.in0(tmp03_6_35), .in1(tmp03_7_35), .out(tmp04_3_35));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004561(.in0(tmp03_8_35), .in1(tmp03_9_35), .out(tmp04_4_35));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004562(.in0(tmp03_10_35), .in1(tmp03_11_35), .out(tmp04_5_35));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004563(.in0(tmp03_12_35), .in1(tmp03_13_35), .out(tmp04_6_35));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004564(.in0(tmp03_14_35), .in1(tmp03_15_35), .out(tmp04_7_35));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004565(.in0(tmp04_0_35), .in1(tmp04_1_35), .out(tmp05_0_35));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004566(.in0(tmp04_2_35), .in1(tmp04_3_35), .out(tmp05_1_35));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004567(.in0(tmp04_4_35), .in1(tmp04_5_35), .out(tmp05_2_35));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004568(.in0(tmp04_6_35), .in1(tmp04_7_35), .out(tmp05_3_35));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004569(.in0(tmp05_0_35), .in1(tmp05_1_35), .out(tmp06_0_35));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004570(.in0(tmp05_2_35), .in1(tmp05_3_35), .out(tmp06_1_35));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add004571(.in0(tmp06_0_35), .in1(tmp06_1_35), .out(tmp07_0_35));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004572(.in0(tmp00_0_36), .in1(tmp00_1_36), .out(tmp01_0_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004573(.in0(tmp00_2_36), .in1(tmp00_3_36), .out(tmp01_1_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004574(.in0(tmp00_4_36), .in1(tmp00_5_36), .out(tmp01_2_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004575(.in0(tmp00_6_36), .in1(tmp00_7_36), .out(tmp01_3_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004576(.in0(tmp00_8_36), .in1(tmp00_9_36), .out(tmp01_4_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004577(.in0(tmp00_10_36), .in1(tmp00_11_36), .out(tmp01_5_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004578(.in0(tmp00_12_36), .in1(tmp00_13_36), .out(tmp01_6_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004579(.in0(tmp00_14_36), .in1(tmp00_15_36), .out(tmp01_7_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004580(.in0(tmp00_16_36), .in1(tmp00_17_36), .out(tmp01_8_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004581(.in0(tmp00_18_36), .in1(tmp00_19_36), .out(tmp01_9_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004582(.in0(tmp00_20_36), .in1(tmp00_21_36), .out(tmp01_10_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004583(.in0(tmp00_22_36), .in1(tmp00_23_36), .out(tmp01_11_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004584(.in0(tmp00_24_36), .in1(tmp00_25_36), .out(tmp01_12_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004585(.in0(tmp00_26_36), .in1(tmp00_27_36), .out(tmp01_13_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004586(.in0(tmp00_28_36), .in1(tmp00_29_36), .out(tmp01_14_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004587(.in0(tmp00_30_36), .in1(tmp00_31_36), .out(tmp01_15_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004588(.in0(tmp00_32_36), .in1(tmp00_33_36), .out(tmp01_16_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004589(.in0(tmp00_34_36), .in1(tmp00_35_36), .out(tmp01_17_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004590(.in0(tmp00_36_36), .in1(tmp00_37_36), .out(tmp01_18_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004591(.in0(tmp00_38_36), .in1(tmp00_39_36), .out(tmp01_19_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004592(.in0(tmp00_40_36), .in1(tmp00_41_36), .out(tmp01_20_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004593(.in0(tmp00_42_36), .in1(tmp00_43_36), .out(tmp01_21_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004594(.in0(tmp00_44_36), .in1(tmp00_45_36), .out(tmp01_22_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004595(.in0(tmp00_46_36), .in1(tmp00_47_36), .out(tmp01_23_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004596(.in0(tmp00_48_36), .in1(tmp00_49_36), .out(tmp01_24_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004597(.in0(tmp00_50_36), .in1(tmp00_51_36), .out(tmp01_25_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004598(.in0(tmp00_52_36), .in1(tmp00_53_36), .out(tmp01_26_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004599(.in0(tmp00_54_36), .in1(tmp00_55_36), .out(tmp01_27_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004600(.in0(tmp00_56_36), .in1(tmp00_57_36), .out(tmp01_28_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004601(.in0(tmp00_58_36), .in1(tmp00_59_36), .out(tmp01_29_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004602(.in0(tmp00_60_36), .in1(tmp00_61_36), .out(tmp01_30_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004603(.in0(tmp00_62_36), .in1(tmp00_63_36), .out(tmp01_31_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004604(.in0(tmp00_64_36), .in1(tmp00_65_36), .out(tmp01_32_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004605(.in0(tmp00_66_36), .in1(tmp00_67_36), .out(tmp01_33_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004606(.in0(tmp00_68_36), .in1(tmp00_69_36), .out(tmp01_34_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004607(.in0(tmp00_70_36), .in1(tmp00_71_36), .out(tmp01_35_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004608(.in0(tmp00_72_36), .in1(tmp00_73_36), .out(tmp01_36_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004609(.in0(tmp00_74_36), .in1(tmp00_75_36), .out(tmp01_37_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004610(.in0(tmp00_76_36), .in1(tmp00_77_36), .out(tmp01_38_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004611(.in0(tmp00_78_36), .in1(tmp00_79_36), .out(tmp01_39_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004612(.in0(tmp00_80_36), .in1(tmp00_81_36), .out(tmp01_40_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004613(.in0(tmp00_82_36), .in1(tmp00_83_36), .out(tmp01_41_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004614(.in0(tmp00_84_36), .in1(tmp00_85_36), .out(tmp01_42_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004615(.in0(tmp00_86_36), .in1(tmp00_87_36), .out(tmp01_43_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004616(.in0(tmp00_88_36), .in1(tmp00_89_36), .out(tmp01_44_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004617(.in0(tmp00_90_36), .in1(tmp00_91_36), .out(tmp01_45_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004618(.in0(tmp00_92_36), .in1(tmp00_93_36), .out(tmp01_46_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004619(.in0(tmp00_94_36), .in1(tmp00_95_36), .out(tmp01_47_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004620(.in0(tmp00_96_36), .in1(tmp00_97_36), .out(tmp01_48_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004621(.in0(tmp00_98_36), .in1(tmp00_99_36), .out(tmp01_49_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004622(.in0(tmp00_100_36), .in1(tmp00_101_36), .out(tmp01_50_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004623(.in0(tmp00_102_36), .in1(tmp00_103_36), .out(tmp01_51_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004624(.in0(tmp00_104_36), .in1(tmp00_105_36), .out(tmp01_52_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004625(.in0(tmp00_106_36), .in1(tmp00_107_36), .out(tmp01_53_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004626(.in0(tmp00_108_36), .in1(tmp00_109_36), .out(tmp01_54_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004627(.in0(tmp00_110_36), .in1(tmp00_111_36), .out(tmp01_55_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004628(.in0(tmp00_112_36), .in1(tmp00_113_36), .out(tmp01_56_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004629(.in0(tmp00_114_36), .in1(tmp00_115_36), .out(tmp01_57_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004630(.in0(tmp00_116_36), .in1(tmp00_117_36), .out(tmp01_58_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004631(.in0(tmp00_118_36), .in1(tmp00_119_36), .out(tmp01_59_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004632(.in0(tmp00_120_36), .in1(tmp00_121_36), .out(tmp01_60_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004633(.in0(tmp00_122_36), .in1(tmp00_123_36), .out(tmp01_61_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004634(.in0(tmp00_124_36), .in1(tmp00_125_36), .out(tmp01_62_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004635(.in0(tmp00_126_36), .in1(tmp00_127_36), .out(tmp01_63_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004636(.in0(tmp01_0_36), .in1(tmp01_1_36), .out(tmp02_0_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004637(.in0(tmp01_2_36), .in1(tmp01_3_36), .out(tmp02_1_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004638(.in0(tmp01_4_36), .in1(tmp01_5_36), .out(tmp02_2_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004639(.in0(tmp01_6_36), .in1(tmp01_7_36), .out(tmp02_3_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004640(.in0(tmp01_8_36), .in1(tmp01_9_36), .out(tmp02_4_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004641(.in0(tmp01_10_36), .in1(tmp01_11_36), .out(tmp02_5_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004642(.in0(tmp01_12_36), .in1(tmp01_13_36), .out(tmp02_6_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004643(.in0(tmp01_14_36), .in1(tmp01_15_36), .out(tmp02_7_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004644(.in0(tmp01_16_36), .in1(tmp01_17_36), .out(tmp02_8_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004645(.in0(tmp01_18_36), .in1(tmp01_19_36), .out(tmp02_9_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004646(.in0(tmp01_20_36), .in1(tmp01_21_36), .out(tmp02_10_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004647(.in0(tmp01_22_36), .in1(tmp01_23_36), .out(tmp02_11_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004648(.in0(tmp01_24_36), .in1(tmp01_25_36), .out(tmp02_12_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004649(.in0(tmp01_26_36), .in1(tmp01_27_36), .out(tmp02_13_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004650(.in0(tmp01_28_36), .in1(tmp01_29_36), .out(tmp02_14_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004651(.in0(tmp01_30_36), .in1(tmp01_31_36), .out(tmp02_15_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004652(.in0(tmp01_32_36), .in1(tmp01_33_36), .out(tmp02_16_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004653(.in0(tmp01_34_36), .in1(tmp01_35_36), .out(tmp02_17_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004654(.in0(tmp01_36_36), .in1(tmp01_37_36), .out(tmp02_18_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004655(.in0(tmp01_38_36), .in1(tmp01_39_36), .out(tmp02_19_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004656(.in0(tmp01_40_36), .in1(tmp01_41_36), .out(tmp02_20_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004657(.in0(tmp01_42_36), .in1(tmp01_43_36), .out(tmp02_21_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004658(.in0(tmp01_44_36), .in1(tmp01_45_36), .out(tmp02_22_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004659(.in0(tmp01_46_36), .in1(tmp01_47_36), .out(tmp02_23_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004660(.in0(tmp01_48_36), .in1(tmp01_49_36), .out(tmp02_24_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004661(.in0(tmp01_50_36), .in1(tmp01_51_36), .out(tmp02_25_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004662(.in0(tmp01_52_36), .in1(tmp01_53_36), .out(tmp02_26_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004663(.in0(tmp01_54_36), .in1(tmp01_55_36), .out(tmp02_27_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004664(.in0(tmp01_56_36), .in1(tmp01_57_36), .out(tmp02_28_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004665(.in0(tmp01_58_36), .in1(tmp01_59_36), .out(tmp02_29_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004666(.in0(tmp01_60_36), .in1(tmp01_61_36), .out(tmp02_30_36));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004667(.in0(tmp01_62_36), .in1(tmp01_63_36), .out(tmp02_31_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004668(.in0(tmp02_0_36), .in1(tmp02_1_36), .out(tmp03_0_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004669(.in0(tmp02_2_36), .in1(tmp02_3_36), .out(tmp03_1_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004670(.in0(tmp02_4_36), .in1(tmp02_5_36), .out(tmp03_2_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004671(.in0(tmp02_6_36), .in1(tmp02_7_36), .out(tmp03_3_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004672(.in0(tmp02_8_36), .in1(tmp02_9_36), .out(tmp03_4_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004673(.in0(tmp02_10_36), .in1(tmp02_11_36), .out(tmp03_5_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004674(.in0(tmp02_12_36), .in1(tmp02_13_36), .out(tmp03_6_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004675(.in0(tmp02_14_36), .in1(tmp02_15_36), .out(tmp03_7_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004676(.in0(tmp02_16_36), .in1(tmp02_17_36), .out(tmp03_8_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004677(.in0(tmp02_18_36), .in1(tmp02_19_36), .out(tmp03_9_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004678(.in0(tmp02_20_36), .in1(tmp02_21_36), .out(tmp03_10_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004679(.in0(tmp02_22_36), .in1(tmp02_23_36), .out(tmp03_11_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004680(.in0(tmp02_24_36), .in1(tmp02_25_36), .out(tmp03_12_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004681(.in0(tmp02_26_36), .in1(tmp02_27_36), .out(tmp03_13_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004682(.in0(tmp02_28_36), .in1(tmp02_29_36), .out(tmp03_14_36));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004683(.in0(tmp02_30_36), .in1(tmp02_31_36), .out(tmp03_15_36));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004684(.in0(tmp03_0_36), .in1(tmp03_1_36), .out(tmp04_0_36));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004685(.in0(tmp03_2_36), .in1(tmp03_3_36), .out(tmp04_1_36));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004686(.in0(tmp03_4_36), .in1(tmp03_5_36), .out(tmp04_2_36));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004687(.in0(tmp03_6_36), .in1(tmp03_7_36), .out(tmp04_3_36));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004688(.in0(tmp03_8_36), .in1(tmp03_9_36), .out(tmp04_4_36));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004689(.in0(tmp03_10_36), .in1(tmp03_11_36), .out(tmp04_5_36));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004690(.in0(tmp03_12_36), .in1(tmp03_13_36), .out(tmp04_6_36));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004691(.in0(tmp03_14_36), .in1(tmp03_15_36), .out(tmp04_7_36));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004692(.in0(tmp04_0_36), .in1(tmp04_1_36), .out(tmp05_0_36));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004693(.in0(tmp04_2_36), .in1(tmp04_3_36), .out(tmp05_1_36));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004694(.in0(tmp04_4_36), .in1(tmp04_5_36), .out(tmp05_2_36));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004695(.in0(tmp04_6_36), .in1(tmp04_7_36), .out(tmp05_3_36));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004696(.in0(tmp05_0_36), .in1(tmp05_1_36), .out(tmp06_0_36));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004697(.in0(tmp05_2_36), .in1(tmp05_3_36), .out(tmp06_1_36));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add004698(.in0(tmp06_0_36), .in1(tmp06_1_36), .out(tmp07_0_36));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004699(.in0(tmp00_0_37), .in1(tmp00_1_37), .out(tmp01_0_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004700(.in0(tmp00_2_37), .in1(tmp00_3_37), .out(tmp01_1_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004701(.in0(tmp00_4_37), .in1(tmp00_5_37), .out(tmp01_2_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004702(.in0(tmp00_6_37), .in1(tmp00_7_37), .out(tmp01_3_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004703(.in0(tmp00_8_37), .in1(tmp00_9_37), .out(tmp01_4_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004704(.in0(tmp00_10_37), .in1(tmp00_11_37), .out(tmp01_5_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004705(.in0(tmp00_12_37), .in1(tmp00_13_37), .out(tmp01_6_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004706(.in0(tmp00_14_37), .in1(tmp00_15_37), .out(tmp01_7_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004707(.in0(tmp00_16_37), .in1(tmp00_17_37), .out(tmp01_8_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004708(.in0(tmp00_18_37), .in1(tmp00_19_37), .out(tmp01_9_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004709(.in0(tmp00_20_37), .in1(tmp00_21_37), .out(tmp01_10_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004710(.in0(tmp00_22_37), .in1(tmp00_23_37), .out(tmp01_11_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004711(.in0(tmp00_24_37), .in1(tmp00_25_37), .out(tmp01_12_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004712(.in0(tmp00_26_37), .in1(tmp00_27_37), .out(tmp01_13_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004713(.in0(tmp00_28_37), .in1(tmp00_29_37), .out(tmp01_14_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004714(.in0(tmp00_30_37), .in1(tmp00_31_37), .out(tmp01_15_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004715(.in0(tmp00_32_37), .in1(tmp00_33_37), .out(tmp01_16_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004716(.in0(tmp00_34_37), .in1(tmp00_35_37), .out(tmp01_17_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004717(.in0(tmp00_36_37), .in1(tmp00_37_37), .out(tmp01_18_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004718(.in0(tmp00_38_37), .in1(tmp00_39_37), .out(tmp01_19_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004719(.in0(tmp00_40_37), .in1(tmp00_41_37), .out(tmp01_20_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004720(.in0(tmp00_42_37), .in1(tmp00_43_37), .out(tmp01_21_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004721(.in0(tmp00_44_37), .in1(tmp00_45_37), .out(tmp01_22_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004722(.in0(tmp00_46_37), .in1(tmp00_47_37), .out(tmp01_23_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004723(.in0(tmp00_48_37), .in1(tmp00_49_37), .out(tmp01_24_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004724(.in0(tmp00_50_37), .in1(tmp00_51_37), .out(tmp01_25_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004725(.in0(tmp00_52_37), .in1(tmp00_53_37), .out(tmp01_26_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004726(.in0(tmp00_54_37), .in1(tmp00_55_37), .out(tmp01_27_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004727(.in0(tmp00_56_37), .in1(tmp00_57_37), .out(tmp01_28_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004728(.in0(tmp00_58_37), .in1(tmp00_59_37), .out(tmp01_29_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004729(.in0(tmp00_60_37), .in1(tmp00_61_37), .out(tmp01_30_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004730(.in0(tmp00_62_37), .in1(tmp00_63_37), .out(tmp01_31_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004731(.in0(tmp00_64_37), .in1(tmp00_65_37), .out(tmp01_32_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004732(.in0(tmp00_66_37), .in1(tmp00_67_37), .out(tmp01_33_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004733(.in0(tmp00_68_37), .in1(tmp00_69_37), .out(tmp01_34_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004734(.in0(tmp00_70_37), .in1(tmp00_71_37), .out(tmp01_35_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004735(.in0(tmp00_72_37), .in1(tmp00_73_37), .out(tmp01_36_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004736(.in0(tmp00_74_37), .in1(tmp00_75_37), .out(tmp01_37_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004737(.in0(tmp00_76_37), .in1(tmp00_77_37), .out(tmp01_38_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004738(.in0(tmp00_78_37), .in1(tmp00_79_37), .out(tmp01_39_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004739(.in0(tmp00_80_37), .in1(tmp00_81_37), .out(tmp01_40_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004740(.in0(tmp00_82_37), .in1(tmp00_83_37), .out(tmp01_41_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004741(.in0(tmp00_84_37), .in1(tmp00_85_37), .out(tmp01_42_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004742(.in0(tmp00_86_37), .in1(tmp00_87_37), .out(tmp01_43_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004743(.in0(tmp00_88_37), .in1(tmp00_89_37), .out(tmp01_44_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004744(.in0(tmp00_90_37), .in1(tmp00_91_37), .out(tmp01_45_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004745(.in0(tmp00_92_37), .in1(tmp00_93_37), .out(tmp01_46_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004746(.in0(tmp00_94_37), .in1(tmp00_95_37), .out(tmp01_47_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004747(.in0(tmp00_96_37), .in1(tmp00_97_37), .out(tmp01_48_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004748(.in0(tmp00_98_37), .in1(tmp00_99_37), .out(tmp01_49_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004749(.in0(tmp00_100_37), .in1(tmp00_101_37), .out(tmp01_50_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004750(.in0(tmp00_102_37), .in1(tmp00_103_37), .out(tmp01_51_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004751(.in0(tmp00_104_37), .in1(tmp00_105_37), .out(tmp01_52_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004752(.in0(tmp00_106_37), .in1(tmp00_107_37), .out(tmp01_53_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004753(.in0(tmp00_108_37), .in1(tmp00_109_37), .out(tmp01_54_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004754(.in0(tmp00_110_37), .in1(tmp00_111_37), .out(tmp01_55_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004755(.in0(tmp00_112_37), .in1(tmp00_113_37), .out(tmp01_56_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004756(.in0(tmp00_114_37), .in1(tmp00_115_37), .out(tmp01_57_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004757(.in0(tmp00_116_37), .in1(tmp00_117_37), .out(tmp01_58_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004758(.in0(tmp00_118_37), .in1(tmp00_119_37), .out(tmp01_59_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004759(.in0(tmp00_120_37), .in1(tmp00_121_37), .out(tmp01_60_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004760(.in0(tmp00_122_37), .in1(tmp00_123_37), .out(tmp01_61_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004761(.in0(tmp00_124_37), .in1(tmp00_125_37), .out(tmp01_62_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004762(.in0(tmp00_126_37), .in1(tmp00_127_37), .out(tmp01_63_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004763(.in0(tmp01_0_37), .in1(tmp01_1_37), .out(tmp02_0_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004764(.in0(tmp01_2_37), .in1(tmp01_3_37), .out(tmp02_1_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004765(.in0(tmp01_4_37), .in1(tmp01_5_37), .out(tmp02_2_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004766(.in0(tmp01_6_37), .in1(tmp01_7_37), .out(tmp02_3_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004767(.in0(tmp01_8_37), .in1(tmp01_9_37), .out(tmp02_4_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004768(.in0(tmp01_10_37), .in1(tmp01_11_37), .out(tmp02_5_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004769(.in0(tmp01_12_37), .in1(tmp01_13_37), .out(tmp02_6_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004770(.in0(tmp01_14_37), .in1(tmp01_15_37), .out(tmp02_7_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004771(.in0(tmp01_16_37), .in1(tmp01_17_37), .out(tmp02_8_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004772(.in0(tmp01_18_37), .in1(tmp01_19_37), .out(tmp02_9_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004773(.in0(tmp01_20_37), .in1(tmp01_21_37), .out(tmp02_10_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004774(.in0(tmp01_22_37), .in1(tmp01_23_37), .out(tmp02_11_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004775(.in0(tmp01_24_37), .in1(tmp01_25_37), .out(tmp02_12_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004776(.in0(tmp01_26_37), .in1(tmp01_27_37), .out(tmp02_13_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004777(.in0(tmp01_28_37), .in1(tmp01_29_37), .out(tmp02_14_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004778(.in0(tmp01_30_37), .in1(tmp01_31_37), .out(tmp02_15_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004779(.in0(tmp01_32_37), .in1(tmp01_33_37), .out(tmp02_16_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004780(.in0(tmp01_34_37), .in1(tmp01_35_37), .out(tmp02_17_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004781(.in0(tmp01_36_37), .in1(tmp01_37_37), .out(tmp02_18_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004782(.in0(tmp01_38_37), .in1(tmp01_39_37), .out(tmp02_19_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004783(.in0(tmp01_40_37), .in1(tmp01_41_37), .out(tmp02_20_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004784(.in0(tmp01_42_37), .in1(tmp01_43_37), .out(tmp02_21_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004785(.in0(tmp01_44_37), .in1(tmp01_45_37), .out(tmp02_22_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004786(.in0(tmp01_46_37), .in1(tmp01_47_37), .out(tmp02_23_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004787(.in0(tmp01_48_37), .in1(tmp01_49_37), .out(tmp02_24_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004788(.in0(tmp01_50_37), .in1(tmp01_51_37), .out(tmp02_25_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004789(.in0(tmp01_52_37), .in1(tmp01_53_37), .out(tmp02_26_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004790(.in0(tmp01_54_37), .in1(tmp01_55_37), .out(tmp02_27_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004791(.in0(tmp01_56_37), .in1(tmp01_57_37), .out(tmp02_28_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004792(.in0(tmp01_58_37), .in1(tmp01_59_37), .out(tmp02_29_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004793(.in0(tmp01_60_37), .in1(tmp01_61_37), .out(tmp02_30_37));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004794(.in0(tmp01_62_37), .in1(tmp01_63_37), .out(tmp02_31_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004795(.in0(tmp02_0_37), .in1(tmp02_1_37), .out(tmp03_0_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004796(.in0(tmp02_2_37), .in1(tmp02_3_37), .out(tmp03_1_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004797(.in0(tmp02_4_37), .in1(tmp02_5_37), .out(tmp03_2_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004798(.in0(tmp02_6_37), .in1(tmp02_7_37), .out(tmp03_3_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004799(.in0(tmp02_8_37), .in1(tmp02_9_37), .out(tmp03_4_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004800(.in0(tmp02_10_37), .in1(tmp02_11_37), .out(tmp03_5_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004801(.in0(tmp02_12_37), .in1(tmp02_13_37), .out(tmp03_6_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004802(.in0(tmp02_14_37), .in1(tmp02_15_37), .out(tmp03_7_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004803(.in0(tmp02_16_37), .in1(tmp02_17_37), .out(tmp03_8_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004804(.in0(tmp02_18_37), .in1(tmp02_19_37), .out(tmp03_9_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004805(.in0(tmp02_20_37), .in1(tmp02_21_37), .out(tmp03_10_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004806(.in0(tmp02_22_37), .in1(tmp02_23_37), .out(tmp03_11_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004807(.in0(tmp02_24_37), .in1(tmp02_25_37), .out(tmp03_12_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004808(.in0(tmp02_26_37), .in1(tmp02_27_37), .out(tmp03_13_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004809(.in0(tmp02_28_37), .in1(tmp02_29_37), .out(tmp03_14_37));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004810(.in0(tmp02_30_37), .in1(tmp02_31_37), .out(tmp03_15_37));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004811(.in0(tmp03_0_37), .in1(tmp03_1_37), .out(tmp04_0_37));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004812(.in0(tmp03_2_37), .in1(tmp03_3_37), .out(tmp04_1_37));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004813(.in0(tmp03_4_37), .in1(tmp03_5_37), .out(tmp04_2_37));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004814(.in0(tmp03_6_37), .in1(tmp03_7_37), .out(tmp04_3_37));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004815(.in0(tmp03_8_37), .in1(tmp03_9_37), .out(tmp04_4_37));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004816(.in0(tmp03_10_37), .in1(tmp03_11_37), .out(tmp04_5_37));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004817(.in0(tmp03_12_37), .in1(tmp03_13_37), .out(tmp04_6_37));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004818(.in0(tmp03_14_37), .in1(tmp03_15_37), .out(tmp04_7_37));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004819(.in0(tmp04_0_37), .in1(tmp04_1_37), .out(tmp05_0_37));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004820(.in0(tmp04_2_37), .in1(tmp04_3_37), .out(tmp05_1_37));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004821(.in0(tmp04_4_37), .in1(tmp04_5_37), .out(tmp05_2_37));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004822(.in0(tmp04_6_37), .in1(tmp04_7_37), .out(tmp05_3_37));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004823(.in0(tmp05_0_37), .in1(tmp05_1_37), .out(tmp06_0_37));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004824(.in0(tmp05_2_37), .in1(tmp05_3_37), .out(tmp06_1_37));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add004825(.in0(tmp06_0_37), .in1(tmp06_1_37), .out(tmp07_0_37));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004826(.in0(tmp00_0_38), .in1(tmp00_1_38), .out(tmp01_0_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004827(.in0(tmp00_2_38), .in1(tmp00_3_38), .out(tmp01_1_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004828(.in0(tmp00_4_38), .in1(tmp00_5_38), .out(tmp01_2_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004829(.in0(tmp00_6_38), .in1(tmp00_7_38), .out(tmp01_3_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004830(.in0(tmp00_8_38), .in1(tmp00_9_38), .out(tmp01_4_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004831(.in0(tmp00_10_38), .in1(tmp00_11_38), .out(tmp01_5_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004832(.in0(tmp00_12_38), .in1(tmp00_13_38), .out(tmp01_6_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004833(.in0(tmp00_14_38), .in1(tmp00_15_38), .out(tmp01_7_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004834(.in0(tmp00_16_38), .in1(tmp00_17_38), .out(tmp01_8_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004835(.in0(tmp00_18_38), .in1(tmp00_19_38), .out(tmp01_9_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004836(.in0(tmp00_20_38), .in1(tmp00_21_38), .out(tmp01_10_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004837(.in0(tmp00_22_38), .in1(tmp00_23_38), .out(tmp01_11_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004838(.in0(tmp00_24_38), .in1(tmp00_25_38), .out(tmp01_12_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004839(.in0(tmp00_26_38), .in1(tmp00_27_38), .out(tmp01_13_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004840(.in0(tmp00_28_38), .in1(tmp00_29_38), .out(tmp01_14_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004841(.in0(tmp00_30_38), .in1(tmp00_31_38), .out(tmp01_15_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004842(.in0(tmp00_32_38), .in1(tmp00_33_38), .out(tmp01_16_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004843(.in0(tmp00_34_38), .in1(tmp00_35_38), .out(tmp01_17_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004844(.in0(tmp00_36_38), .in1(tmp00_37_38), .out(tmp01_18_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004845(.in0(tmp00_38_38), .in1(tmp00_39_38), .out(tmp01_19_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004846(.in0(tmp00_40_38), .in1(tmp00_41_38), .out(tmp01_20_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004847(.in0(tmp00_42_38), .in1(tmp00_43_38), .out(tmp01_21_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004848(.in0(tmp00_44_38), .in1(tmp00_45_38), .out(tmp01_22_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004849(.in0(tmp00_46_38), .in1(tmp00_47_38), .out(tmp01_23_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004850(.in0(tmp00_48_38), .in1(tmp00_49_38), .out(tmp01_24_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004851(.in0(tmp00_50_38), .in1(tmp00_51_38), .out(tmp01_25_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004852(.in0(tmp00_52_38), .in1(tmp00_53_38), .out(tmp01_26_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004853(.in0(tmp00_54_38), .in1(tmp00_55_38), .out(tmp01_27_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004854(.in0(tmp00_56_38), .in1(tmp00_57_38), .out(tmp01_28_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004855(.in0(tmp00_58_38), .in1(tmp00_59_38), .out(tmp01_29_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004856(.in0(tmp00_60_38), .in1(tmp00_61_38), .out(tmp01_30_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004857(.in0(tmp00_62_38), .in1(tmp00_63_38), .out(tmp01_31_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004858(.in0(tmp00_64_38), .in1(tmp00_65_38), .out(tmp01_32_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004859(.in0(tmp00_66_38), .in1(tmp00_67_38), .out(tmp01_33_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004860(.in0(tmp00_68_38), .in1(tmp00_69_38), .out(tmp01_34_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004861(.in0(tmp00_70_38), .in1(tmp00_71_38), .out(tmp01_35_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004862(.in0(tmp00_72_38), .in1(tmp00_73_38), .out(tmp01_36_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004863(.in0(tmp00_74_38), .in1(tmp00_75_38), .out(tmp01_37_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004864(.in0(tmp00_76_38), .in1(tmp00_77_38), .out(tmp01_38_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004865(.in0(tmp00_78_38), .in1(tmp00_79_38), .out(tmp01_39_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004866(.in0(tmp00_80_38), .in1(tmp00_81_38), .out(tmp01_40_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004867(.in0(tmp00_82_38), .in1(tmp00_83_38), .out(tmp01_41_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004868(.in0(tmp00_84_38), .in1(tmp00_85_38), .out(tmp01_42_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004869(.in0(tmp00_86_38), .in1(tmp00_87_38), .out(tmp01_43_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004870(.in0(tmp00_88_38), .in1(tmp00_89_38), .out(tmp01_44_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004871(.in0(tmp00_90_38), .in1(tmp00_91_38), .out(tmp01_45_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004872(.in0(tmp00_92_38), .in1(tmp00_93_38), .out(tmp01_46_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004873(.in0(tmp00_94_38), .in1(tmp00_95_38), .out(tmp01_47_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004874(.in0(tmp00_96_38), .in1(tmp00_97_38), .out(tmp01_48_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004875(.in0(tmp00_98_38), .in1(tmp00_99_38), .out(tmp01_49_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004876(.in0(tmp00_100_38), .in1(tmp00_101_38), .out(tmp01_50_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004877(.in0(tmp00_102_38), .in1(tmp00_103_38), .out(tmp01_51_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004878(.in0(tmp00_104_38), .in1(tmp00_105_38), .out(tmp01_52_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004879(.in0(tmp00_106_38), .in1(tmp00_107_38), .out(tmp01_53_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004880(.in0(tmp00_108_38), .in1(tmp00_109_38), .out(tmp01_54_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004881(.in0(tmp00_110_38), .in1(tmp00_111_38), .out(tmp01_55_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004882(.in0(tmp00_112_38), .in1(tmp00_113_38), .out(tmp01_56_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004883(.in0(tmp00_114_38), .in1(tmp00_115_38), .out(tmp01_57_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004884(.in0(tmp00_116_38), .in1(tmp00_117_38), .out(tmp01_58_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004885(.in0(tmp00_118_38), .in1(tmp00_119_38), .out(tmp01_59_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004886(.in0(tmp00_120_38), .in1(tmp00_121_38), .out(tmp01_60_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004887(.in0(tmp00_122_38), .in1(tmp00_123_38), .out(tmp01_61_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004888(.in0(tmp00_124_38), .in1(tmp00_125_38), .out(tmp01_62_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004889(.in0(tmp00_126_38), .in1(tmp00_127_38), .out(tmp01_63_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004890(.in0(tmp01_0_38), .in1(tmp01_1_38), .out(tmp02_0_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004891(.in0(tmp01_2_38), .in1(tmp01_3_38), .out(tmp02_1_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004892(.in0(tmp01_4_38), .in1(tmp01_5_38), .out(tmp02_2_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004893(.in0(tmp01_6_38), .in1(tmp01_7_38), .out(tmp02_3_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004894(.in0(tmp01_8_38), .in1(tmp01_9_38), .out(tmp02_4_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004895(.in0(tmp01_10_38), .in1(tmp01_11_38), .out(tmp02_5_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004896(.in0(tmp01_12_38), .in1(tmp01_13_38), .out(tmp02_6_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004897(.in0(tmp01_14_38), .in1(tmp01_15_38), .out(tmp02_7_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004898(.in0(tmp01_16_38), .in1(tmp01_17_38), .out(tmp02_8_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004899(.in0(tmp01_18_38), .in1(tmp01_19_38), .out(tmp02_9_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004900(.in0(tmp01_20_38), .in1(tmp01_21_38), .out(tmp02_10_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004901(.in0(tmp01_22_38), .in1(tmp01_23_38), .out(tmp02_11_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004902(.in0(tmp01_24_38), .in1(tmp01_25_38), .out(tmp02_12_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004903(.in0(tmp01_26_38), .in1(tmp01_27_38), .out(tmp02_13_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004904(.in0(tmp01_28_38), .in1(tmp01_29_38), .out(tmp02_14_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004905(.in0(tmp01_30_38), .in1(tmp01_31_38), .out(tmp02_15_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004906(.in0(tmp01_32_38), .in1(tmp01_33_38), .out(tmp02_16_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004907(.in0(tmp01_34_38), .in1(tmp01_35_38), .out(tmp02_17_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004908(.in0(tmp01_36_38), .in1(tmp01_37_38), .out(tmp02_18_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004909(.in0(tmp01_38_38), .in1(tmp01_39_38), .out(tmp02_19_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004910(.in0(tmp01_40_38), .in1(tmp01_41_38), .out(tmp02_20_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004911(.in0(tmp01_42_38), .in1(tmp01_43_38), .out(tmp02_21_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004912(.in0(tmp01_44_38), .in1(tmp01_45_38), .out(tmp02_22_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004913(.in0(tmp01_46_38), .in1(tmp01_47_38), .out(tmp02_23_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004914(.in0(tmp01_48_38), .in1(tmp01_49_38), .out(tmp02_24_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004915(.in0(tmp01_50_38), .in1(tmp01_51_38), .out(tmp02_25_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004916(.in0(tmp01_52_38), .in1(tmp01_53_38), .out(tmp02_26_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004917(.in0(tmp01_54_38), .in1(tmp01_55_38), .out(tmp02_27_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004918(.in0(tmp01_56_38), .in1(tmp01_57_38), .out(tmp02_28_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004919(.in0(tmp01_58_38), .in1(tmp01_59_38), .out(tmp02_29_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004920(.in0(tmp01_60_38), .in1(tmp01_61_38), .out(tmp02_30_38));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add004921(.in0(tmp01_62_38), .in1(tmp01_63_38), .out(tmp02_31_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004922(.in0(tmp02_0_38), .in1(tmp02_1_38), .out(tmp03_0_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004923(.in0(tmp02_2_38), .in1(tmp02_3_38), .out(tmp03_1_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004924(.in0(tmp02_4_38), .in1(tmp02_5_38), .out(tmp03_2_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004925(.in0(tmp02_6_38), .in1(tmp02_7_38), .out(tmp03_3_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004926(.in0(tmp02_8_38), .in1(tmp02_9_38), .out(tmp03_4_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004927(.in0(tmp02_10_38), .in1(tmp02_11_38), .out(tmp03_5_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004928(.in0(tmp02_12_38), .in1(tmp02_13_38), .out(tmp03_6_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004929(.in0(tmp02_14_38), .in1(tmp02_15_38), .out(tmp03_7_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004930(.in0(tmp02_16_38), .in1(tmp02_17_38), .out(tmp03_8_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004931(.in0(tmp02_18_38), .in1(tmp02_19_38), .out(tmp03_9_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004932(.in0(tmp02_20_38), .in1(tmp02_21_38), .out(tmp03_10_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004933(.in0(tmp02_22_38), .in1(tmp02_23_38), .out(tmp03_11_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004934(.in0(tmp02_24_38), .in1(tmp02_25_38), .out(tmp03_12_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004935(.in0(tmp02_26_38), .in1(tmp02_27_38), .out(tmp03_13_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004936(.in0(tmp02_28_38), .in1(tmp02_29_38), .out(tmp03_14_38));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add004937(.in0(tmp02_30_38), .in1(tmp02_31_38), .out(tmp03_15_38));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004938(.in0(tmp03_0_38), .in1(tmp03_1_38), .out(tmp04_0_38));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004939(.in0(tmp03_2_38), .in1(tmp03_3_38), .out(tmp04_1_38));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004940(.in0(tmp03_4_38), .in1(tmp03_5_38), .out(tmp04_2_38));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004941(.in0(tmp03_6_38), .in1(tmp03_7_38), .out(tmp04_3_38));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004942(.in0(tmp03_8_38), .in1(tmp03_9_38), .out(tmp04_4_38));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004943(.in0(tmp03_10_38), .in1(tmp03_11_38), .out(tmp04_5_38));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004944(.in0(tmp03_12_38), .in1(tmp03_13_38), .out(tmp04_6_38));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add004945(.in0(tmp03_14_38), .in1(tmp03_15_38), .out(tmp04_7_38));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004946(.in0(tmp04_0_38), .in1(tmp04_1_38), .out(tmp05_0_38));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004947(.in0(tmp04_2_38), .in1(tmp04_3_38), .out(tmp05_1_38));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004948(.in0(tmp04_4_38), .in1(tmp04_5_38), .out(tmp05_2_38));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add004949(.in0(tmp04_6_38), .in1(tmp04_7_38), .out(tmp05_3_38));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004950(.in0(tmp05_0_38), .in1(tmp05_1_38), .out(tmp06_0_38));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add004951(.in0(tmp05_2_38), .in1(tmp05_3_38), .out(tmp06_1_38));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add004952(.in0(tmp06_0_38), .in1(tmp06_1_38), .out(tmp07_0_38));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004953(.in0(tmp00_0_39), .in1(tmp00_1_39), .out(tmp01_0_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004954(.in0(tmp00_2_39), .in1(tmp00_3_39), .out(tmp01_1_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004955(.in0(tmp00_4_39), .in1(tmp00_5_39), .out(tmp01_2_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004956(.in0(tmp00_6_39), .in1(tmp00_7_39), .out(tmp01_3_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004957(.in0(tmp00_8_39), .in1(tmp00_9_39), .out(tmp01_4_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004958(.in0(tmp00_10_39), .in1(tmp00_11_39), .out(tmp01_5_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004959(.in0(tmp00_12_39), .in1(tmp00_13_39), .out(tmp01_6_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004960(.in0(tmp00_14_39), .in1(tmp00_15_39), .out(tmp01_7_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004961(.in0(tmp00_16_39), .in1(tmp00_17_39), .out(tmp01_8_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004962(.in0(tmp00_18_39), .in1(tmp00_19_39), .out(tmp01_9_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004963(.in0(tmp00_20_39), .in1(tmp00_21_39), .out(tmp01_10_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004964(.in0(tmp00_22_39), .in1(tmp00_23_39), .out(tmp01_11_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004965(.in0(tmp00_24_39), .in1(tmp00_25_39), .out(tmp01_12_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004966(.in0(tmp00_26_39), .in1(tmp00_27_39), .out(tmp01_13_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004967(.in0(tmp00_28_39), .in1(tmp00_29_39), .out(tmp01_14_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004968(.in0(tmp00_30_39), .in1(tmp00_31_39), .out(tmp01_15_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004969(.in0(tmp00_32_39), .in1(tmp00_33_39), .out(tmp01_16_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004970(.in0(tmp00_34_39), .in1(tmp00_35_39), .out(tmp01_17_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004971(.in0(tmp00_36_39), .in1(tmp00_37_39), .out(tmp01_18_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004972(.in0(tmp00_38_39), .in1(tmp00_39_39), .out(tmp01_19_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004973(.in0(tmp00_40_39), .in1(tmp00_41_39), .out(tmp01_20_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004974(.in0(tmp00_42_39), .in1(tmp00_43_39), .out(tmp01_21_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004975(.in0(tmp00_44_39), .in1(tmp00_45_39), .out(tmp01_22_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004976(.in0(tmp00_46_39), .in1(tmp00_47_39), .out(tmp01_23_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004977(.in0(tmp00_48_39), .in1(tmp00_49_39), .out(tmp01_24_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004978(.in0(tmp00_50_39), .in1(tmp00_51_39), .out(tmp01_25_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004979(.in0(tmp00_52_39), .in1(tmp00_53_39), .out(tmp01_26_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004980(.in0(tmp00_54_39), .in1(tmp00_55_39), .out(tmp01_27_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004981(.in0(tmp00_56_39), .in1(tmp00_57_39), .out(tmp01_28_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004982(.in0(tmp00_58_39), .in1(tmp00_59_39), .out(tmp01_29_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004983(.in0(tmp00_60_39), .in1(tmp00_61_39), .out(tmp01_30_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004984(.in0(tmp00_62_39), .in1(tmp00_63_39), .out(tmp01_31_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004985(.in0(tmp00_64_39), .in1(tmp00_65_39), .out(tmp01_32_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004986(.in0(tmp00_66_39), .in1(tmp00_67_39), .out(tmp01_33_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004987(.in0(tmp00_68_39), .in1(tmp00_69_39), .out(tmp01_34_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004988(.in0(tmp00_70_39), .in1(tmp00_71_39), .out(tmp01_35_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004989(.in0(tmp00_72_39), .in1(tmp00_73_39), .out(tmp01_36_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004990(.in0(tmp00_74_39), .in1(tmp00_75_39), .out(tmp01_37_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004991(.in0(tmp00_76_39), .in1(tmp00_77_39), .out(tmp01_38_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004992(.in0(tmp00_78_39), .in1(tmp00_79_39), .out(tmp01_39_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004993(.in0(tmp00_80_39), .in1(tmp00_81_39), .out(tmp01_40_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004994(.in0(tmp00_82_39), .in1(tmp00_83_39), .out(tmp01_41_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004995(.in0(tmp00_84_39), .in1(tmp00_85_39), .out(tmp01_42_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004996(.in0(tmp00_86_39), .in1(tmp00_87_39), .out(tmp01_43_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004997(.in0(tmp00_88_39), .in1(tmp00_89_39), .out(tmp01_44_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004998(.in0(tmp00_90_39), .in1(tmp00_91_39), .out(tmp01_45_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add004999(.in0(tmp00_92_39), .in1(tmp00_93_39), .out(tmp01_46_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005000(.in0(tmp00_94_39), .in1(tmp00_95_39), .out(tmp01_47_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005001(.in0(tmp00_96_39), .in1(tmp00_97_39), .out(tmp01_48_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005002(.in0(tmp00_98_39), .in1(tmp00_99_39), .out(tmp01_49_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005003(.in0(tmp00_100_39), .in1(tmp00_101_39), .out(tmp01_50_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005004(.in0(tmp00_102_39), .in1(tmp00_103_39), .out(tmp01_51_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005005(.in0(tmp00_104_39), .in1(tmp00_105_39), .out(tmp01_52_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005006(.in0(tmp00_106_39), .in1(tmp00_107_39), .out(tmp01_53_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005007(.in0(tmp00_108_39), .in1(tmp00_109_39), .out(tmp01_54_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005008(.in0(tmp00_110_39), .in1(tmp00_111_39), .out(tmp01_55_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005009(.in0(tmp00_112_39), .in1(tmp00_113_39), .out(tmp01_56_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005010(.in0(tmp00_114_39), .in1(tmp00_115_39), .out(tmp01_57_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005011(.in0(tmp00_116_39), .in1(tmp00_117_39), .out(tmp01_58_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005012(.in0(tmp00_118_39), .in1(tmp00_119_39), .out(tmp01_59_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005013(.in0(tmp00_120_39), .in1(tmp00_121_39), .out(tmp01_60_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005014(.in0(tmp00_122_39), .in1(tmp00_123_39), .out(tmp01_61_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005015(.in0(tmp00_124_39), .in1(tmp00_125_39), .out(tmp01_62_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005016(.in0(tmp00_126_39), .in1(tmp00_127_39), .out(tmp01_63_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005017(.in0(tmp01_0_39), .in1(tmp01_1_39), .out(tmp02_0_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005018(.in0(tmp01_2_39), .in1(tmp01_3_39), .out(tmp02_1_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005019(.in0(tmp01_4_39), .in1(tmp01_5_39), .out(tmp02_2_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005020(.in0(tmp01_6_39), .in1(tmp01_7_39), .out(tmp02_3_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005021(.in0(tmp01_8_39), .in1(tmp01_9_39), .out(tmp02_4_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005022(.in0(tmp01_10_39), .in1(tmp01_11_39), .out(tmp02_5_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005023(.in0(tmp01_12_39), .in1(tmp01_13_39), .out(tmp02_6_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005024(.in0(tmp01_14_39), .in1(tmp01_15_39), .out(tmp02_7_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005025(.in0(tmp01_16_39), .in1(tmp01_17_39), .out(tmp02_8_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005026(.in0(tmp01_18_39), .in1(tmp01_19_39), .out(tmp02_9_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005027(.in0(tmp01_20_39), .in1(tmp01_21_39), .out(tmp02_10_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005028(.in0(tmp01_22_39), .in1(tmp01_23_39), .out(tmp02_11_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005029(.in0(tmp01_24_39), .in1(tmp01_25_39), .out(tmp02_12_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005030(.in0(tmp01_26_39), .in1(tmp01_27_39), .out(tmp02_13_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005031(.in0(tmp01_28_39), .in1(tmp01_29_39), .out(tmp02_14_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005032(.in0(tmp01_30_39), .in1(tmp01_31_39), .out(tmp02_15_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005033(.in0(tmp01_32_39), .in1(tmp01_33_39), .out(tmp02_16_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005034(.in0(tmp01_34_39), .in1(tmp01_35_39), .out(tmp02_17_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005035(.in0(tmp01_36_39), .in1(tmp01_37_39), .out(tmp02_18_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005036(.in0(tmp01_38_39), .in1(tmp01_39_39), .out(tmp02_19_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005037(.in0(tmp01_40_39), .in1(tmp01_41_39), .out(tmp02_20_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005038(.in0(tmp01_42_39), .in1(tmp01_43_39), .out(tmp02_21_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005039(.in0(tmp01_44_39), .in1(tmp01_45_39), .out(tmp02_22_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005040(.in0(tmp01_46_39), .in1(tmp01_47_39), .out(tmp02_23_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005041(.in0(tmp01_48_39), .in1(tmp01_49_39), .out(tmp02_24_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005042(.in0(tmp01_50_39), .in1(tmp01_51_39), .out(tmp02_25_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005043(.in0(tmp01_52_39), .in1(tmp01_53_39), .out(tmp02_26_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005044(.in0(tmp01_54_39), .in1(tmp01_55_39), .out(tmp02_27_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005045(.in0(tmp01_56_39), .in1(tmp01_57_39), .out(tmp02_28_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005046(.in0(tmp01_58_39), .in1(tmp01_59_39), .out(tmp02_29_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005047(.in0(tmp01_60_39), .in1(tmp01_61_39), .out(tmp02_30_39));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005048(.in0(tmp01_62_39), .in1(tmp01_63_39), .out(tmp02_31_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005049(.in0(tmp02_0_39), .in1(tmp02_1_39), .out(tmp03_0_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005050(.in0(tmp02_2_39), .in1(tmp02_3_39), .out(tmp03_1_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005051(.in0(tmp02_4_39), .in1(tmp02_5_39), .out(tmp03_2_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005052(.in0(tmp02_6_39), .in1(tmp02_7_39), .out(tmp03_3_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005053(.in0(tmp02_8_39), .in1(tmp02_9_39), .out(tmp03_4_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005054(.in0(tmp02_10_39), .in1(tmp02_11_39), .out(tmp03_5_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005055(.in0(tmp02_12_39), .in1(tmp02_13_39), .out(tmp03_6_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005056(.in0(tmp02_14_39), .in1(tmp02_15_39), .out(tmp03_7_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005057(.in0(tmp02_16_39), .in1(tmp02_17_39), .out(tmp03_8_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005058(.in0(tmp02_18_39), .in1(tmp02_19_39), .out(tmp03_9_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005059(.in0(tmp02_20_39), .in1(tmp02_21_39), .out(tmp03_10_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005060(.in0(tmp02_22_39), .in1(tmp02_23_39), .out(tmp03_11_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005061(.in0(tmp02_24_39), .in1(tmp02_25_39), .out(tmp03_12_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005062(.in0(tmp02_26_39), .in1(tmp02_27_39), .out(tmp03_13_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005063(.in0(tmp02_28_39), .in1(tmp02_29_39), .out(tmp03_14_39));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005064(.in0(tmp02_30_39), .in1(tmp02_31_39), .out(tmp03_15_39));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005065(.in0(tmp03_0_39), .in1(tmp03_1_39), .out(tmp04_0_39));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005066(.in0(tmp03_2_39), .in1(tmp03_3_39), .out(tmp04_1_39));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005067(.in0(tmp03_4_39), .in1(tmp03_5_39), .out(tmp04_2_39));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005068(.in0(tmp03_6_39), .in1(tmp03_7_39), .out(tmp04_3_39));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005069(.in0(tmp03_8_39), .in1(tmp03_9_39), .out(tmp04_4_39));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005070(.in0(tmp03_10_39), .in1(tmp03_11_39), .out(tmp04_5_39));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005071(.in0(tmp03_12_39), .in1(tmp03_13_39), .out(tmp04_6_39));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005072(.in0(tmp03_14_39), .in1(tmp03_15_39), .out(tmp04_7_39));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005073(.in0(tmp04_0_39), .in1(tmp04_1_39), .out(tmp05_0_39));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005074(.in0(tmp04_2_39), .in1(tmp04_3_39), .out(tmp05_1_39));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005075(.in0(tmp04_4_39), .in1(tmp04_5_39), .out(tmp05_2_39));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005076(.in0(tmp04_6_39), .in1(tmp04_7_39), .out(tmp05_3_39));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005077(.in0(tmp05_0_39), .in1(tmp05_1_39), .out(tmp06_0_39));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005078(.in0(tmp05_2_39), .in1(tmp05_3_39), .out(tmp06_1_39));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add005079(.in0(tmp06_0_39), .in1(tmp06_1_39), .out(tmp07_0_39));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005080(.in0(tmp00_0_40), .in1(tmp00_1_40), .out(tmp01_0_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005081(.in0(tmp00_2_40), .in1(tmp00_3_40), .out(tmp01_1_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005082(.in0(tmp00_4_40), .in1(tmp00_5_40), .out(tmp01_2_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005083(.in0(tmp00_6_40), .in1(tmp00_7_40), .out(tmp01_3_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005084(.in0(tmp00_8_40), .in1(tmp00_9_40), .out(tmp01_4_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005085(.in0(tmp00_10_40), .in1(tmp00_11_40), .out(tmp01_5_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005086(.in0(tmp00_12_40), .in1(tmp00_13_40), .out(tmp01_6_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005087(.in0(tmp00_14_40), .in1(tmp00_15_40), .out(tmp01_7_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005088(.in0(tmp00_16_40), .in1(tmp00_17_40), .out(tmp01_8_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005089(.in0(tmp00_18_40), .in1(tmp00_19_40), .out(tmp01_9_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005090(.in0(tmp00_20_40), .in1(tmp00_21_40), .out(tmp01_10_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005091(.in0(tmp00_22_40), .in1(tmp00_23_40), .out(tmp01_11_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005092(.in0(tmp00_24_40), .in1(tmp00_25_40), .out(tmp01_12_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005093(.in0(tmp00_26_40), .in1(tmp00_27_40), .out(tmp01_13_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005094(.in0(tmp00_28_40), .in1(tmp00_29_40), .out(tmp01_14_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005095(.in0(tmp00_30_40), .in1(tmp00_31_40), .out(tmp01_15_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005096(.in0(tmp00_32_40), .in1(tmp00_33_40), .out(tmp01_16_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005097(.in0(tmp00_34_40), .in1(tmp00_35_40), .out(tmp01_17_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005098(.in0(tmp00_36_40), .in1(tmp00_37_40), .out(tmp01_18_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005099(.in0(tmp00_38_40), .in1(tmp00_39_40), .out(tmp01_19_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005100(.in0(tmp00_40_40), .in1(tmp00_41_40), .out(tmp01_20_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005101(.in0(tmp00_42_40), .in1(tmp00_43_40), .out(tmp01_21_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005102(.in0(tmp00_44_40), .in1(tmp00_45_40), .out(tmp01_22_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005103(.in0(tmp00_46_40), .in1(tmp00_47_40), .out(tmp01_23_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005104(.in0(tmp00_48_40), .in1(tmp00_49_40), .out(tmp01_24_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005105(.in0(tmp00_50_40), .in1(tmp00_51_40), .out(tmp01_25_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005106(.in0(tmp00_52_40), .in1(tmp00_53_40), .out(tmp01_26_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005107(.in0(tmp00_54_40), .in1(tmp00_55_40), .out(tmp01_27_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005108(.in0(tmp00_56_40), .in1(tmp00_57_40), .out(tmp01_28_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005109(.in0(tmp00_58_40), .in1(tmp00_59_40), .out(tmp01_29_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005110(.in0(tmp00_60_40), .in1(tmp00_61_40), .out(tmp01_30_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005111(.in0(tmp00_62_40), .in1(tmp00_63_40), .out(tmp01_31_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005112(.in0(tmp00_64_40), .in1(tmp00_65_40), .out(tmp01_32_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005113(.in0(tmp00_66_40), .in1(tmp00_67_40), .out(tmp01_33_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005114(.in0(tmp00_68_40), .in1(tmp00_69_40), .out(tmp01_34_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005115(.in0(tmp00_70_40), .in1(tmp00_71_40), .out(tmp01_35_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005116(.in0(tmp00_72_40), .in1(tmp00_73_40), .out(tmp01_36_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005117(.in0(tmp00_74_40), .in1(tmp00_75_40), .out(tmp01_37_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005118(.in0(tmp00_76_40), .in1(tmp00_77_40), .out(tmp01_38_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005119(.in0(tmp00_78_40), .in1(tmp00_79_40), .out(tmp01_39_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005120(.in0(tmp00_80_40), .in1(tmp00_81_40), .out(tmp01_40_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005121(.in0(tmp00_82_40), .in1(tmp00_83_40), .out(tmp01_41_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005122(.in0(tmp00_84_40), .in1(tmp00_85_40), .out(tmp01_42_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005123(.in0(tmp00_86_40), .in1(tmp00_87_40), .out(tmp01_43_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005124(.in0(tmp00_88_40), .in1(tmp00_89_40), .out(tmp01_44_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005125(.in0(tmp00_90_40), .in1(tmp00_91_40), .out(tmp01_45_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005126(.in0(tmp00_92_40), .in1(tmp00_93_40), .out(tmp01_46_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005127(.in0(tmp00_94_40), .in1(tmp00_95_40), .out(tmp01_47_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005128(.in0(tmp00_96_40), .in1(tmp00_97_40), .out(tmp01_48_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005129(.in0(tmp00_98_40), .in1(tmp00_99_40), .out(tmp01_49_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005130(.in0(tmp00_100_40), .in1(tmp00_101_40), .out(tmp01_50_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005131(.in0(tmp00_102_40), .in1(tmp00_103_40), .out(tmp01_51_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005132(.in0(tmp00_104_40), .in1(tmp00_105_40), .out(tmp01_52_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005133(.in0(tmp00_106_40), .in1(tmp00_107_40), .out(tmp01_53_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005134(.in0(tmp00_108_40), .in1(tmp00_109_40), .out(tmp01_54_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005135(.in0(tmp00_110_40), .in1(tmp00_111_40), .out(tmp01_55_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005136(.in0(tmp00_112_40), .in1(tmp00_113_40), .out(tmp01_56_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005137(.in0(tmp00_114_40), .in1(tmp00_115_40), .out(tmp01_57_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005138(.in0(tmp00_116_40), .in1(tmp00_117_40), .out(tmp01_58_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005139(.in0(tmp00_118_40), .in1(tmp00_119_40), .out(tmp01_59_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005140(.in0(tmp00_120_40), .in1(tmp00_121_40), .out(tmp01_60_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005141(.in0(tmp00_122_40), .in1(tmp00_123_40), .out(tmp01_61_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005142(.in0(tmp00_124_40), .in1(tmp00_125_40), .out(tmp01_62_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005143(.in0(tmp00_126_40), .in1(tmp00_127_40), .out(tmp01_63_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005144(.in0(tmp01_0_40), .in1(tmp01_1_40), .out(tmp02_0_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005145(.in0(tmp01_2_40), .in1(tmp01_3_40), .out(tmp02_1_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005146(.in0(tmp01_4_40), .in1(tmp01_5_40), .out(tmp02_2_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005147(.in0(tmp01_6_40), .in1(tmp01_7_40), .out(tmp02_3_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005148(.in0(tmp01_8_40), .in1(tmp01_9_40), .out(tmp02_4_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005149(.in0(tmp01_10_40), .in1(tmp01_11_40), .out(tmp02_5_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005150(.in0(tmp01_12_40), .in1(tmp01_13_40), .out(tmp02_6_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005151(.in0(tmp01_14_40), .in1(tmp01_15_40), .out(tmp02_7_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005152(.in0(tmp01_16_40), .in1(tmp01_17_40), .out(tmp02_8_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005153(.in0(tmp01_18_40), .in1(tmp01_19_40), .out(tmp02_9_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005154(.in0(tmp01_20_40), .in1(tmp01_21_40), .out(tmp02_10_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005155(.in0(tmp01_22_40), .in1(tmp01_23_40), .out(tmp02_11_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005156(.in0(tmp01_24_40), .in1(tmp01_25_40), .out(tmp02_12_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005157(.in0(tmp01_26_40), .in1(tmp01_27_40), .out(tmp02_13_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005158(.in0(tmp01_28_40), .in1(tmp01_29_40), .out(tmp02_14_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005159(.in0(tmp01_30_40), .in1(tmp01_31_40), .out(tmp02_15_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005160(.in0(tmp01_32_40), .in1(tmp01_33_40), .out(tmp02_16_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005161(.in0(tmp01_34_40), .in1(tmp01_35_40), .out(tmp02_17_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005162(.in0(tmp01_36_40), .in1(tmp01_37_40), .out(tmp02_18_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005163(.in0(tmp01_38_40), .in1(tmp01_39_40), .out(tmp02_19_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005164(.in0(tmp01_40_40), .in1(tmp01_41_40), .out(tmp02_20_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005165(.in0(tmp01_42_40), .in1(tmp01_43_40), .out(tmp02_21_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005166(.in0(tmp01_44_40), .in1(tmp01_45_40), .out(tmp02_22_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005167(.in0(tmp01_46_40), .in1(tmp01_47_40), .out(tmp02_23_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005168(.in0(tmp01_48_40), .in1(tmp01_49_40), .out(tmp02_24_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005169(.in0(tmp01_50_40), .in1(tmp01_51_40), .out(tmp02_25_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005170(.in0(tmp01_52_40), .in1(tmp01_53_40), .out(tmp02_26_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005171(.in0(tmp01_54_40), .in1(tmp01_55_40), .out(tmp02_27_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005172(.in0(tmp01_56_40), .in1(tmp01_57_40), .out(tmp02_28_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005173(.in0(tmp01_58_40), .in1(tmp01_59_40), .out(tmp02_29_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005174(.in0(tmp01_60_40), .in1(tmp01_61_40), .out(tmp02_30_40));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005175(.in0(tmp01_62_40), .in1(tmp01_63_40), .out(tmp02_31_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005176(.in0(tmp02_0_40), .in1(tmp02_1_40), .out(tmp03_0_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005177(.in0(tmp02_2_40), .in1(tmp02_3_40), .out(tmp03_1_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005178(.in0(tmp02_4_40), .in1(tmp02_5_40), .out(tmp03_2_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005179(.in0(tmp02_6_40), .in1(tmp02_7_40), .out(tmp03_3_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005180(.in0(tmp02_8_40), .in1(tmp02_9_40), .out(tmp03_4_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005181(.in0(tmp02_10_40), .in1(tmp02_11_40), .out(tmp03_5_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005182(.in0(tmp02_12_40), .in1(tmp02_13_40), .out(tmp03_6_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005183(.in0(tmp02_14_40), .in1(tmp02_15_40), .out(tmp03_7_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005184(.in0(tmp02_16_40), .in1(tmp02_17_40), .out(tmp03_8_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005185(.in0(tmp02_18_40), .in1(tmp02_19_40), .out(tmp03_9_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005186(.in0(tmp02_20_40), .in1(tmp02_21_40), .out(tmp03_10_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005187(.in0(tmp02_22_40), .in1(tmp02_23_40), .out(tmp03_11_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005188(.in0(tmp02_24_40), .in1(tmp02_25_40), .out(tmp03_12_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005189(.in0(tmp02_26_40), .in1(tmp02_27_40), .out(tmp03_13_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005190(.in0(tmp02_28_40), .in1(tmp02_29_40), .out(tmp03_14_40));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005191(.in0(tmp02_30_40), .in1(tmp02_31_40), .out(tmp03_15_40));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005192(.in0(tmp03_0_40), .in1(tmp03_1_40), .out(tmp04_0_40));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005193(.in0(tmp03_2_40), .in1(tmp03_3_40), .out(tmp04_1_40));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005194(.in0(tmp03_4_40), .in1(tmp03_5_40), .out(tmp04_2_40));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005195(.in0(tmp03_6_40), .in1(tmp03_7_40), .out(tmp04_3_40));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005196(.in0(tmp03_8_40), .in1(tmp03_9_40), .out(tmp04_4_40));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005197(.in0(tmp03_10_40), .in1(tmp03_11_40), .out(tmp04_5_40));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005198(.in0(tmp03_12_40), .in1(tmp03_13_40), .out(tmp04_6_40));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005199(.in0(tmp03_14_40), .in1(tmp03_15_40), .out(tmp04_7_40));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005200(.in0(tmp04_0_40), .in1(tmp04_1_40), .out(tmp05_0_40));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005201(.in0(tmp04_2_40), .in1(tmp04_3_40), .out(tmp05_1_40));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005202(.in0(tmp04_4_40), .in1(tmp04_5_40), .out(tmp05_2_40));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005203(.in0(tmp04_6_40), .in1(tmp04_7_40), .out(tmp05_3_40));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005204(.in0(tmp05_0_40), .in1(tmp05_1_40), .out(tmp06_0_40));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005205(.in0(tmp05_2_40), .in1(tmp05_3_40), .out(tmp06_1_40));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add005206(.in0(tmp06_0_40), .in1(tmp06_1_40), .out(tmp07_0_40));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005207(.in0(tmp00_0_41), .in1(tmp00_1_41), .out(tmp01_0_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005208(.in0(tmp00_2_41), .in1(tmp00_3_41), .out(tmp01_1_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005209(.in0(tmp00_4_41), .in1(tmp00_5_41), .out(tmp01_2_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005210(.in0(tmp00_6_41), .in1(tmp00_7_41), .out(tmp01_3_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005211(.in0(tmp00_8_41), .in1(tmp00_9_41), .out(tmp01_4_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005212(.in0(tmp00_10_41), .in1(tmp00_11_41), .out(tmp01_5_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005213(.in0(tmp00_12_41), .in1(tmp00_13_41), .out(tmp01_6_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005214(.in0(tmp00_14_41), .in1(tmp00_15_41), .out(tmp01_7_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005215(.in0(tmp00_16_41), .in1(tmp00_17_41), .out(tmp01_8_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005216(.in0(tmp00_18_41), .in1(tmp00_19_41), .out(tmp01_9_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005217(.in0(tmp00_20_41), .in1(tmp00_21_41), .out(tmp01_10_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005218(.in0(tmp00_22_41), .in1(tmp00_23_41), .out(tmp01_11_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005219(.in0(tmp00_24_41), .in1(tmp00_25_41), .out(tmp01_12_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005220(.in0(tmp00_26_41), .in1(tmp00_27_41), .out(tmp01_13_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005221(.in0(tmp00_28_41), .in1(tmp00_29_41), .out(tmp01_14_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005222(.in0(tmp00_30_41), .in1(tmp00_31_41), .out(tmp01_15_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005223(.in0(tmp00_32_41), .in1(tmp00_33_41), .out(tmp01_16_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005224(.in0(tmp00_34_41), .in1(tmp00_35_41), .out(tmp01_17_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005225(.in0(tmp00_36_41), .in1(tmp00_37_41), .out(tmp01_18_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005226(.in0(tmp00_38_41), .in1(tmp00_39_41), .out(tmp01_19_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005227(.in0(tmp00_40_41), .in1(tmp00_41_41), .out(tmp01_20_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005228(.in0(tmp00_42_41), .in1(tmp00_43_41), .out(tmp01_21_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005229(.in0(tmp00_44_41), .in1(tmp00_45_41), .out(tmp01_22_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005230(.in0(tmp00_46_41), .in1(tmp00_47_41), .out(tmp01_23_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005231(.in0(tmp00_48_41), .in1(tmp00_49_41), .out(tmp01_24_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005232(.in0(tmp00_50_41), .in1(tmp00_51_41), .out(tmp01_25_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005233(.in0(tmp00_52_41), .in1(tmp00_53_41), .out(tmp01_26_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005234(.in0(tmp00_54_41), .in1(tmp00_55_41), .out(tmp01_27_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005235(.in0(tmp00_56_41), .in1(tmp00_57_41), .out(tmp01_28_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005236(.in0(tmp00_58_41), .in1(tmp00_59_41), .out(tmp01_29_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005237(.in0(tmp00_60_41), .in1(tmp00_61_41), .out(tmp01_30_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005238(.in0(tmp00_62_41), .in1(tmp00_63_41), .out(tmp01_31_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005239(.in0(tmp00_64_41), .in1(tmp00_65_41), .out(tmp01_32_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005240(.in0(tmp00_66_41), .in1(tmp00_67_41), .out(tmp01_33_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005241(.in0(tmp00_68_41), .in1(tmp00_69_41), .out(tmp01_34_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005242(.in0(tmp00_70_41), .in1(tmp00_71_41), .out(tmp01_35_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005243(.in0(tmp00_72_41), .in1(tmp00_73_41), .out(tmp01_36_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005244(.in0(tmp00_74_41), .in1(tmp00_75_41), .out(tmp01_37_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005245(.in0(tmp00_76_41), .in1(tmp00_77_41), .out(tmp01_38_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005246(.in0(tmp00_78_41), .in1(tmp00_79_41), .out(tmp01_39_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005247(.in0(tmp00_80_41), .in1(tmp00_81_41), .out(tmp01_40_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005248(.in0(tmp00_82_41), .in1(tmp00_83_41), .out(tmp01_41_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005249(.in0(tmp00_84_41), .in1(tmp00_85_41), .out(tmp01_42_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005250(.in0(tmp00_86_41), .in1(tmp00_87_41), .out(tmp01_43_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005251(.in0(tmp00_88_41), .in1(tmp00_89_41), .out(tmp01_44_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005252(.in0(tmp00_90_41), .in1(tmp00_91_41), .out(tmp01_45_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005253(.in0(tmp00_92_41), .in1(tmp00_93_41), .out(tmp01_46_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005254(.in0(tmp00_94_41), .in1(tmp00_95_41), .out(tmp01_47_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005255(.in0(tmp00_96_41), .in1(tmp00_97_41), .out(tmp01_48_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005256(.in0(tmp00_98_41), .in1(tmp00_99_41), .out(tmp01_49_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005257(.in0(tmp00_100_41), .in1(tmp00_101_41), .out(tmp01_50_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005258(.in0(tmp00_102_41), .in1(tmp00_103_41), .out(tmp01_51_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005259(.in0(tmp00_104_41), .in1(tmp00_105_41), .out(tmp01_52_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005260(.in0(tmp00_106_41), .in1(tmp00_107_41), .out(tmp01_53_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005261(.in0(tmp00_108_41), .in1(tmp00_109_41), .out(tmp01_54_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005262(.in0(tmp00_110_41), .in1(tmp00_111_41), .out(tmp01_55_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005263(.in0(tmp00_112_41), .in1(tmp00_113_41), .out(tmp01_56_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005264(.in0(tmp00_114_41), .in1(tmp00_115_41), .out(tmp01_57_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005265(.in0(tmp00_116_41), .in1(tmp00_117_41), .out(tmp01_58_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005266(.in0(tmp00_118_41), .in1(tmp00_119_41), .out(tmp01_59_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005267(.in0(tmp00_120_41), .in1(tmp00_121_41), .out(tmp01_60_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005268(.in0(tmp00_122_41), .in1(tmp00_123_41), .out(tmp01_61_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005269(.in0(tmp00_124_41), .in1(tmp00_125_41), .out(tmp01_62_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005270(.in0(tmp00_126_41), .in1(tmp00_127_41), .out(tmp01_63_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005271(.in0(tmp01_0_41), .in1(tmp01_1_41), .out(tmp02_0_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005272(.in0(tmp01_2_41), .in1(tmp01_3_41), .out(tmp02_1_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005273(.in0(tmp01_4_41), .in1(tmp01_5_41), .out(tmp02_2_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005274(.in0(tmp01_6_41), .in1(tmp01_7_41), .out(tmp02_3_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005275(.in0(tmp01_8_41), .in1(tmp01_9_41), .out(tmp02_4_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005276(.in0(tmp01_10_41), .in1(tmp01_11_41), .out(tmp02_5_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005277(.in0(tmp01_12_41), .in1(tmp01_13_41), .out(tmp02_6_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005278(.in0(tmp01_14_41), .in1(tmp01_15_41), .out(tmp02_7_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005279(.in0(tmp01_16_41), .in1(tmp01_17_41), .out(tmp02_8_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005280(.in0(tmp01_18_41), .in1(tmp01_19_41), .out(tmp02_9_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005281(.in0(tmp01_20_41), .in1(tmp01_21_41), .out(tmp02_10_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005282(.in0(tmp01_22_41), .in1(tmp01_23_41), .out(tmp02_11_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005283(.in0(tmp01_24_41), .in1(tmp01_25_41), .out(tmp02_12_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005284(.in0(tmp01_26_41), .in1(tmp01_27_41), .out(tmp02_13_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005285(.in0(tmp01_28_41), .in1(tmp01_29_41), .out(tmp02_14_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005286(.in0(tmp01_30_41), .in1(tmp01_31_41), .out(tmp02_15_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005287(.in0(tmp01_32_41), .in1(tmp01_33_41), .out(tmp02_16_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005288(.in0(tmp01_34_41), .in1(tmp01_35_41), .out(tmp02_17_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005289(.in0(tmp01_36_41), .in1(tmp01_37_41), .out(tmp02_18_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005290(.in0(tmp01_38_41), .in1(tmp01_39_41), .out(tmp02_19_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005291(.in0(tmp01_40_41), .in1(tmp01_41_41), .out(tmp02_20_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005292(.in0(tmp01_42_41), .in1(tmp01_43_41), .out(tmp02_21_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005293(.in0(tmp01_44_41), .in1(tmp01_45_41), .out(tmp02_22_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005294(.in0(tmp01_46_41), .in1(tmp01_47_41), .out(tmp02_23_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005295(.in0(tmp01_48_41), .in1(tmp01_49_41), .out(tmp02_24_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005296(.in0(tmp01_50_41), .in1(tmp01_51_41), .out(tmp02_25_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005297(.in0(tmp01_52_41), .in1(tmp01_53_41), .out(tmp02_26_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005298(.in0(tmp01_54_41), .in1(tmp01_55_41), .out(tmp02_27_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005299(.in0(tmp01_56_41), .in1(tmp01_57_41), .out(tmp02_28_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005300(.in0(tmp01_58_41), .in1(tmp01_59_41), .out(tmp02_29_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005301(.in0(tmp01_60_41), .in1(tmp01_61_41), .out(tmp02_30_41));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005302(.in0(tmp01_62_41), .in1(tmp01_63_41), .out(tmp02_31_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005303(.in0(tmp02_0_41), .in1(tmp02_1_41), .out(tmp03_0_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005304(.in0(tmp02_2_41), .in1(tmp02_3_41), .out(tmp03_1_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005305(.in0(tmp02_4_41), .in1(tmp02_5_41), .out(tmp03_2_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005306(.in0(tmp02_6_41), .in1(tmp02_7_41), .out(tmp03_3_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005307(.in0(tmp02_8_41), .in1(tmp02_9_41), .out(tmp03_4_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005308(.in0(tmp02_10_41), .in1(tmp02_11_41), .out(tmp03_5_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005309(.in0(tmp02_12_41), .in1(tmp02_13_41), .out(tmp03_6_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005310(.in0(tmp02_14_41), .in1(tmp02_15_41), .out(tmp03_7_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005311(.in0(tmp02_16_41), .in1(tmp02_17_41), .out(tmp03_8_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005312(.in0(tmp02_18_41), .in1(tmp02_19_41), .out(tmp03_9_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005313(.in0(tmp02_20_41), .in1(tmp02_21_41), .out(tmp03_10_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005314(.in0(tmp02_22_41), .in1(tmp02_23_41), .out(tmp03_11_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005315(.in0(tmp02_24_41), .in1(tmp02_25_41), .out(tmp03_12_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005316(.in0(tmp02_26_41), .in1(tmp02_27_41), .out(tmp03_13_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005317(.in0(tmp02_28_41), .in1(tmp02_29_41), .out(tmp03_14_41));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005318(.in0(tmp02_30_41), .in1(tmp02_31_41), .out(tmp03_15_41));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005319(.in0(tmp03_0_41), .in1(tmp03_1_41), .out(tmp04_0_41));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005320(.in0(tmp03_2_41), .in1(tmp03_3_41), .out(tmp04_1_41));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005321(.in0(tmp03_4_41), .in1(tmp03_5_41), .out(tmp04_2_41));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005322(.in0(tmp03_6_41), .in1(tmp03_7_41), .out(tmp04_3_41));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005323(.in0(tmp03_8_41), .in1(tmp03_9_41), .out(tmp04_4_41));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005324(.in0(tmp03_10_41), .in1(tmp03_11_41), .out(tmp04_5_41));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005325(.in0(tmp03_12_41), .in1(tmp03_13_41), .out(tmp04_6_41));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005326(.in0(tmp03_14_41), .in1(tmp03_15_41), .out(tmp04_7_41));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005327(.in0(tmp04_0_41), .in1(tmp04_1_41), .out(tmp05_0_41));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005328(.in0(tmp04_2_41), .in1(tmp04_3_41), .out(tmp05_1_41));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005329(.in0(tmp04_4_41), .in1(tmp04_5_41), .out(tmp05_2_41));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005330(.in0(tmp04_6_41), .in1(tmp04_7_41), .out(tmp05_3_41));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005331(.in0(tmp05_0_41), .in1(tmp05_1_41), .out(tmp06_0_41));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005332(.in0(tmp05_2_41), .in1(tmp05_3_41), .out(tmp06_1_41));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add005333(.in0(tmp06_0_41), .in1(tmp06_1_41), .out(tmp07_0_41));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005334(.in0(tmp00_0_42), .in1(tmp00_1_42), .out(tmp01_0_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005335(.in0(tmp00_2_42), .in1(tmp00_3_42), .out(tmp01_1_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005336(.in0(tmp00_4_42), .in1(tmp00_5_42), .out(tmp01_2_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005337(.in0(tmp00_6_42), .in1(tmp00_7_42), .out(tmp01_3_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005338(.in0(tmp00_8_42), .in1(tmp00_9_42), .out(tmp01_4_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005339(.in0(tmp00_10_42), .in1(tmp00_11_42), .out(tmp01_5_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005340(.in0(tmp00_12_42), .in1(tmp00_13_42), .out(tmp01_6_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005341(.in0(tmp00_14_42), .in1(tmp00_15_42), .out(tmp01_7_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005342(.in0(tmp00_16_42), .in1(tmp00_17_42), .out(tmp01_8_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005343(.in0(tmp00_18_42), .in1(tmp00_19_42), .out(tmp01_9_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005344(.in0(tmp00_20_42), .in1(tmp00_21_42), .out(tmp01_10_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005345(.in0(tmp00_22_42), .in1(tmp00_23_42), .out(tmp01_11_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005346(.in0(tmp00_24_42), .in1(tmp00_25_42), .out(tmp01_12_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005347(.in0(tmp00_26_42), .in1(tmp00_27_42), .out(tmp01_13_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005348(.in0(tmp00_28_42), .in1(tmp00_29_42), .out(tmp01_14_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005349(.in0(tmp00_30_42), .in1(tmp00_31_42), .out(tmp01_15_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005350(.in0(tmp00_32_42), .in1(tmp00_33_42), .out(tmp01_16_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005351(.in0(tmp00_34_42), .in1(tmp00_35_42), .out(tmp01_17_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005352(.in0(tmp00_36_42), .in1(tmp00_37_42), .out(tmp01_18_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005353(.in0(tmp00_38_42), .in1(tmp00_39_42), .out(tmp01_19_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005354(.in0(tmp00_40_42), .in1(tmp00_41_42), .out(tmp01_20_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005355(.in0(tmp00_42_42), .in1(tmp00_43_42), .out(tmp01_21_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005356(.in0(tmp00_44_42), .in1(tmp00_45_42), .out(tmp01_22_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005357(.in0(tmp00_46_42), .in1(tmp00_47_42), .out(tmp01_23_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005358(.in0(tmp00_48_42), .in1(tmp00_49_42), .out(tmp01_24_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005359(.in0(tmp00_50_42), .in1(tmp00_51_42), .out(tmp01_25_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005360(.in0(tmp00_52_42), .in1(tmp00_53_42), .out(tmp01_26_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005361(.in0(tmp00_54_42), .in1(tmp00_55_42), .out(tmp01_27_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005362(.in0(tmp00_56_42), .in1(tmp00_57_42), .out(tmp01_28_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005363(.in0(tmp00_58_42), .in1(tmp00_59_42), .out(tmp01_29_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005364(.in0(tmp00_60_42), .in1(tmp00_61_42), .out(tmp01_30_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005365(.in0(tmp00_62_42), .in1(tmp00_63_42), .out(tmp01_31_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005366(.in0(tmp00_64_42), .in1(tmp00_65_42), .out(tmp01_32_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005367(.in0(tmp00_66_42), .in1(tmp00_67_42), .out(tmp01_33_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005368(.in0(tmp00_68_42), .in1(tmp00_69_42), .out(tmp01_34_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005369(.in0(tmp00_70_42), .in1(tmp00_71_42), .out(tmp01_35_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005370(.in0(tmp00_72_42), .in1(tmp00_73_42), .out(tmp01_36_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005371(.in0(tmp00_74_42), .in1(tmp00_75_42), .out(tmp01_37_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005372(.in0(tmp00_76_42), .in1(tmp00_77_42), .out(tmp01_38_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005373(.in0(tmp00_78_42), .in1(tmp00_79_42), .out(tmp01_39_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005374(.in0(tmp00_80_42), .in1(tmp00_81_42), .out(tmp01_40_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005375(.in0(tmp00_82_42), .in1(tmp00_83_42), .out(tmp01_41_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005376(.in0(tmp00_84_42), .in1(tmp00_85_42), .out(tmp01_42_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005377(.in0(tmp00_86_42), .in1(tmp00_87_42), .out(tmp01_43_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005378(.in0(tmp00_88_42), .in1(tmp00_89_42), .out(tmp01_44_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005379(.in0(tmp00_90_42), .in1(tmp00_91_42), .out(tmp01_45_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005380(.in0(tmp00_92_42), .in1(tmp00_93_42), .out(tmp01_46_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005381(.in0(tmp00_94_42), .in1(tmp00_95_42), .out(tmp01_47_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005382(.in0(tmp00_96_42), .in1(tmp00_97_42), .out(tmp01_48_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005383(.in0(tmp00_98_42), .in1(tmp00_99_42), .out(tmp01_49_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005384(.in0(tmp00_100_42), .in1(tmp00_101_42), .out(tmp01_50_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005385(.in0(tmp00_102_42), .in1(tmp00_103_42), .out(tmp01_51_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005386(.in0(tmp00_104_42), .in1(tmp00_105_42), .out(tmp01_52_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005387(.in0(tmp00_106_42), .in1(tmp00_107_42), .out(tmp01_53_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005388(.in0(tmp00_108_42), .in1(tmp00_109_42), .out(tmp01_54_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005389(.in0(tmp00_110_42), .in1(tmp00_111_42), .out(tmp01_55_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005390(.in0(tmp00_112_42), .in1(tmp00_113_42), .out(tmp01_56_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005391(.in0(tmp00_114_42), .in1(tmp00_115_42), .out(tmp01_57_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005392(.in0(tmp00_116_42), .in1(tmp00_117_42), .out(tmp01_58_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005393(.in0(tmp00_118_42), .in1(tmp00_119_42), .out(tmp01_59_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005394(.in0(tmp00_120_42), .in1(tmp00_121_42), .out(tmp01_60_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005395(.in0(tmp00_122_42), .in1(tmp00_123_42), .out(tmp01_61_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005396(.in0(tmp00_124_42), .in1(tmp00_125_42), .out(tmp01_62_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005397(.in0(tmp00_126_42), .in1(tmp00_127_42), .out(tmp01_63_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005398(.in0(tmp01_0_42), .in1(tmp01_1_42), .out(tmp02_0_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005399(.in0(tmp01_2_42), .in1(tmp01_3_42), .out(tmp02_1_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005400(.in0(tmp01_4_42), .in1(tmp01_5_42), .out(tmp02_2_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005401(.in0(tmp01_6_42), .in1(tmp01_7_42), .out(tmp02_3_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005402(.in0(tmp01_8_42), .in1(tmp01_9_42), .out(tmp02_4_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005403(.in0(tmp01_10_42), .in1(tmp01_11_42), .out(tmp02_5_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005404(.in0(tmp01_12_42), .in1(tmp01_13_42), .out(tmp02_6_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005405(.in0(tmp01_14_42), .in1(tmp01_15_42), .out(tmp02_7_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005406(.in0(tmp01_16_42), .in1(tmp01_17_42), .out(tmp02_8_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005407(.in0(tmp01_18_42), .in1(tmp01_19_42), .out(tmp02_9_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005408(.in0(tmp01_20_42), .in1(tmp01_21_42), .out(tmp02_10_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005409(.in0(tmp01_22_42), .in1(tmp01_23_42), .out(tmp02_11_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005410(.in0(tmp01_24_42), .in1(tmp01_25_42), .out(tmp02_12_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005411(.in0(tmp01_26_42), .in1(tmp01_27_42), .out(tmp02_13_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005412(.in0(tmp01_28_42), .in1(tmp01_29_42), .out(tmp02_14_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005413(.in0(tmp01_30_42), .in1(tmp01_31_42), .out(tmp02_15_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005414(.in0(tmp01_32_42), .in1(tmp01_33_42), .out(tmp02_16_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005415(.in0(tmp01_34_42), .in1(tmp01_35_42), .out(tmp02_17_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005416(.in0(tmp01_36_42), .in1(tmp01_37_42), .out(tmp02_18_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005417(.in0(tmp01_38_42), .in1(tmp01_39_42), .out(tmp02_19_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005418(.in0(tmp01_40_42), .in1(tmp01_41_42), .out(tmp02_20_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005419(.in0(tmp01_42_42), .in1(tmp01_43_42), .out(tmp02_21_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005420(.in0(tmp01_44_42), .in1(tmp01_45_42), .out(tmp02_22_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005421(.in0(tmp01_46_42), .in1(tmp01_47_42), .out(tmp02_23_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005422(.in0(tmp01_48_42), .in1(tmp01_49_42), .out(tmp02_24_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005423(.in0(tmp01_50_42), .in1(tmp01_51_42), .out(tmp02_25_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005424(.in0(tmp01_52_42), .in1(tmp01_53_42), .out(tmp02_26_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005425(.in0(tmp01_54_42), .in1(tmp01_55_42), .out(tmp02_27_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005426(.in0(tmp01_56_42), .in1(tmp01_57_42), .out(tmp02_28_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005427(.in0(tmp01_58_42), .in1(tmp01_59_42), .out(tmp02_29_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005428(.in0(tmp01_60_42), .in1(tmp01_61_42), .out(tmp02_30_42));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005429(.in0(tmp01_62_42), .in1(tmp01_63_42), .out(tmp02_31_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005430(.in0(tmp02_0_42), .in1(tmp02_1_42), .out(tmp03_0_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005431(.in0(tmp02_2_42), .in1(tmp02_3_42), .out(tmp03_1_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005432(.in0(tmp02_4_42), .in1(tmp02_5_42), .out(tmp03_2_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005433(.in0(tmp02_6_42), .in1(tmp02_7_42), .out(tmp03_3_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005434(.in0(tmp02_8_42), .in1(tmp02_9_42), .out(tmp03_4_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005435(.in0(tmp02_10_42), .in1(tmp02_11_42), .out(tmp03_5_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005436(.in0(tmp02_12_42), .in1(tmp02_13_42), .out(tmp03_6_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005437(.in0(tmp02_14_42), .in1(tmp02_15_42), .out(tmp03_7_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005438(.in0(tmp02_16_42), .in1(tmp02_17_42), .out(tmp03_8_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005439(.in0(tmp02_18_42), .in1(tmp02_19_42), .out(tmp03_9_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005440(.in0(tmp02_20_42), .in1(tmp02_21_42), .out(tmp03_10_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005441(.in0(tmp02_22_42), .in1(tmp02_23_42), .out(tmp03_11_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005442(.in0(tmp02_24_42), .in1(tmp02_25_42), .out(tmp03_12_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005443(.in0(tmp02_26_42), .in1(tmp02_27_42), .out(tmp03_13_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005444(.in0(tmp02_28_42), .in1(tmp02_29_42), .out(tmp03_14_42));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005445(.in0(tmp02_30_42), .in1(tmp02_31_42), .out(tmp03_15_42));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005446(.in0(tmp03_0_42), .in1(tmp03_1_42), .out(tmp04_0_42));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005447(.in0(tmp03_2_42), .in1(tmp03_3_42), .out(tmp04_1_42));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005448(.in0(tmp03_4_42), .in1(tmp03_5_42), .out(tmp04_2_42));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005449(.in0(tmp03_6_42), .in1(tmp03_7_42), .out(tmp04_3_42));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005450(.in0(tmp03_8_42), .in1(tmp03_9_42), .out(tmp04_4_42));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005451(.in0(tmp03_10_42), .in1(tmp03_11_42), .out(tmp04_5_42));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005452(.in0(tmp03_12_42), .in1(tmp03_13_42), .out(tmp04_6_42));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005453(.in0(tmp03_14_42), .in1(tmp03_15_42), .out(tmp04_7_42));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005454(.in0(tmp04_0_42), .in1(tmp04_1_42), .out(tmp05_0_42));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005455(.in0(tmp04_2_42), .in1(tmp04_3_42), .out(tmp05_1_42));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005456(.in0(tmp04_4_42), .in1(tmp04_5_42), .out(tmp05_2_42));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005457(.in0(tmp04_6_42), .in1(tmp04_7_42), .out(tmp05_3_42));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005458(.in0(tmp05_0_42), .in1(tmp05_1_42), .out(tmp06_0_42));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005459(.in0(tmp05_2_42), .in1(tmp05_3_42), .out(tmp06_1_42));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add005460(.in0(tmp06_0_42), .in1(tmp06_1_42), .out(tmp07_0_42));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005461(.in0(tmp00_0_43), .in1(tmp00_1_43), .out(tmp01_0_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005462(.in0(tmp00_2_43), .in1(tmp00_3_43), .out(tmp01_1_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005463(.in0(tmp00_4_43), .in1(tmp00_5_43), .out(tmp01_2_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005464(.in0(tmp00_6_43), .in1(tmp00_7_43), .out(tmp01_3_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005465(.in0(tmp00_8_43), .in1(tmp00_9_43), .out(tmp01_4_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005466(.in0(tmp00_10_43), .in1(tmp00_11_43), .out(tmp01_5_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005467(.in0(tmp00_12_43), .in1(tmp00_13_43), .out(tmp01_6_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005468(.in0(tmp00_14_43), .in1(tmp00_15_43), .out(tmp01_7_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005469(.in0(tmp00_16_43), .in1(tmp00_17_43), .out(tmp01_8_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005470(.in0(tmp00_18_43), .in1(tmp00_19_43), .out(tmp01_9_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005471(.in0(tmp00_20_43), .in1(tmp00_21_43), .out(tmp01_10_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005472(.in0(tmp00_22_43), .in1(tmp00_23_43), .out(tmp01_11_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005473(.in0(tmp00_24_43), .in1(tmp00_25_43), .out(tmp01_12_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005474(.in0(tmp00_26_43), .in1(tmp00_27_43), .out(tmp01_13_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005475(.in0(tmp00_28_43), .in1(tmp00_29_43), .out(tmp01_14_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005476(.in0(tmp00_30_43), .in1(tmp00_31_43), .out(tmp01_15_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005477(.in0(tmp00_32_43), .in1(tmp00_33_43), .out(tmp01_16_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005478(.in0(tmp00_34_43), .in1(tmp00_35_43), .out(tmp01_17_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005479(.in0(tmp00_36_43), .in1(tmp00_37_43), .out(tmp01_18_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005480(.in0(tmp00_38_43), .in1(tmp00_39_43), .out(tmp01_19_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005481(.in0(tmp00_40_43), .in1(tmp00_41_43), .out(tmp01_20_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005482(.in0(tmp00_42_43), .in1(tmp00_43_43), .out(tmp01_21_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005483(.in0(tmp00_44_43), .in1(tmp00_45_43), .out(tmp01_22_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005484(.in0(tmp00_46_43), .in1(tmp00_47_43), .out(tmp01_23_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005485(.in0(tmp00_48_43), .in1(tmp00_49_43), .out(tmp01_24_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005486(.in0(tmp00_50_43), .in1(tmp00_51_43), .out(tmp01_25_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005487(.in0(tmp00_52_43), .in1(tmp00_53_43), .out(tmp01_26_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005488(.in0(tmp00_54_43), .in1(tmp00_55_43), .out(tmp01_27_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005489(.in0(tmp00_56_43), .in1(tmp00_57_43), .out(tmp01_28_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005490(.in0(tmp00_58_43), .in1(tmp00_59_43), .out(tmp01_29_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005491(.in0(tmp00_60_43), .in1(tmp00_61_43), .out(tmp01_30_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005492(.in0(tmp00_62_43), .in1(tmp00_63_43), .out(tmp01_31_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005493(.in0(tmp00_64_43), .in1(tmp00_65_43), .out(tmp01_32_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005494(.in0(tmp00_66_43), .in1(tmp00_67_43), .out(tmp01_33_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005495(.in0(tmp00_68_43), .in1(tmp00_69_43), .out(tmp01_34_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005496(.in0(tmp00_70_43), .in1(tmp00_71_43), .out(tmp01_35_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005497(.in0(tmp00_72_43), .in1(tmp00_73_43), .out(tmp01_36_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005498(.in0(tmp00_74_43), .in1(tmp00_75_43), .out(tmp01_37_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005499(.in0(tmp00_76_43), .in1(tmp00_77_43), .out(tmp01_38_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005500(.in0(tmp00_78_43), .in1(tmp00_79_43), .out(tmp01_39_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005501(.in0(tmp00_80_43), .in1(tmp00_81_43), .out(tmp01_40_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005502(.in0(tmp00_82_43), .in1(tmp00_83_43), .out(tmp01_41_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005503(.in0(tmp00_84_43), .in1(tmp00_85_43), .out(tmp01_42_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005504(.in0(tmp00_86_43), .in1(tmp00_87_43), .out(tmp01_43_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005505(.in0(tmp00_88_43), .in1(tmp00_89_43), .out(tmp01_44_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005506(.in0(tmp00_90_43), .in1(tmp00_91_43), .out(tmp01_45_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005507(.in0(tmp00_92_43), .in1(tmp00_93_43), .out(tmp01_46_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005508(.in0(tmp00_94_43), .in1(tmp00_95_43), .out(tmp01_47_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005509(.in0(tmp00_96_43), .in1(tmp00_97_43), .out(tmp01_48_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005510(.in0(tmp00_98_43), .in1(tmp00_99_43), .out(tmp01_49_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005511(.in0(tmp00_100_43), .in1(tmp00_101_43), .out(tmp01_50_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005512(.in0(tmp00_102_43), .in1(tmp00_103_43), .out(tmp01_51_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005513(.in0(tmp00_104_43), .in1(tmp00_105_43), .out(tmp01_52_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005514(.in0(tmp00_106_43), .in1(tmp00_107_43), .out(tmp01_53_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005515(.in0(tmp00_108_43), .in1(tmp00_109_43), .out(tmp01_54_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005516(.in0(tmp00_110_43), .in1(tmp00_111_43), .out(tmp01_55_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005517(.in0(tmp00_112_43), .in1(tmp00_113_43), .out(tmp01_56_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005518(.in0(tmp00_114_43), .in1(tmp00_115_43), .out(tmp01_57_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005519(.in0(tmp00_116_43), .in1(tmp00_117_43), .out(tmp01_58_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005520(.in0(tmp00_118_43), .in1(tmp00_119_43), .out(tmp01_59_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005521(.in0(tmp00_120_43), .in1(tmp00_121_43), .out(tmp01_60_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005522(.in0(tmp00_122_43), .in1(tmp00_123_43), .out(tmp01_61_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005523(.in0(tmp00_124_43), .in1(tmp00_125_43), .out(tmp01_62_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005524(.in0(tmp00_126_43), .in1(tmp00_127_43), .out(tmp01_63_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005525(.in0(tmp01_0_43), .in1(tmp01_1_43), .out(tmp02_0_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005526(.in0(tmp01_2_43), .in1(tmp01_3_43), .out(tmp02_1_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005527(.in0(tmp01_4_43), .in1(tmp01_5_43), .out(tmp02_2_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005528(.in0(tmp01_6_43), .in1(tmp01_7_43), .out(tmp02_3_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005529(.in0(tmp01_8_43), .in1(tmp01_9_43), .out(tmp02_4_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005530(.in0(tmp01_10_43), .in1(tmp01_11_43), .out(tmp02_5_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005531(.in0(tmp01_12_43), .in1(tmp01_13_43), .out(tmp02_6_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005532(.in0(tmp01_14_43), .in1(tmp01_15_43), .out(tmp02_7_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005533(.in0(tmp01_16_43), .in1(tmp01_17_43), .out(tmp02_8_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005534(.in0(tmp01_18_43), .in1(tmp01_19_43), .out(tmp02_9_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005535(.in0(tmp01_20_43), .in1(tmp01_21_43), .out(tmp02_10_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005536(.in0(tmp01_22_43), .in1(tmp01_23_43), .out(tmp02_11_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005537(.in0(tmp01_24_43), .in1(tmp01_25_43), .out(tmp02_12_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005538(.in0(tmp01_26_43), .in1(tmp01_27_43), .out(tmp02_13_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005539(.in0(tmp01_28_43), .in1(tmp01_29_43), .out(tmp02_14_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005540(.in0(tmp01_30_43), .in1(tmp01_31_43), .out(tmp02_15_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005541(.in0(tmp01_32_43), .in1(tmp01_33_43), .out(tmp02_16_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005542(.in0(tmp01_34_43), .in1(tmp01_35_43), .out(tmp02_17_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005543(.in0(tmp01_36_43), .in1(tmp01_37_43), .out(tmp02_18_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005544(.in0(tmp01_38_43), .in1(tmp01_39_43), .out(tmp02_19_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005545(.in0(tmp01_40_43), .in1(tmp01_41_43), .out(tmp02_20_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005546(.in0(tmp01_42_43), .in1(tmp01_43_43), .out(tmp02_21_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005547(.in0(tmp01_44_43), .in1(tmp01_45_43), .out(tmp02_22_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005548(.in0(tmp01_46_43), .in1(tmp01_47_43), .out(tmp02_23_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005549(.in0(tmp01_48_43), .in1(tmp01_49_43), .out(tmp02_24_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005550(.in0(tmp01_50_43), .in1(tmp01_51_43), .out(tmp02_25_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005551(.in0(tmp01_52_43), .in1(tmp01_53_43), .out(tmp02_26_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005552(.in0(tmp01_54_43), .in1(tmp01_55_43), .out(tmp02_27_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005553(.in0(tmp01_56_43), .in1(tmp01_57_43), .out(tmp02_28_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005554(.in0(tmp01_58_43), .in1(tmp01_59_43), .out(tmp02_29_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005555(.in0(tmp01_60_43), .in1(tmp01_61_43), .out(tmp02_30_43));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005556(.in0(tmp01_62_43), .in1(tmp01_63_43), .out(tmp02_31_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005557(.in0(tmp02_0_43), .in1(tmp02_1_43), .out(tmp03_0_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005558(.in0(tmp02_2_43), .in1(tmp02_3_43), .out(tmp03_1_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005559(.in0(tmp02_4_43), .in1(tmp02_5_43), .out(tmp03_2_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005560(.in0(tmp02_6_43), .in1(tmp02_7_43), .out(tmp03_3_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005561(.in0(tmp02_8_43), .in1(tmp02_9_43), .out(tmp03_4_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005562(.in0(tmp02_10_43), .in1(tmp02_11_43), .out(tmp03_5_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005563(.in0(tmp02_12_43), .in1(tmp02_13_43), .out(tmp03_6_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005564(.in0(tmp02_14_43), .in1(tmp02_15_43), .out(tmp03_7_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005565(.in0(tmp02_16_43), .in1(tmp02_17_43), .out(tmp03_8_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005566(.in0(tmp02_18_43), .in1(tmp02_19_43), .out(tmp03_9_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005567(.in0(tmp02_20_43), .in1(tmp02_21_43), .out(tmp03_10_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005568(.in0(tmp02_22_43), .in1(tmp02_23_43), .out(tmp03_11_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005569(.in0(tmp02_24_43), .in1(tmp02_25_43), .out(tmp03_12_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005570(.in0(tmp02_26_43), .in1(tmp02_27_43), .out(tmp03_13_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005571(.in0(tmp02_28_43), .in1(tmp02_29_43), .out(tmp03_14_43));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005572(.in0(tmp02_30_43), .in1(tmp02_31_43), .out(tmp03_15_43));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005573(.in0(tmp03_0_43), .in1(tmp03_1_43), .out(tmp04_0_43));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005574(.in0(tmp03_2_43), .in1(tmp03_3_43), .out(tmp04_1_43));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005575(.in0(tmp03_4_43), .in1(tmp03_5_43), .out(tmp04_2_43));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005576(.in0(tmp03_6_43), .in1(tmp03_7_43), .out(tmp04_3_43));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005577(.in0(tmp03_8_43), .in1(tmp03_9_43), .out(tmp04_4_43));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005578(.in0(tmp03_10_43), .in1(tmp03_11_43), .out(tmp04_5_43));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005579(.in0(tmp03_12_43), .in1(tmp03_13_43), .out(tmp04_6_43));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005580(.in0(tmp03_14_43), .in1(tmp03_15_43), .out(tmp04_7_43));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005581(.in0(tmp04_0_43), .in1(tmp04_1_43), .out(tmp05_0_43));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005582(.in0(tmp04_2_43), .in1(tmp04_3_43), .out(tmp05_1_43));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005583(.in0(tmp04_4_43), .in1(tmp04_5_43), .out(tmp05_2_43));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005584(.in0(tmp04_6_43), .in1(tmp04_7_43), .out(tmp05_3_43));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005585(.in0(tmp05_0_43), .in1(tmp05_1_43), .out(tmp06_0_43));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005586(.in0(tmp05_2_43), .in1(tmp05_3_43), .out(tmp06_1_43));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add005587(.in0(tmp06_0_43), .in1(tmp06_1_43), .out(tmp07_0_43));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005588(.in0(tmp00_0_44), .in1(tmp00_1_44), .out(tmp01_0_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005589(.in0(tmp00_2_44), .in1(tmp00_3_44), .out(tmp01_1_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005590(.in0(tmp00_4_44), .in1(tmp00_5_44), .out(tmp01_2_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005591(.in0(tmp00_6_44), .in1(tmp00_7_44), .out(tmp01_3_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005592(.in0(tmp00_8_44), .in1(tmp00_9_44), .out(tmp01_4_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005593(.in0(tmp00_10_44), .in1(tmp00_11_44), .out(tmp01_5_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005594(.in0(tmp00_12_44), .in1(tmp00_13_44), .out(tmp01_6_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005595(.in0(tmp00_14_44), .in1(tmp00_15_44), .out(tmp01_7_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005596(.in0(tmp00_16_44), .in1(tmp00_17_44), .out(tmp01_8_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005597(.in0(tmp00_18_44), .in1(tmp00_19_44), .out(tmp01_9_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005598(.in0(tmp00_20_44), .in1(tmp00_21_44), .out(tmp01_10_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005599(.in0(tmp00_22_44), .in1(tmp00_23_44), .out(tmp01_11_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005600(.in0(tmp00_24_44), .in1(tmp00_25_44), .out(tmp01_12_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005601(.in0(tmp00_26_44), .in1(tmp00_27_44), .out(tmp01_13_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005602(.in0(tmp00_28_44), .in1(tmp00_29_44), .out(tmp01_14_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005603(.in0(tmp00_30_44), .in1(tmp00_31_44), .out(tmp01_15_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005604(.in0(tmp00_32_44), .in1(tmp00_33_44), .out(tmp01_16_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005605(.in0(tmp00_34_44), .in1(tmp00_35_44), .out(tmp01_17_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005606(.in0(tmp00_36_44), .in1(tmp00_37_44), .out(tmp01_18_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005607(.in0(tmp00_38_44), .in1(tmp00_39_44), .out(tmp01_19_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005608(.in0(tmp00_40_44), .in1(tmp00_41_44), .out(tmp01_20_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005609(.in0(tmp00_42_44), .in1(tmp00_43_44), .out(tmp01_21_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005610(.in0(tmp00_44_44), .in1(tmp00_45_44), .out(tmp01_22_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005611(.in0(tmp00_46_44), .in1(tmp00_47_44), .out(tmp01_23_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005612(.in0(tmp00_48_44), .in1(tmp00_49_44), .out(tmp01_24_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005613(.in0(tmp00_50_44), .in1(tmp00_51_44), .out(tmp01_25_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005614(.in0(tmp00_52_44), .in1(tmp00_53_44), .out(tmp01_26_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005615(.in0(tmp00_54_44), .in1(tmp00_55_44), .out(tmp01_27_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005616(.in0(tmp00_56_44), .in1(tmp00_57_44), .out(tmp01_28_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005617(.in0(tmp00_58_44), .in1(tmp00_59_44), .out(tmp01_29_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005618(.in0(tmp00_60_44), .in1(tmp00_61_44), .out(tmp01_30_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005619(.in0(tmp00_62_44), .in1(tmp00_63_44), .out(tmp01_31_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005620(.in0(tmp00_64_44), .in1(tmp00_65_44), .out(tmp01_32_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005621(.in0(tmp00_66_44), .in1(tmp00_67_44), .out(tmp01_33_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005622(.in0(tmp00_68_44), .in1(tmp00_69_44), .out(tmp01_34_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005623(.in0(tmp00_70_44), .in1(tmp00_71_44), .out(tmp01_35_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005624(.in0(tmp00_72_44), .in1(tmp00_73_44), .out(tmp01_36_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005625(.in0(tmp00_74_44), .in1(tmp00_75_44), .out(tmp01_37_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005626(.in0(tmp00_76_44), .in1(tmp00_77_44), .out(tmp01_38_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005627(.in0(tmp00_78_44), .in1(tmp00_79_44), .out(tmp01_39_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005628(.in0(tmp00_80_44), .in1(tmp00_81_44), .out(tmp01_40_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005629(.in0(tmp00_82_44), .in1(tmp00_83_44), .out(tmp01_41_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005630(.in0(tmp00_84_44), .in1(tmp00_85_44), .out(tmp01_42_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005631(.in0(tmp00_86_44), .in1(tmp00_87_44), .out(tmp01_43_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005632(.in0(tmp00_88_44), .in1(tmp00_89_44), .out(tmp01_44_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005633(.in0(tmp00_90_44), .in1(tmp00_91_44), .out(tmp01_45_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005634(.in0(tmp00_92_44), .in1(tmp00_93_44), .out(tmp01_46_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005635(.in0(tmp00_94_44), .in1(tmp00_95_44), .out(tmp01_47_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005636(.in0(tmp00_96_44), .in1(tmp00_97_44), .out(tmp01_48_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005637(.in0(tmp00_98_44), .in1(tmp00_99_44), .out(tmp01_49_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005638(.in0(tmp00_100_44), .in1(tmp00_101_44), .out(tmp01_50_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005639(.in0(tmp00_102_44), .in1(tmp00_103_44), .out(tmp01_51_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005640(.in0(tmp00_104_44), .in1(tmp00_105_44), .out(tmp01_52_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005641(.in0(tmp00_106_44), .in1(tmp00_107_44), .out(tmp01_53_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005642(.in0(tmp00_108_44), .in1(tmp00_109_44), .out(tmp01_54_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005643(.in0(tmp00_110_44), .in1(tmp00_111_44), .out(tmp01_55_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005644(.in0(tmp00_112_44), .in1(tmp00_113_44), .out(tmp01_56_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005645(.in0(tmp00_114_44), .in1(tmp00_115_44), .out(tmp01_57_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005646(.in0(tmp00_116_44), .in1(tmp00_117_44), .out(tmp01_58_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005647(.in0(tmp00_118_44), .in1(tmp00_119_44), .out(tmp01_59_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005648(.in0(tmp00_120_44), .in1(tmp00_121_44), .out(tmp01_60_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005649(.in0(tmp00_122_44), .in1(tmp00_123_44), .out(tmp01_61_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005650(.in0(tmp00_124_44), .in1(tmp00_125_44), .out(tmp01_62_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005651(.in0(tmp00_126_44), .in1(tmp00_127_44), .out(tmp01_63_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005652(.in0(tmp01_0_44), .in1(tmp01_1_44), .out(tmp02_0_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005653(.in0(tmp01_2_44), .in1(tmp01_3_44), .out(tmp02_1_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005654(.in0(tmp01_4_44), .in1(tmp01_5_44), .out(tmp02_2_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005655(.in0(tmp01_6_44), .in1(tmp01_7_44), .out(tmp02_3_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005656(.in0(tmp01_8_44), .in1(tmp01_9_44), .out(tmp02_4_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005657(.in0(tmp01_10_44), .in1(tmp01_11_44), .out(tmp02_5_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005658(.in0(tmp01_12_44), .in1(tmp01_13_44), .out(tmp02_6_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005659(.in0(tmp01_14_44), .in1(tmp01_15_44), .out(tmp02_7_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005660(.in0(tmp01_16_44), .in1(tmp01_17_44), .out(tmp02_8_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005661(.in0(tmp01_18_44), .in1(tmp01_19_44), .out(tmp02_9_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005662(.in0(tmp01_20_44), .in1(tmp01_21_44), .out(tmp02_10_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005663(.in0(tmp01_22_44), .in1(tmp01_23_44), .out(tmp02_11_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005664(.in0(tmp01_24_44), .in1(tmp01_25_44), .out(tmp02_12_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005665(.in0(tmp01_26_44), .in1(tmp01_27_44), .out(tmp02_13_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005666(.in0(tmp01_28_44), .in1(tmp01_29_44), .out(tmp02_14_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005667(.in0(tmp01_30_44), .in1(tmp01_31_44), .out(tmp02_15_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005668(.in0(tmp01_32_44), .in1(tmp01_33_44), .out(tmp02_16_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005669(.in0(tmp01_34_44), .in1(tmp01_35_44), .out(tmp02_17_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005670(.in0(tmp01_36_44), .in1(tmp01_37_44), .out(tmp02_18_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005671(.in0(tmp01_38_44), .in1(tmp01_39_44), .out(tmp02_19_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005672(.in0(tmp01_40_44), .in1(tmp01_41_44), .out(tmp02_20_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005673(.in0(tmp01_42_44), .in1(tmp01_43_44), .out(tmp02_21_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005674(.in0(tmp01_44_44), .in1(tmp01_45_44), .out(tmp02_22_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005675(.in0(tmp01_46_44), .in1(tmp01_47_44), .out(tmp02_23_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005676(.in0(tmp01_48_44), .in1(tmp01_49_44), .out(tmp02_24_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005677(.in0(tmp01_50_44), .in1(tmp01_51_44), .out(tmp02_25_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005678(.in0(tmp01_52_44), .in1(tmp01_53_44), .out(tmp02_26_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005679(.in0(tmp01_54_44), .in1(tmp01_55_44), .out(tmp02_27_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005680(.in0(tmp01_56_44), .in1(tmp01_57_44), .out(tmp02_28_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005681(.in0(tmp01_58_44), .in1(tmp01_59_44), .out(tmp02_29_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005682(.in0(tmp01_60_44), .in1(tmp01_61_44), .out(tmp02_30_44));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005683(.in0(tmp01_62_44), .in1(tmp01_63_44), .out(tmp02_31_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005684(.in0(tmp02_0_44), .in1(tmp02_1_44), .out(tmp03_0_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005685(.in0(tmp02_2_44), .in1(tmp02_3_44), .out(tmp03_1_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005686(.in0(tmp02_4_44), .in1(tmp02_5_44), .out(tmp03_2_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005687(.in0(tmp02_6_44), .in1(tmp02_7_44), .out(tmp03_3_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005688(.in0(tmp02_8_44), .in1(tmp02_9_44), .out(tmp03_4_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005689(.in0(tmp02_10_44), .in1(tmp02_11_44), .out(tmp03_5_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005690(.in0(tmp02_12_44), .in1(tmp02_13_44), .out(tmp03_6_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005691(.in0(tmp02_14_44), .in1(tmp02_15_44), .out(tmp03_7_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005692(.in0(tmp02_16_44), .in1(tmp02_17_44), .out(tmp03_8_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005693(.in0(tmp02_18_44), .in1(tmp02_19_44), .out(tmp03_9_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005694(.in0(tmp02_20_44), .in1(tmp02_21_44), .out(tmp03_10_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005695(.in0(tmp02_22_44), .in1(tmp02_23_44), .out(tmp03_11_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005696(.in0(tmp02_24_44), .in1(tmp02_25_44), .out(tmp03_12_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005697(.in0(tmp02_26_44), .in1(tmp02_27_44), .out(tmp03_13_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005698(.in0(tmp02_28_44), .in1(tmp02_29_44), .out(tmp03_14_44));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005699(.in0(tmp02_30_44), .in1(tmp02_31_44), .out(tmp03_15_44));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005700(.in0(tmp03_0_44), .in1(tmp03_1_44), .out(tmp04_0_44));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005701(.in0(tmp03_2_44), .in1(tmp03_3_44), .out(tmp04_1_44));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005702(.in0(tmp03_4_44), .in1(tmp03_5_44), .out(tmp04_2_44));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005703(.in0(tmp03_6_44), .in1(tmp03_7_44), .out(tmp04_3_44));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005704(.in0(tmp03_8_44), .in1(tmp03_9_44), .out(tmp04_4_44));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005705(.in0(tmp03_10_44), .in1(tmp03_11_44), .out(tmp04_5_44));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005706(.in0(tmp03_12_44), .in1(tmp03_13_44), .out(tmp04_6_44));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005707(.in0(tmp03_14_44), .in1(tmp03_15_44), .out(tmp04_7_44));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005708(.in0(tmp04_0_44), .in1(tmp04_1_44), .out(tmp05_0_44));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005709(.in0(tmp04_2_44), .in1(tmp04_3_44), .out(tmp05_1_44));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005710(.in0(tmp04_4_44), .in1(tmp04_5_44), .out(tmp05_2_44));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005711(.in0(tmp04_6_44), .in1(tmp04_7_44), .out(tmp05_3_44));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005712(.in0(tmp05_0_44), .in1(tmp05_1_44), .out(tmp06_0_44));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005713(.in0(tmp05_2_44), .in1(tmp05_3_44), .out(tmp06_1_44));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add005714(.in0(tmp06_0_44), .in1(tmp06_1_44), .out(tmp07_0_44));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005715(.in0(tmp00_0_45), .in1(tmp00_1_45), .out(tmp01_0_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005716(.in0(tmp00_2_45), .in1(tmp00_3_45), .out(tmp01_1_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005717(.in0(tmp00_4_45), .in1(tmp00_5_45), .out(tmp01_2_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005718(.in0(tmp00_6_45), .in1(tmp00_7_45), .out(tmp01_3_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005719(.in0(tmp00_8_45), .in1(tmp00_9_45), .out(tmp01_4_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005720(.in0(tmp00_10_45), .in1(tmp00_11_45), .out(tmp01_5_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005721(.in0(tmp00_12_45), .in1(tmp00_13_45), .out(tmp01_6_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005722(.in0(tmp00_14_45), .in1(tmp00_15_45), .out(tmp01_7_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005723(.in0(tmp00_16_45), .in1(tmp00_17_45), .out(tmp01_8_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005724(.in0(tmp00_18_45), .in1(tmp00_19_45), .out(tmp01_9_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005725(.in0(tmp00_20_45), .in1(tmp00_21_45), .out(tmp01_10_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005726(.in0(tmp00_22_45), .in1(tmp00_23_45), .out(tmp01_11_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005727(.in0(tmp00_24_45), .in1(tmp00_25_45), .out(tmp01_12_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005728(.in0(tmp00_26_45), .in1(tmp00_27_45), .out(tmp01_13_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005729(.in0(tmp00_28_45), .in1(tmp00_29_45), .out(tmp01_14_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005730(.in0(tmp00_30_45), .in1(tmp00_31_45), .out(tmp01_15_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005731(.in0(tmp00_32_45), .in1(tmp00_33_45), .out(tmp01_16_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005732(.in0(tmp00_34_45), .in1(tmp00_35_45), .out(tmp01_17_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005733(.in0(tmp00_36_45), .in1(tmp00_37_45), .out(tmp01_18_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005734(.in0(tmp00_38_45), .in1(tmp00_39_45), .out(tmp01_19_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005735(.in0(tmp00_40_45), .in1(tmp00_41_45), .out(tmp01_20_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005736(.in0(tmp00_42_45), .in1(tmp00_43_45), .out(tmp01_21_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005737(.in0(tmp00_44_45), .in1(tmp00_45_45), .out(tmp01_22_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005738(.in0(tmp00_46_45), .in1(tmp00_47_45), .out(tmp01_23_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005739(.in0(tmp00_48_45), .in1(tmp00_49_45), .out(tmp01_24_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005740(.in0(tmp00_50_45), .in1(tmp00_51_45), .out(tmp01_25_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005741(.in0(tmp00_52_45), .in1(tmp00_53_45), .out(tmp01_26_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005742(.in0(tmp00_54_45), .in1(tmp00_55_45), .out(tmp01_27_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005743(.in0(tmp00_56_45), .in1(tmp00_57_45), .out(tmp01_28_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005744(.in0(tmp00_58_45), .in1(tmp00_59_45), .out(tmp01_29_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005745(.in0(tmp00_60_45), .in1(tmp00_61_45), .out(tmp01_30_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005746(.in0(tmp00_62_45), .in1(tmp00_63_45), .out(tmp01_31_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005747(.in0(tmp00_64_45), .in1(tmp00_65_45), .out(tmp01_32_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005748(.in0(tmp00_66_45), .in1(tmp00_67_45), .out(tmp01_33_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005749(.in0(tmp00_68_45), .in1(tmp00_69_45), .out(tmp01_34_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005750(.in0(tmp00_70_45), .in1(tmp00_71_45), .out(tmp01_35_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005751(.in0(tmp00_72_45), .in1(tmp00_73_45), .out(tmp01_36_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005752(.in0(tmp00_74_45), .in1(tmp00_75_45), .out(tmp01_37_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005753(.in0(tmp00_76_45), .in1(tmp00_77_45), .out(tmp01_38_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005754(.in0(tmp00_78_45), .in1(tmp00_79_45), .out(tmp01_39_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005755(.in0(tmp00_80_45), .in1(tmp00_81_45), .out(tmp01_40_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005756(.in0(tmp00_82_45), .in1(tmp00_83_45), .out(tmp01_41_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005757(.in0(tmp00_84_45), .in1(tmp00_85_45), .out(tmp01_42_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005758(.in0(tmp00_86_45), .in1(tmp00_87_45), .out(tmp01_43_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005759(.in0(tmp00_88_45), .in1(tmp00_89_45), .out(tmp01_44_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005760(.in0(tmp00_90_45), .in1(tmp00_91_45), .out(tmp01_45_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005761(.in0(tmp00_92_45), .in1(tmp00_93_45), .out(tmp01_46_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005762(.in0(tmp00_94_45), .in1(tmp00_95_45), .out(tmp01_47_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005763(.in0(tmp00_96_45), .in1(tmp00_97_45), .out(tmp01_48_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005764(.in0(tmp00_98_45), .in1(tmp00_99_45), .out(tmp01_49_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005765(.in0(tmp00_100_45), .in1(tmp00_101_45), .out(tmp01_50_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005766(.in0(tmp00_102_45), .in1(tmp00_103_45), .out(tmp01_51_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005767(.in0(tmp00_104_45), .in1(tmp00_105_45), .out(tmp01_52_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005768(.in0(tmp00_106_45), .in1(tmp00_107_45), .out(tmp01_53_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005769(.in0(tmp00_108_45), .in1(tmp00_109_45), .out(tmp01_54_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005770(.in0(tmp00_110_45), .in1(tmp00_111_45), .out(tmp01_55_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005771(.in0(tmp00_112_45), .in1(tmp00_113_45), .out(tmp01_56_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005772(.in0(tmp00_114_45), .in1(tmp00_115_45), .out(tmp01_57_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005773(.in0(tmp00_116_45), .in1(tmp00_117_45), .out(tmp01_58_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005774(.in0(tmp00_118_45), .in1(tmp00_119_45), .out(tmp01_59_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005775(.in0(tmp00_120_45), .in1(tmp00_121_45), .out(tmp01_60_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005776(.in0(tmp00_122_45), .in1(tmp00_123_45), .out(tmp01_61_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005777(.in0(tmp00_124_45), .in1(tmp00_125_45), .out(tmp01_62_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005778(.in0(tmp00_126_45), .in1(tmp00_127_45), .out(tmp01_63_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005779(.in0(tmp01_0_45), .in1(tmp01_1_45), .out(tmp02_0_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005780(.in0(tmp01_2_45), .in1(tmp01_3_45), .out(tmp02_1_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005781(.in0(tmp01_4_45), .in1(tmp01_5_45), .out(tmp02_2_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005782(.in0(tmp01_6_45), .in1(tmp01_7_45), .out(tmp02_3_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005783(.in0(tmp01_8_45), .in1(tmp01_9_45), .out(tmp02_4_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005784(.in0(tmp01_10_45), .in1(tmp01_11_45), .out(tmp02_5_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005785(.in0(tmp01_12_45), .in1(tmp01_13_45), .out(tmp02_6_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005786(.in0(tmp01_14_45), .in1(tmp01_15_45), .out(tmp02_7_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005787(.in0(tmp01_16_45), .in1(tmp01_17_45), .out(tmp02_8_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005788(.in0(tmp01_18_45), .in1(tmp01_19_45), .out(tmp02_9_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005789(.in0(tmp01_20_45), .in1(tmp01_21_45), .out(tmp02_10_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005790(.in0(tmp01_22_45), .in1(tmp01_23_45), .out(tmp02_11_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005791(.in0(tmp01_24_45), .in1(tmp01_25_45), .out(tmp02_12_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005792(.in0(tmp01_26_45), .in1(tmp01_27_45), .out(tmp02_13_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005793(.in0(tmp01_28_45), .in1(tmp01_29_45), .out(tmp02_14_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005794(.in0(tmp01_30_45), .in1(tmp01_31_45), .out(tmp02_15_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005795(.in0(tmp01_32_45), .in1(tmp01_33_45), .out(tmp02_16_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005796(.in0(tmp01_34_45), .in1(tmp01_35_45), .out(tmp02_17_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005797(.in0(tmp01_36_45), .in1(tmp01_37_45), .out(tmp02_18_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005798(.in0(tmp01_38_45), .in1(tmp01_39_45), .out(tmp02_19_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005799(.in0(tmp01_40_45), .in1(tmp01_41_45), .out(tmp02_20_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005800(.in0(tmp01_42_45), .in1(tmp01_43_45), .out(tmp02_21_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005801(.in0(tmp01_44_45), .in1(tmp01_45_45), .out(tmp02_22_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005802(.in0(tmp01_46_45), .in1(tmp01_47_45), .out(tmp02_23_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005803(.in0(tmp01_48_45), .in1(tmp01_49_45), .out(tmp02_24_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005804(.in0(tmp01_50_45), .in1(tmp01_51_45), .out(tmp02_25_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005805(.in0(tmp01_52_45), .in1(tmp01_53_45), .out(tmp02_26_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005806(.in0(tmp01_54_45), .in1(tmp01_55_45), .out(tmp02_27_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005807(.in0(tmp01_56_45), .in1(tmp01_57_45), .out(tmp02_28_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005808(.in0(tmp01_58_45), .in1(tmp01_59_45), .out(tmp02_29_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005809(.in0(tmp01_60_45), .in1(tmp01_61_45), .out(tmp02_30_45));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005810(.in0(tmp01_62_45), .in1(tmp01_63_45), .out(tmp02_31_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005811(.in0(tmp02_0_45), .in1(tmp02_1_45), .out(tmp03_0_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005812(.in0(tmp02_2_45), .in1(tmp02_3_45), .out(tmp03_1_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005813(.in0(tmp02_4_45), .in1(tmp02_5_45), .out(tmp03_2_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005814(.in0(tmp02_6_45), .in1(tmp02_7_45), .out(tmp03_3_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005815(.in0(tmp02_8_45), .in1(tmp02_9_45), .out(tmp03_4_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005816(.in0(tmp02_10_45), .in1(tmp02_11_45), .out(tmp03_5_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005817(.in0(tmp02_12_45), .in1(tmp02_13_45), .out(tmp03_6_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005818(.in0(tmp02_14_45), .in1(tmp02_15_45), .out(tmp03_7_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005819(.in0(tmp02_16_45), .in1(tmp02_17_45), .out(tmp03_8_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005820(.in0(tmp02_18_45), .in1(tmp02_19_45), .out(tmp03_9_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005821(.in0(tmp02_20_45), .in1(tmp02_21_45), .out(tmp03_10_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005822(.in0(tmp02_22_45), .in1(tmp02_23_45), .out(tmp03_11_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005823(.in0(tmp02_24_45), .in1(tmp02_25_45), .out(tmp03_12_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005824(.in0(tmp02_26_45), .in1(tmp02_27_45), .out(tmp03_13_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005825(.in0(tmp02_28_45), .in1(tmp02_29_45), .out(tmp03_14_45));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005826(.in0(tmp02_30_45), .in1(tmp02_31_45), .out(tmp03_15_45));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005827(.in0(tmp03_0_45), .in1(tmp03_1_45), .out(tmp04_0_45));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005828(.in0(tmp03_2_45), .in1(tmp03_3_45), .out(tmp04_1_45));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005829(.in0(tmp03_4_45), .in1(tmp03_5_45), .out(tmp04_2_45));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005830(.in0(tmp03_6_45), .in1(tmp03_7_45), .out(tmp04_3_45));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005831(.in0(tmp03_8_45), .in1(tmp03_9_45), .out(tmp04_4_45));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005832(.in0(tmp03_10_45), .in1(tmp03_11_45), .out(tmp04_5_45));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005833(.in0(tmp03_12_45), .in1(tmp03_13_45), .out(tmp04_6_45));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005834(.in0(tmp03_14_45), .in1(tmp03_15_45), .out(tmp04_7_45));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005835(.in0(tmp04_0_45), .in1(tmp04_1_45), .out(tmp05_0_45));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005836(.in0(tmp04_2_45), .in1(tmp04_3_45), .out(tmp05_1_45));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005837(.in0(tmp04_4_45), .in1(tmp04_5_45), .out(tmp05_2_45));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005838(.in0(tmp04_6_45), .in1(tmp04_7_45), .out(tmp05_3_45));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005839(.in0(tmp05_0_45), .in1(tmp05_1_45), .out(tmp06_0_45));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005840(.in0(tmp05_2_45), .in1(tmp05_3_45), .out(tmp06_1_45));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add005841(.in0(tmp06_0_45), .in1(tmp06_1_45), .out(tmp07_0_45));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005842(.in0(tmp00_0_46), .in1(tmp00_1_46), .out(tmp01_0_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005843(.in0(tmp00_2_46), .in1(tmp00_3_46), .out(tmp01_1_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005844(.in0(tmp00_4_46), .in1(tmp00_5_46), .out(tmp01_2_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005845(.in0(tmp00_6_46), .in1(tmp00_7_46), .out(tmp01_3_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005846(.in0(tmp00_8_46), .in1(tmp00_9_46), .out(tmp01_4_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005847(.in0(tmp00_10_46), .in1(tmp00_11_46), .out(tmp01_5_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005848(.in0(tmp00_12_46), .in1(tmp00_13_46), .out(tmp01_6_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005849(.in0(tmp00_14_46), .in1(tmp00_15_46), .out(tmp01_7_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005850(.in0(tmp00_16_46), .in1(tmp00_17_46), .out(tmp01_8_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005851(.in0(tmp00_18_46), .in1(tmp00_19_46), .out(tmp01_9_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005852(.in0(tmp00_20_46), .in1(tmp00_21_46), .out(tmp01_10_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005853(.in0(tmp00_22_46), .in1(tmp00_23_46), .out(tmp01_11_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005854(.in0(tmp00_24_46), .in1(tmp00_25_46), .out(tmp01_12_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005855(.in0(tmp00_26_46), .in1(tmp00_27_46), .out(tmp01_13_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005856(.in0(tmp00_28_46), .in1(tmp00_29_46), .out(tmp01_14_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005857(.in0(tmp00_30_46), .in1(tmp00_31_46), .out(tmp01_15_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005858(.in0(tmp00_32_46), .in1(tmp00_33_46), .out(tmp01_16_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005859(.in0(tmp00_34_46), .in1(tmp00_35_46), .out(tmp01_17_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005860(.in0(tmp00_36_46), .in1(tmp00_37_46), .out(tmp01_18_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005861(.in0(tmp00_38_46), .in1(tmp00_39_46), .out(tmp01_19_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005862(.in0(tmp00_40_46), .in1(tmp00_41_46), .out(tmp01_20_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005863(.in0(tmp00_42_46), .in1(tmp00_43_46), .out(tmp01_21_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005864(.in0(tmp00_44_46), .in1(tmp00_45_46), .out(tmp01_22_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005865(.in0(tmp00_46_46), .in1(tmp00_47_46), .out(tmp01_23_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005866(.in0(tmp00_48_46), .in1(tmp00_49_46), .out(tmp01_24_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005867(.in0(tmp00_50_46), .in1(tmp00_51_46), .out(tmp01_25_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005868(.in0(tmp00_52_46), .in1(tmp00_53_46), .out(tmp01_26_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005869(.in0(tmp00_54_46), .in1(tmp00_55_46), .out(tmp01_27_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005870(.in0(tmp00_56_46), .in1(tmp00_57_46), .out(tmp01_28_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005871(.in0(tmp00_58_46), .in1(tmp00_59_46), .out(tmp01_29_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005872(.in0(tmp00_60_46), .in1(tmp00_61_46), .out(tmp01_30_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005873(.in0(tmp00_62_46), .in1(tmp00_63_46), .out(tmp01_31_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005874(.in0(tmp00_64_46), .in1(tmp00_65_46), .out(tmp01_32_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005875(.in0(tmp00_66_46), .in1(tmp00_67_46), .out(tmp01_33_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005876(.in0(tmp00_68_46), .in1(tmp00_69_46), .out(tmp01_34_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005877(.in0(tmp00_70_46), .in1(tmp00_71_46), .out(tmp01_35_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005878(.in0(tmp00_72_46), .in1(tmp00_73_46), .out(tmp01_36_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005879(.in0(tmp00_74_46), .in1(tmp00_75_46), .out(tmp01_37_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005880(.in0(tmp00_76_46), .in1(tmp00_77_46), .out(tmp01_38_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005881(.in0(tmp00_78_46), .in1(tmp00_79_46), .out(tmp01_39_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005882(.in0(tmp00_80_46), .in1(tmp00_81_46), .out(tmp01_40_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005883(.in0(tmp00_82_46), .in1(tmp00_83_46), .out(tmp01_41_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005884(.in0(tmp00_84_46), .in1(tmp00_85_46), .out(tmp01_42_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005885(.in0(tmp00_86_46), .in1(tmp00_87_46), .out(tmp01_43_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005886(.in0(tmp00_88_46), .in1(tmp00_89_46), .out(tmp01_44_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005887(.in0(tmp00_90_46), .in1(tmp00_91_46), .out(tmp01_45_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005888(.in0(tmp00_92_46), .in1(tmp00_93_46), .out(tmp01_46_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005889(.in0(tmp00_94_46), .in1(tmp00_95_46), .out(tmp01_47_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005890(.in0(tmp00_96_46), .in1(tmp00_97_46), .out(tmp01_48_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005891(.in0(tmp00_98_46), .in1(tmp00_99_46), .out(tmp01_49_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005892(.in0(tmp00_100_46), .in1(tmp00_101_46), .out(tmp01_50_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005893(.in0(tmp00_102_46), .in1(tmp00_103_46), .out(tmp01_51_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005894(.in0(tmp00_104_46), .in1(tmp00_105_46), .out(tmp01_52_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005895(.in0(tmp00_106_46), .in1(tmp00_107_46), .out(tmp01_53_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005896(.in0(tmp00_108_46), .in1(tmp00_109_46), .out(tmp01_54_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005897(.in0(tmp00_110_46), .in1(tmp00_111_46), .out(tmp01_55_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005898(.in0(tmp00_112_46), .in1(tmp00_113_46), .out(tmp01_56_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005899(.in0(tmp00_114_46), .in1(tmp00_115_46), .out(tmp01_57_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005900(.in0(tmp00_116_46), .in1(tmp00_117_46), .out(tmp01_58_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005901(.in0(tmp00_118_46), .in1(tmp00_119_46), .out(tmp01_59_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005902(.in0(tmp00_120_46), .in1(tmp00_121_46), .out(tmp01_60_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005903(.in0(tmp00_122_46), .in1(tmp00_123_46), .out(tmp01_61_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005904(.in0(tmp00_124_46), .in1(tmp00_125_46), .out(tmp01_62_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005905(.in0(tmp00_126_46), .in1(tmp00_127_46), .out(tmp01_63_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005906(.in0(tmp01_0_46), .in1(tmp01_1_46), .out(tmp02_0_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005907(.in0(tmp01_2_46), .in1(tmp01_3_46), .out(tmp02_1_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005908(.in0(tmp01_4_46), .in1(tmp01_5_46), .out(tmp02_2_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005909(.in0(tmp01_6_46), .in1(tmp01_7_46), .out(tmp02_3_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005910(.in0(tmp01_8_46), .in1(tmp01_9_46), .out(tmp02_4_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005911(.in0(tmp01_10_46), .in1(tmp01_11_46), .out(tmp02_5_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005912(.in0(tmp01_12_46), .in1(tmp01_13_46), .out(tmp02_6_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005913(.in0(tmp01_14_46), .in1(tmp01_15_46), .out(tmp02_7_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005914(.in0(tmp01_16_46), .in1(tmp01_17_46), .out(tmp02_8_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005915(.in0(tmp01_18_46), .in1(tmp01_19_46), .out(tmp02_9_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005916(.in0(tmp01_20_46), .in1(tmp01_21_46), .out(tmp02_10_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005917(.in0(tmp01_22_46), .in1(tmp01_23_46), .out(tmp02_11_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005918(.in0(tmp01_24_46), .in1(tmp01_25_46), .out(tmp02_12_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005919(.in0(tmp01_26_46), .in1(tmp01_27_46), .out(tmp02_13_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005920(.in0(tmp01_28_46), .in1(tmp01_29_46), .out(tmp02_14_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005921(.in0(tmp01_30_46), .in1(tmp01_31_46), .out(tmp02_15_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005922(.in0(tmp01_32_46), .in1(tmp01_33_46), .out(tmp02_16_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005923(.in0(tmp01_34_46), .in1(tmp01_35_46), .out(tmp02_17_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005924(.in0(tmp01_36_46), .in1(tmp01_37_46), .out(tmp02_18_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005925(.in0(tmp01_38_46), .in1(tmp01_39_46), .out(tmp02_19_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005926(.in0(tmp01_40_46), .in1(tmp01_41_46), .out(tmp02_20_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005927(.in0(tmp01_42_46), .in1(tmp01_43_46), .out(tmp02_21_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005928(.in0(tmp01_44_46), .in1(tmp01_45_46), .out(tmp02_22_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005929(.in0(tmp01_46_46), .in1(tmp01_47_46), .out(tmp02_23_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005930(.in0(tmp01_48_46), .in1(tmp01_49_46), .out(tmp02_24_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005931(.in0(tmp01_50_46), .in1(tmp01_51_46), .out(tmp02_25_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005932(.in0(tmp01_52_46), .in1(tmp01_53_46), .out(tmp02_26_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005933(.in0(tmp01_54_46), .in1(tmp01_55_46), .out(tmp02_27_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005934(.in0(tmp01_56_46), .in1(tmp01_57_46), .out(tmp02_28_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005935(.in0(tmp01_58_46), .in1(tmp01_59_46), .out(tmp02_29_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005936(.in0(tmp01_60_46), .in1(tmp01_61_46), .out(tmp02_30_46));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add005937(.in0(tmp01_62_46), .in1(tmp01_63_46), .out(tmp02_31_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005938(.in0(tmp02_0_46), .in1(tmp02_1_46), .out(tmp03_0_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005939(.in0(tmp02_2_46), .in1(tmp02_3_46), .out(tmp03_1_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005940(.in0(tmp02_4_46), .in1(tmp02_5_46), .out(tmp03_2_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005941(.in0(tmp02_6_46), .in1(tmp02_7_46), .out(tmp03_3_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005942(.in0(tmp02_8_46), .in1(tmp02_9_46), .out(tmp03_4_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005943(.in0(tmp02_10_46), .in1(tmp02_11_46), .out(tmp03_5_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005944(.in0(tmp02_12_46), .in1(tmp02_13_46), .out(tmp03_6_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005945(.in0(tmp02_14_46), .in1(tmp02_15_46), .out(tmp03_7_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005946(.in0(tmp02_16_46), .in1(tmp02_17_46), .out(tmp03_8_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005947(.in0(tmp02_18_46), .in1(tmp02_19_46), .out(tmp03_9_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005948(.in0(tmp02_20_46), .in1(tmp02_21_46), .out(tmp03_10_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005949(.in0(tmp02_22_46), .in1(tmp02_23_46), .out(tmp03_11_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005950(.in0(tmp02_24_46), .in1(tmp02_25_46), .out(tmp03_12_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005951(.in0(tmp02_26_46), .in1(tmp02_27_46), .out(tmp03_13_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005952(.in0(tmp02_28_46), .in1(tmp02_29_46), .out(tmp03_14_46));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add005953(.in0(tmp02_30_46), .in1(tmp02_31_46), .out(tmp03_15_46));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005954(.in0(tmp03_0_46), .in1(tmp03_1_46), .out(tmp04_0_46));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005955(.in0(tmp03_2_46), .in1(tmp03_3_46), .out(tmp04_1_46));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005956(.in0(tmp03_4_46), .in1(tmp03_5_46), .out(tmp04_2_46));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005957(.in0(tmp03_6_46), .in1(tmp03_7_46), .out(tmp04_3_46));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005958(.in0(tmp03_8_46), .in1(tmp03_9_46), .out(tmp04_4_46));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005959(.in0(tmp03_10_46), .in1(tmp03_11_46), .out(tmp04_5_46));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005960(.in0(tmp03_12_46), .in1(tmp03_13_46), .out(tmp04_6_46));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add005961(.in0(tmp03_14_46), .in1(tmp03_15_46), .out(tmp04_7_46));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005962(.in0(tmp04_0_46), .in1(tmp04_1_46), .out(tmp05_0_46));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005963(.in0(tmp04_2_46), .in1(tmp04_3_46), .out(tmp05_1_46));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005964(.in0(tmp04_4_46), .in1(tmp04_5_46), .out(tmp05_2_46));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add005965(.in0(tmp04_6_46), .in1(tmp04_7_46), .out(tmp05_3_46));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005966(.in0(tmp05_0_46), .in1(tmp05_1_46), .out(tmp06_0_46));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add005967(.in0(tmp05_2_46), .in1(tmp05_3_46), .out(tmp06_1_46));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add005968(.in0(tmp06_0_46), .in1(tmp06_1_46), .out(tmp07_0_46));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005969(.in0(tmp00_0_47), .in1(tmp00_1_47), .out(tmp01_0_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005970(.in0(tmp00_2_47), .in1(tmp00_3_47), .out(tmp01_1_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005971(.in0(tmp00_4_47), .in1(tmp00_5_47), .out(tmp01_2_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005972(.in0(tmp00_6_47), .in1(tmp00_7_47), .out(tmp01_3_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005973(.in0(tmp00_8_47), .in1(tmp00_9_47), .out(tmp01_4_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005974(.in0(tmp00_10_47), .in1(tmp00_11_47), .out(tmp01_5_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005975(.in0(tmp00_12_47), .in1(tmp00_13_47), .out(tmp01_6_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005976(.in0(tmp00_14_47), .in1(tmp00_15_47), .out(tmp01_7_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005977(.in0(tmp00_16_47), .in1(tmp00_17_47), .out(tmp01_8_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005978(.in0(tmp00_18_47), .in1(tmp00_19_47), .out(tmp01_9_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005979(.in0(tmp00_20_47), .in1(tmp00_21_47), .out(tmp01_10_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005980(.in0(tmp00_22_47), .in1(tmp00_23_47), .out(tmp01_11_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005981(.in0(tmp00_24_47), .in1(tmp00_25_47), .out(tmp01_12_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005982(.in0(tmp00_26_47), .in1(tmp00_27_47), .out(tmp01_13_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005983(.in0(tmp00_28_47), .in1(tmp00_29_47), .out(tmp01_14_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005984(.in0(tmp00_30_47), .in1(tmp00_31_47), .out(tmp01_15_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005985(.in0(tmp00_32_47), .in1(tmp00_33_47), .out(tmp01_16_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005986(.in0(tmp00_34_47), .in1(tmp00_35_47), .out(tmp01_17_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005987(.in0(tmp00_36_47), .in1(tmp00_37_47), .out(tmp01_18_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005988(.in0(tmp00_38_47), .in1(tmp00_39_47), .out(tmp01_19_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005989(.in0(tmp00_40_47), .in1(tmp00_41_47), .out(tmp01_20_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005990(.in0(tmp00_42_47), .in1(tmp00_43_47), .out(tmp01_21_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005991(.in0(tmp00_44_47), .in1(tmp00_45_47), .out(tmp01_22_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005992(.in0(tmp00_46_47), .in1(tmp00_47_47), .out(tmp01_23_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005993(.in0(tmp00_48_47), .in1(tmp00_49_47), .out(tmp01_24_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005994(.in0(tmp00_50_47), .in1(tmp00_51_47), .out(tmp01_25_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005995(.in0(tmp00_52_47), .in1(tmp00_53_47), .out(tmp01_26_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005996(.in0(tmp00_54_47), .in1(tmp00_55_47), .out(tmp01_27_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005997(.in0(tmp00_56_47), .in1(tmp00_57_47), .out(tmp01_28_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005998(.in0(tmp00_58_47), .in1(tmp00_59_47), .out(tmp01_29_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add005999(.in0(tmp00_60_47), .in1(tmp00_61_47), .out(tmp01_30_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006000(.in0(tmp00_62_47), .in1(tmp00_63_47), .out(tmp01_31_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006001(.in0(tmp00_64_47), .in1(tmp00_65_47), .out(tmp01_32_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006002(.in0(tmp00_66_47), .in1(tmp00_67_47), .out(tmp01_33_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006003(.in0(tmp00_68_47), .in1(tmp00_69_47), .out(tmp01_34_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006004(.in0(tmp00_70_47), .in1(tmp00_71_47), .out(tmp01_35_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006005(.in0(tmp00_72_47), .in1(tmp00_73_47), .out(tmp01_36_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006006(.in0(tmp00_74_47), .in1(tmp00_75_47), .out(tmp01_37_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006007(.in0(tmp00_76_47), .in1(tmp00_77_47), .out(tmp01_38_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006008(.in0(tmp00_78_47), .in1(tmp00_79_47), .out(tmp01_39_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006009(.in0(tmp00_80_47), .in1(tmp00_81_47), .out(tmp01_40_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006010(.in0(tmp00_82_47), .in1(tmp00_83_47), .out(tmp01_41_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006011(.in0(tmp00_84_47), .in1(tmp00_85_47), .out(tmp01_42_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006012(.in0(tmp00_86_47), .in1(tmp00_87_47), .out(tmp01_43_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006013(.in0(tmp00_88_47), .in1(tmp00_89_47), .out(tmp01_44_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006014(.in0(tmp00_90_47), .in1(tmp00_91_47), .out(tmp01_45_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006015(.in0(tmp00_92_47), .in1(tmp00_93_47), .out(tmp01_46_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006016(.in0(tmp00_94_47), .in1(tmp00_95_47), .out(tmp01_47_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006017(.in0(tmp00_96_47), .in1(tmp00_97_47), .out(tmp01_48_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006018(.in0(tmp00_98_47), .in1(tmp00_99_47), .out(tmp01_49_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006019(.in0(tmp00_100_47), .in1(tmp00_101_47), .out(tmp01_50_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006020(.in0(tmp00_102_47), .in1(tmp00_103_47), .out(tmp01_51_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006021(.in0(tmp00_104_47), .in1(tmp00_105_47), .out(tmp01_52_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006022(.in0(tmp00_106_47), .in1(tmp00_107_47), .out(tmp01_53_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006023(.in0(tmp00_108_47), .in1(tmp00_109_47), .out(tmp01_54_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006024(.in0(tmp00_110_47), .in1(tmp00_111_47), .out(tmp01_55_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006025(.in0(tmp00_112_47), .in1(tmp00_113_47), .out(tmp01_56_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006026(.in0(tmp00_114_47), .in1(tmp00_115_47), .out(tmp01_57_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006027(.in0(tmp00_116_47), .in1(tmp00_117_47), .out(tmp01_58_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006028(.in0(tmp00_118_47), .in1(tmp00_119_47), .out(tmp01_59_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006029(.in0(tmp00_120_47), .in1(tmp00_121_47), .out(tmp01_60_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006030(.in0(tmp00_122_47), .in1(tmp00_123_47), .out(tmp01_61_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006031(.in0(tmp00_124_47), .in1(tmp00_125_47), .out(tmp01_62_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006032(.in0(tmp00_126_47), .in1(tmp00_127_47), .out(tmp01_63_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006033(.in0(tmp01_0_47), .in1(tmp01_1_47), .out(tmp02_0_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006034(.in0(tmp01_2_47), .in1(tmp01_3_47), .out(tmp02_1_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006035(.in0(tmp01_4_47), .in1(tmp01_5_47), .out(tmp02_2_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006036(.in0(tmp01_6_47), .in1(tmp01_7_47), .out(tmp02_3_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006037(.in0(tmp01_8_47), .in1(tmp01_9_47), .out(tmp02_4_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006038(.in0(tmp01_10_47), .in1(tmp01_11_47), .out(tmp02_5_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006039(.in0(tmp01_12_47), .in1(tmp01_13_47), .out(tmp02_6_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006040(.in0(tmp01_14_47), .in1(tmp01_15_47), .out(tmp02_7_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006041(.in0(tmp01_16_47), .in1(tmp01_17_47), .out(tmp02_8_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006042(.in0(tmp01_18_47), .in1(tmp01_19_47), .out(tmp02_9_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006043(.in0(tmp01_20_47), .in1(tmp01_21_47), .out(tmp02_10_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006044(.in0(tmp01_22_47), .in1(tmp01_23_47), .out(tmp02_11_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006045(.in0(tmp01_24_47), .in1(tmp01_25_47), .out(tmp02_12_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006046(.in0(tmp01_26_47), .in1(tmp01_27_47), .out(tmp02_13_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006047(.in0(tmp01_28_47), .in1(tmp01_29_47), .out(tmp02_14_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006048(.in0(tmp01_30_47), .in1(tmp01_31_47), .out(tmp02_15_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006049(.in0(tmp01_32_47), .in1(tmp01_33_47), .out(tmp02_16_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006050(.in0(tmp01_34_47), .in1(tmp01_35_47), .out(tmp02_17_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006051(.in0(tmp01_36_47), .in1(tmp01_37_47), .out(tmp02_18_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006052(.in0(tmp01_38_47), .in1(tmp01_39_47), .out(tmp02_19_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006053(.in0(tmp01_40_47), .in1(tmp01_41_47), .out(tmp02_20_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006054(.in0(tmp01_42_47), .in1(tmp01_43_47), .out(tmp02_21_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006055(.in0(tmp01_44_47), .in1(tmp01_45_47), .out(tmp02_22_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006056(.in0(tmp01_46_47), .in1(tmp01_47_47), .out(tmp02_23_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006057(.in0(tmp01_48_47), .in1(tmp01_49_47), .out(tmp02_24_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006058(.in0(tmp01_50_47), .in1(tmp01_51_47), .out(tmp02_25_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006059(.in0(tmp01_52_47), .in1(tmp01_53_47), .out(tmp02_26_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006060(.in0(tmp01_54_47), .in1(tmp01_55_47), .out(tmp02_27_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006061(.in0(tmp01_56_47), .in1(tmp01_57_47), .out(tmp02_28_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006062(.in0(tmp01_58_47), .in1(tmp01_59_47), .out(tmp02_29_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006063(.in0(tmp01_60_47), .in1(tmp01_61_47), .out(tmp02_30_47));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006064(.in0(tmp01_62_47), .in1(tmp01_63_47), .out(tmp02_31_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006065(.in0(tmp02_0_47), .in1(tmp02_1_47), .out(tmp03_0_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006066(.in0(tmp02_2_47), .in1(tmp02_3_47), .out(tmp03_1_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006067(.in0(tmp02_4_47), .in1(tmp02_5_47), .out(tmp03_2_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006068(.in0(tmp02_6_47), .in1(tmp02_7_47), .out(tmp03_3_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006069(.in0(tmp02_8_47), .in1(tmp02_9_47), .out(tmp03_4_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006070(.in0(tmp02_10_47), .in1(tmp02_11_47), .out(tmp03_5_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006071(.in0(tmp02_12_47), .in1(tmp02_13_47), .out(tmp03_6_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006072(.in0(tmp02_14_47), .in1(tmp02_15_47), .out(tmp03_7_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006073(.in0(tmp02_16_47), .in1(tmp02_17_47), .out(tmp03_8_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006074(.in0(tmp02_18_47), .in1(tmp02_19_47), .out(tmp03_9_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006075(.in0(tmp02_20_47), .in1(tmp02_21_47), .out(tmp03_10_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006076(.in0(tmp02_22_47), .in1(tmp02_23_47), .out(tmp03_11_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006077(.in0(tmp02_24_47), .in1(tmp02_25_47), .out(tmp03_12_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006078(.in0(tmp02_26_47), .in1(tmp02_27_47), .out(tmp03_13_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006079(.in0(tmp02_28_47), .in1(tmp02_29_47), .out(tmp03_14_47));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006080(.in0(tmp02_30_47), .in1(tmp02_31_47), .out(tmp03_15_47));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006081(.in0(tmp03_0_47), .in1(tmp03_1_47), .out(tmp04_0_47));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006082(.in0(tmp03_2_47), .in1(tmp03_3_47), .out(tmp04_1_47));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006083(.in0(tmp03_4_47), .in1(tmp03_5_47), .out(tmp04_2_47));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006084(.in0(tmp03_6_47), .in1(tmp03_7_47), .out(tmp04_3_47));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006085(.in0(tmp03_8_47), .in1(tmp03_9_47), .out(tmp04_4_47));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006086(.in0(tmp03_10_47), .in1(tmp03_11_47), .out(tmp04_5_47));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006087(.in0(tmp03_12_47), .in1(tmp03_13_47), .out(tmp04_6_47));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006088(.in0(tmp03_14_47), .in1(tmp03_15_47), .out(tmp04_7_47));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006089(.in0(tmp04_0_47), .in1(tmp04_1_47), .out(tmp05_0_47));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006090(.in0(tmp04_2_47), .in1(tmp04_3_47), .out(tmp05_1_47));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006091(.in0(tmp04_4_47), .in1(tmp04_5_47), .out(tmp05_2_47));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006092(.in0(tmp04_6_47), .in1(tmp04_7_47), .out(tmp05_3_47));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006093(.in0(tmp05_0_47), .in1(tmp05_1_47), .out(tmp06_0_47));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006094(.in0(tmp05_2_47), .in1(tmp05_3_47), .out(tmp06_1_47));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add006095(.in0(tmp06_0_47), .in1(tmp06_1_47), .out(tmp07_0_47));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006096(.in0(tmp00_0_48), .in1(tmp00_1_48), .out(tmp01_0_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006097(.in0(tmp00_2_48), .in1(tmp00_3_48), .out(tmp01_1_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006098(.in0(tmp00_4_48), .in1(tmp00_5_48), .out(tmp01_2_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006099(.in0(tmp00_6_48), .in1(tmp00_7_48), .out(tmp01_3_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006100(.in0(tmp00_8_48), .in1(tmp00_9_48), .out(tmp01_4_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006101(.in0(tmp00_10_48), .in1(tmp00_11_48), .out(tmp01_5_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006102(.in0(tmp00_12_48), .in1(tmp00_13_48), .out(tmp01_6_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006103(.in0(tmp00_14_48), .in1(tmp00_15_48), .out(tmp01_7_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006104(.in0(tmp00_16_48), .in1(tmp00_17_48), .out(tmp01_8_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006105(.in0(tmp00_18_48), .in1(tmp00_19_48), .out(tmp01_9_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006106(.in0(tmp00_20_48), .in1(tmp00_21_48), .out(tmp01_10_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006107(.in0(tmp00_22_48), .in1(tmp00_23_48), .out(tmp01_11_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006108(.in0(tmp00_24_48), .in1(tmp00_25_48), .out(tmp01_12_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006109(.in0(tmp00_26_48), .in1(tmp00_27_48), .out(tmp01_13_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006110(.in0(tmp00_28_48), .in1(tmp00_29_48), .out(tmp01_14_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006111(.in0(tmp00_30_48), .in1(tmp00_31_48), .out(tmp01_15_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006112(.in0(tmp00_32_48), .in1(tmp00_33_48), .out(tmp01_16_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006113(.in0(tmp00_34_48), .in1(tmp00_35_48), .out(tmp01_17_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006114(.in0(tmp00_36_48), .in1(tmp00_37_48), .out(tmp01_18_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006115(.in0(tmp00_38_48), .in1(tmp00_39_48), .out(tmp01_19_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006116(.in0(tmp00_40_48), .in1(tmp00_41_48), .out(tmp01_20_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006117(.in0(tmp00_42_48), .in1(tmp00_43_48), .out(tmp01_21_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006118(.in0(tmp00_44_48), .in1(tmp00_45_48), .out(tmp01_22_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006119(.in0(tmp00_46_48), .in1(tmp00_47_48), .out(tmp01_23_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006120(.in0(tmp00_48_48), .in1(tmp00_49_48), .out(tmp01_24_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006121(.in0(tmp00_50_48), .in1(tmp00_51_48), .out(tmp01_25_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006122(.in0(tmp00_52_48), .in1(tmp00_53_48), .out(tmp01_26_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006123(.in0(tmp00_54_48), .in1(tmp00_55_48), .out(tmp01_27_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006124(.in0(tmp00_56_48), .in1(tmp00_57_48), .out(tmp01_28_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006125(.in0(tmp00_58_48), .in1(tmp00_59_48), .out(tmp01_29_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006126(.in0(tmp00_60_48), .in1(tmp00_61_48), .out(tmp01_30_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006127(.in0(tmp00_62_48), .in1(tmp00_63_48), .out(tmp01_31_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006128(.in0(tmp00_64_48), .in1(tmp00_65_48), .out(tmp01_32_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006129(.in0(tmp00_66_48), .in1(tmp00_67_48), .out(tmp01_33_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006130(.in0(tmp00_68_48), .in1(tmp00_69_48), .out(tmp01_34_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006131(.in0(tmp00_70_48), .in1(tmp00_71_48), .out(tmp01_35_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006132(.in0(tmp00_72_48), .in1(tmp00_73_48), .out(tmp01_36_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006133(.in0(tmp00_74_48), .in1(tmp00_75_48), .out(tmp01_37_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006134(.in0(tmp00_76_48), .in1(tmp00_77_48), .out(tmp01_38_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006135(.in0(tmp00_78_48), .in1(tmp00_79_48), .out(tmp01_39_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006136(.in0(tmp00_80_48), .in1(tmp00_81_48), .out(tmp01_40_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006137(.in0(tmp00_82_48), .in1(tmp00_83_48), .out(tmp01_41_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006138(.in0(tmp00_84_48), .in1(tmp00_85_48), .out(tmp01_42_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006139(.in0(tmp00_86_48), .in1(tmp00_87_48), .out(tmp01_43_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006140(.in0(tmp00_88_48), .in1(tmp00_89_48), .out(tmp01_44_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006141(.in0(tmp00_90_48), .in1(tmp00_91_48), .out(tmp01_45_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006142(.in0(tmp00_92_48), .in1(tmp00_93_48), .out(tmp01_46_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006143(.in0(tmp00_94_48), .in1(tmp00_95_48), .out(tmp01_47_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006144(.in0(tmp00_96_48), .in1(tmp00_97_48), .out(tmp01_48_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006145(.in0(tmp00_98_48), .in1(tmp00_99_48), .out(tmp01_49_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006146(.in0(tmp00_100_48), .in1(tmp00_101_48), .out(tmp01_50_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006147(.in0(tmp00_102_48), .in1(tmp00_103_48), .out(tmp01_51_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006148(.in0(tmp00_104_48), .in1(tmp00_105_48), .out(tmp01_52_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006149(.in0(tmp00_106_48), .in1(tmp00_107_48), .out(tmp01_53_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006150(.in0(tmp00_108_48), .in1(tmp00_109_48), .out(tmp01_54_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006151(.in0(tmp00_110_48), .in1(tmp00_111_48), .out(tmp01_55_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006152(.in0(tmp00_112_48), .in1(tmp00_113_48), .out(tmp01_56_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006153(.in0(tmp00_114_48), .in1(tmp00_115_48), .out(tmp01_57_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006154(.in0(tmp00_116_48), .in1(tmp00_117_48), .out(tmp01_58_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006155(.in0(tmp00_118_48), .in1(tmp00_119_48), .out(tmp01_59_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006156(.in0(tmp00_120_48), .in1(tmp00_121_48), .out(tmp01_60_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006157(.in0(tmp00_122_48), .in1(tmp00_123_48), .out(tmp01_61_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006158(.in0(tmp00_124_48), .in1(tmp00_125_48), .out(tmp01_62_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006159(.in0(tmp00_126_48), .in1(tmp00_127_48), .out(tmp01_63_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006160(.in0(tmp01_0_48), .in1(tmp01_1_48), .out(tmp02_0_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006161(.in0(tmp01_2_48), .in1(tmp01_3_48), .out(tmp02_1_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006162(.in0(tmp01_4_48), .in1(tmp01_5_48), .out(tmp02_2_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006163(.in0(tmp01_6_48), .in1(tmp01_7_48), .out(tmp02_3_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006164(.in0(tmp01_8_48), .in1(tmp01_9_48), .out(tmp02_4_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006165(.in0(tmp01_10_48), .in1(tmp01_11_48), .out(tmp02_5_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006166(.in0(tmp01_12_48), .in1(tmp01_13_48), .out(tmp02_6_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006167(.in0(tmp01_14_48), .in1(tmp01_15_48), .out(tmp02_7_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006168(.in0(tmp01_16_48), .in1(tmp01_17_48), .out(tmp02_8_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006169(.in0(tmp01_18_48), .in1(tmp01_19_48), .out(tmp02_9_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006170(.in0(tmp01_20_48), .in1(tmp01_21_48), .out(tmp02_10_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006171(.in0(tmp01_22_48), .in1(tmp01_23_48), .out(tmp02_11_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006172(.in0(tmp01_24_48), .in1(tmp01_25_48), .out(tmp02_12_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006173(.in0(tmp01_26_48), .in1(tmp01_27_48), .out(tmp02_13_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006174(.in0(tmp01_28_48), .in1(tmp01_29_48), .out(tmp02_14_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006175(.in0(tmp01_30_48), .in1(tmp01_31_48), .out(tmp02_15_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006176(.in0(tmp01_32_48), .in1(tmp01_33_48), .out(tmp02_16_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006177(.in0(tmp01_34_48), .in1(tmp01_35_48), .out(tmp02_17_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006178(.in0(tmp01_36_48), .in1(tmp01_37_48), .out(tmp02_18_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006179(.in0(tmp01_38_48), .in1(tmp01_39_48), .out(tmp02_19_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006180(.in0(tmp01_40_48), .in1(tmp01_41_48), .out(tmp02_20_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006181(.in0(tmp01_42_48), .in1(tmp01_43_48), .out(tmp02_21_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006182(.in0(tmp01_44_48), .in1(tmp01_45_48), .out(tmp02_22_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006183(.in0(tmp01_46_48), .in1(tmp01_47_48), .out(tmp02_23_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006184(.in0(tmp01_48_48), .in1(tmp01_49_48), .out(tmp02_24_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006185(.in0(tmp01_50_48), .in1(tmp01_51_48), .out(tmp02_25_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006186(.in0(tmp01_52_48), .in1(tmp01_53_48), .out(tmp02_26_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006187(.in0(tmp01_54_48), .in1(tmp01_55_48), .out(tmp02_27_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006188(.in0(tmp01_56_48), .in1(tmp01_57_48), .out(tmp02_28_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006189(.in0(tmp01_58_48), .in1(tmp01_59_48), .out(tmp02_29_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006190(.in0(tmp01_60_48), .in1(tmp01_61_48), .out(tmp02_30_48));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006191(.in0(tmp01_62_48), .in1(tmp01_63_48), .out(tmp02_31_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006192(.in0(tmp02_0_48), .in1(tmp02_1_48), .out(tmp03_0_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006193(.in0(tmp02_2_48), .in1(tmp02_3_48), .out(tmp03_1_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006194(.in0(tmp02_4_48), .in1(tmp02_5_48), .out(tmp03_2_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006195(.in0(tmp02_6_48), .in1(tmp02_7_48), .out(tmp03_3_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006196(.in0(tmp02_8_48), .in1(tmp02_9_48), .out(tmp03_4_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006197(.in0(tmp02_10_48), .in1(tmp02_11_48), .out(tmp03_5_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006198(.in0(tmp02_12_48), .in1(tmp02_13_48), .out(tmp03_6_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006199(.in0(tmp02_14_48), .in1(tmp02_15_48), .out(tmp03_7_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006200(.in0(tmp02_16_48), .in1(tmp02_17_48), .out(tmp03_8_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006201(.in0(tmp02_18_48), .in1(tmp02_19_48), .out(tmp03_9_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006202(.in0(tmp02_20_48), .in1(tmp02_21_48), .out(tmp03_10_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006203(.in0(tmp02_22_48), .in1(tmp02_23_48), .out(tmp03_11_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006204(.in0(tmp02_24_48), .in1(tmp02_25_48), .out(tmp03_12_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006205(.in0(tmp02_26_48), .in1(tmp02_27_48), .out(tmp03_13_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006206(.in0(tmp02_28_48), .in1(tmp02_29_48), .out(tmp03_14_48));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006207(.in0(tmp02_30_48), .in1(tmp02_31_48), .out(tmp03_15_48));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006208(.in0(tmp03_0_48), .in1(tmp03_1_48), .out(tmp04_0_48));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006209(.in0(tmp03_2_48), .in1(tmp03_3_48), .out(tmp04_1_48));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006210(.in0(tmp03_4_48), .in1(tmp03_5_48), .out(tmp04_2_48));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006211(.in0(tmp03_6_48), .in1(tmp03_7_48), .out(tmp04_3_48));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006212(.in0(tmp03_8_48), .in1(tmp03_9_48), .out(tmp04_4_48));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006213(.in0(tmp03_10_48), .in1(tmp03_11_48), .out(tmp04_5_48));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006214(.in0(tmp03_12_48), .in1(tmp03_13_48), .out(tmp04_6_48));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006215(.in0(tmp03_14_48), .in1(tmp03_15_48), .out(tmp04_7_48));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006216(.in0(tmp04_0_48), .in1(tmp04_1_48), .out(tmp05_0_48));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006217(.in0(tmp04_2_48), .in1(tmp04_3_48), .out(tmp05_1_48));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006218(.in0(tmp04_4_48), .in1(tmp04_5_48), .out(tmp05_2_48));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006219(.in0(tmp04_6_48), .in1(tmp04_7_48), .out(tmp05_3_48));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006220(.in0(tmp05_0_48), .in1(tmp05_1_48), .out(tmp06_0_48));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006221(.in0(tmp05_2_48), .in1(tmp05_3_48), .out(tmp06_1_48));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add006222(.in0(tmp06_0_48), .in1(tmp06_1_48), .out(tmp07_0_48));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006223(.in0(tmp00_0_49), .in1(tmp00_1_49), .out(tmp01_0_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006224(.in0(tmp00_2_49), .in1(tmp00_3_49), .out(tmp01_1_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006225(.in0(tmp00_4_49), .in1(tmp00_5_49), .out(tmp01_2_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006226(.in0(tmp00_6_49), .in1(tmp00_7_49), .out(tmp01_3_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006227(.in0(tmp00_8_49), .in1(tmp00_9_49), .out(tmp01_4_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006228(.in0(tmp00_10_49), .in1(tmp00_11_49), .out(tmp01_5_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006229(.in0(tmp00_12_49), .in1(tmp00_13_49), .out(tmp01_6_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006230(.in0(tmp00_14_49), .in1(tmp00_15_49), .out(tmp01_7_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006231(.in0(tmp00_16_49), .in1(tmp00_17_49), .out(tmp01_8_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006232(.in0(tmp00_18_49), .in1(tmp00_19_49), .out(tmp01_9_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006233(.in0(tmp00_20_49), .in1(tmp00_21_49), .out(tmp01_10_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006234(.in0(tmp00_22_49), .in1(tmp00_23_49), .out(tmp01_11_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006235(.in0(tmp00_24_49), .in1(tmp00_25_49), .out(tmp01_12_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006236(.in0(tmp00_26_49), .in1(tmp00_27_49), .out(tmp01_13_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006237(.in0(tmp00_28_49), .in1(tmp00_29_49), .out(tmp01_14_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006238(.in0(tmp00_30_49), .in1(tmp00_31_49), .out(tmp01_15_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006239(.in0(tmp00_32_49), .in1(tmp00_33_49), .out(tmp01_16_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006240(.in0(tmp00_34_49), .in1(tmp00_35_49), .out(tmp01_17_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006241(.in0(tmp00_36_49), .in1(tmp00_37_49), .out(tmp01_18_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006242(.in0(tmp00_38_49), .in1(tmp00_39_49), .out(tmp01_19_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006243(.in0(tmp00_40_49), .in1(tmp00_41_49), .out(tmp01_20_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006244(.in0(tmp00_42_49), .in1(tmp00_43_49), .out(tmp01_21_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006245(.in0(tmp00_44_49), .in1(tmp00_45_49), .out(tmp01_22_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006246(.in0(tmp00_46_49), .in1(tmp00_47_49), .out(tmp01_23_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006247(.in0(tmp00_48_49), .in1(tmp00_49_49), .out(tmp01_24_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006248(.in0(tmp00_50_49), .in1(tmp00_51_49), .out(tmp01_25_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006249(.in0(tmp00_52_49), .in1(tmp00_53_49), .out(tmp01_26_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006250(.in0(tmp00_54_49), .in1(tmp00_55_49), .out(tmp01_27_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006251(.in0(tmp00_56_49), .in1(tmp00_57_49), .out(tmp01_28_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006252(.in0(tmp00_58_49), .in1(tmp00_59_49), .out(tmp01_29_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006253(.in0(tmp00_60_49), .in1(tmp00_61_49), .out(tmp01_30_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006254(.in0(tmp00_62_49), .in1(tmp00_63_49), .out(tmp01_31_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006255(.in0(tmp00_64_49), .in1(tmp00_65_49), .out(tmp01_32_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006256(.in0(tmp00_66_49), .in1(tmp00_67_49), .out(tmp01_33_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006257(.in0(tmp00_68_49), .in1(tmp00_69_49), .out(tmp01_34_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006258(.in0(tmp00_70_49), .in1(tmp00_71_49), .out(tmp01_35_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006259(.in0(tmp00_72_49), .in1(tmp00_73_49), .out(tmp01_36_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006260(.in0(tmp00_74_49), .in1(tmp00_75_49), .out(tmp01_37_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006261(.in0(tmp00_76_49), .in1(tmp00_77_49), .out(tmp01_38_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006262(.in0(tmp00_78_49), .in1(tmp00_79_49), .out(tmp01_39_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006263(.in0(tmp00_80_49), .in1(tmp00_81_49), .out(tmp01_40_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006264(.in0(tmp00_82_49), .in1(tmp00_83_49), .out(tmp01_41_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006265(.in0(tmp00_84_49), .in1(tmp00_85_49), .out(tmp01_42_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006266(.in0(tmp00_86_49), .in1(tmp00_87_49), .out(tmp01_43_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006267(.in0(tmp00_88_49), .in1(tmp00_89_49), .out(tmp01_44_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006268(.in0(tmp00_90_49), .in1(tmp00_91_49), .out(tmp01_45_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006269(.in0(tmp00_92_49), .in1(tmp00_93_49), .out(tmp01_46_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006270(.in0(tmp00_94_49), .in1(tmp00_95_49), .out(tmp01_47_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006271(.in0(tmp00_96_49), .in1(tmp00_97_49), .out(tmp01_48_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006272(.in0(tmp00_98_49), .in1(tmp00_99_49), .out(tmp01_49_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006273(.in0(tmp00_100_49), .in1(tmp00_101_49), .out(tmp01_50_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006274(.in0(tmp00_102_49), .in1(tmp00_103_49), .out(tmp01_51_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006275(.in0(tmp00_104_49), .in1(tmp00_105_49), .out(tmp01_52_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006276(.in0(tmp00_106_49), .in1(tmp00_107_49), .out(tmp01_53_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006277(.in0(tmp00_108_49), .in1(tmp00_109_49), .out(tmp01_54_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006278(.in0(tmp00_110_49), .in1(tmp00_111_49), .out(tmp01_55_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006279(.in0(tmp00_112_49), .in1(tmp00_113_49), .out(tmp01_56_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006280(.in0(tmp00_114_49), .in1(tmp00_115_49), .out(tmp01_57_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006281(.in0(tmp00_116_49), .in1(tmp00_117_49), .out(tmp01_58_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006282(.in0(tmp00_118_49), .in1(tmp00_119_49), .out(tmp01_59_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006283(.in0(tmp00_120_49), .in1(tmp00_121_49), .out(tmp01_60_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006284(.in0(tmp00_122_49), .in1(tmp00_123_49), .out(tmp01_61_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006285(.in0(tmp00_124_49), .in1(tmp00_125_49), .out(tmp01_62_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006286(.in0(tmp00_126_49), .in1(tmp00_127_49), .out(tmp01_63_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006287(.in0(tmp01_0_49), .in1(tmp01_1_49), .out(tmp02_0_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006288(.in0(tmp01_2_49), .in1(tmp01_3_49), .out(tmp02_1_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006289(.in0(tmp01_4_49), .in1(tmp01_5_49), .out(tmp02_2_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006290(.in0(tmp01_6_49), .in1(tmp01_7_49), .out(tmp02_3_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006291(.in0(tmp01_8_49), .in1(tmp01_9_49), .out(tmp02_4_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006292(.in0(tmp01_10_49), .in1(tmp01_11_49), .out(tmp02_5_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006293(.in0(tmp01_12_49), .in1(tmp01_13_49), .out(tmp02_6_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006294(.in0(tmp01_14_49), .in1(tmp01_15_49), .out(tmp02_7_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006295(.in0(tmp01_16_49), .in1(tmp01_17_49), .out(tmp02_8_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006296(.in0(tmp01_18_49), .in1(tmp01_19_49), .out(tmp02_9_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006297(.in0(tmp01_20_49), .in1(tmp01_21_49), .out(tmp02_10_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006298(.in0(tmp01_22_49), .in1(tmp01_23_49), .out(tmp02_11_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006299(.in0(tmp01_24_49), .in1(tmp01_25_49), .out(tmp02_12_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006300(.in0(tmp01_26_49), .in1(tmp01_27_49), .out(tmp02_13_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006301(.in0(tmp01_28_49), .in1(tmp01_29_49), .out(tmp02_14_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006302(.in0(tmp01_30_49), .in1(tmp01_31_49), .out(tmp02_15_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006303(.in0(tmp01_32_49), .in1(tmp01_33_49), .out(tmp02_16_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006304(.in0(tmp01_34_49), .in1(tmp01_35_49), .out(tmp02_17_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006305(.in0(tmp01_36_49), .in1(tmp01_37_49), .out(tmp02_18_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006306(.in0(tmp01_38_49), .in1(tmp01_39_49), .out(tmp02_19_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006307(.in0(tmp01_40_49), .in1(tmp01_41_49), .out(tmp02_20_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006308(.in0(tmp01_42_49), .in1(tmp01_43_49), .out(tmp02_21_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006309(.in0(tmp01_44_49), .in1(tmp01_45_49), .out(tmp02_22_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006310(.in0(tmp01_46_49), .in1(tmp01_47_49), .out(tmp02_23_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006311(.in0(tmp01_48_49), .in1(tmp01_49_49), .out(tmp02_24_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006312(.in0(tmp01_50_49), .in1(tmp01_51_49), .out(tmp02_25_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006313(.in0(tmp01_52_49), .in1(tmp01_53_49), .out(tmp02_26_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006314(.in0(tmp01_54_49), .in1(tmp01_55_49), .out(tmp02_27_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006315(.in0(tmp01_56_49), .in1(tmp01_57_49), .out(tmp02_28_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006316(.in0(tmp01_58_49), .in1(tmp01_59_49), .out(tmp02_29_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006317(.in0(tmp01_60_49), .in1(tmp01_61_49), .out(tmp02_30_49));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006318(.in0(tmp01_62_49), .in1(tmp01_63_49), .out(tmp02_31_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006319(.in0(tmp02_0_49), .in1(tmp02_1_49), .out(tmp03_0_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006320(.in0(tmp02_2_49), .in1(tmp02_3_49), .out(tmp03_1_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006321(.in0(tmp02_4_49), .in1(tmp02_5_49), .out(tmp03_2_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006322(.in0(tmp02_6_49), .in1(tmp02_7_49), .out(tmp03_3_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006323(.in0(tmp02_8_49), .in1(tmp02_9_49), .out(tmp03_4_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006324(.in0(tmp02_10_49), .in1(tmp02_11_49), .out(tmp03_5_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006325(.in0(tmp02_12_49), .in1(tmp02_13_49), .out(tmp03_6_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006326(.in0(tmp02_14_49), .in1(tmp02_15_49), .out(tmp03_7_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006327(.in0(tmp02_16_49), .in1(tmp02_17_49), .out(tmp03_8_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006328(.in0(tmp02_18_49), .in1(tmp02_19_49), .out(tmp03_9_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006329(.in0(tmp02_20_49), .in1(tmp02_21_49), .out(tmp03_10_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006330(.in0(tmp02_22_49), .in1(tmp02_23_49), .out(tmp03_11_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006331(.in0(tmp02_24_49), .in1(tmp02_25_49), .out(tmp03_12_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006332(.in0(tmp02_26_49), .in1(tmp02_27_49), .out(tmp03_13_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006333(.in0(tmp02_28_49), .in1(tmp02_29_49), .out(tmp03_14_49));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006334(.in0(tmp02_30_49), .in1(tmp02_31_49), .out(tmp03_15_49));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006335(.in0(tmp03_0_49), .in1(tmp03_1_49), .out(tmp04_0_49));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006336(.in0(tmp03_2_49), .in1(tmp03_3_49), .out(tmp04_1_49));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006337(.in0(tmp03_4_49), .in1(tmp03_5_49), .out(tmp04_2_49));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006338(.in0(tmp03_6_49), .in1(tmp03_7_49), .out(tmp04_3_49));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006339(.in0(tmp03_8_49), .in1(tmp03_9_49), .out(tmp04_4_49));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006340(.in0(tmp03_10_49), .in1(tmp03_11_49), .out(tmp04_5_49));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006341(.in0(tmp03_12_49), .in1(tmp03_13_49), .out(tmp04_6_49));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006342(.in0(tmp03_14_49), .in1(tmp03_15_49), .out(tmp04_7_49));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006343(.in0(tmp04_0_49), .in1(tmp04_1_49), .out(tmp05_0_49));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006344(.in0(tmp04_2_49), .in1(tmp04_3_49), .out(tmp05_1_49));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006345(.in0(tmp04_4_49), .in1(tmp04_5_49), .out(tmp05_2_49));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006346(.in0(tmp04_6_49), .in1(tmp04_7_49), .out(tmp05_3_49));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006347(.in0(tmp05_0_49), .in1(tmp05_1_49), .out(tmp06_0_49));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006348(.in0(tmp05_2_49), .in1(tmp05_3_49), .out(tmp06_1_49));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add006349(.in0(tmp06_0_49), .in1(tmp06_1_49), .out(tmp07_0_49));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006350(.in0(tmp00_0_50), .in1(tmp00_1_50), .out(tmp01_0_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006351(.in0(tmp00_2_50), .in1(tmp00_3_50), .out(tmp01_1_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006352(.in0(tmp00_4_50), .in1(tmp00_5_50), .out(tmp01_2_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006353(.in0(tmp00_6_50), .in1(tmp00_7_50), .out(tmp01_3_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006354(.in0(tmp00_8_50), .in1(tmp00_9_50), .out(tmp01_4_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006355(.in0(tmp00_10_50), .in1(tmp00_11_50), .out(tmp01_5_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006356(.in0(tmp00_12_50), .in1(tmp00_13_50), .out(tmp01_6_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006357(.in0(tmp00_14_50), .in1(tmp00_15_50), .out(tmp01_7_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006358(.in0(tmp00_16_50), .in1(tmp00_17_50), .out(tmp01_8_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006359(.in0(tmp00_18_50), .in1(tmp00_19_50), .out(tmp01_9_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006360(.in0(tmp00_20_50), .in1(tmp00_21_50), .out(tmp01_10_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006361(.in0(tmp00_22_50), .in1(tmp00_23_50), .out(tmp01_11_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006362(.in0(tmp00_24_50), .in1(tmp00_25_50), .out(tmp01_12_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006363(.in0(tmp00_26_50), .in1(tmp00_27_50), .out(tmp01_13_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006364(.in0(tmp00_28_50), .in1(tmp00_29_50), .out(tmp01_14_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006365(.in0(tmp00_30_50), .in1(tmp00_31_50), .out(tmp01_15_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006366(.in0(tmp00_32_50), .in1(tmp00_33_50), .out(tmp01_16_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006367(.in0(tmp00_34_50), .in1(tmp00_35_50), .out(tmp01_17_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006368(.in0(tmp00_36_50), .in1(tmp00_37_50), .out(tmp01_18_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006369(.in0(tmp00_38_50), .in1(tmp00_39_50), .out(tmp01_19_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006370(.in0(tmp00_40_50), .in1(tmp00_41_50), .out(tmp01_20_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006371(.in0(tmp00_42_50), .in1(tmp00_43_50), .out(tmp01_21_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006372(.in0(tmp00_44_50), .in1(tmp00_45_50), .out(tmp01_22_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006373(.in0(tmp00_46_50), .in1(tmp00_47_50), .out(tmp01_23_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006374(.in0(tmp00_48_50), .in1(tmp00_49_50), .out(tmp01_24_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006375(.in0(tmp00_50_50), .in1(tmp00_51_50), .out(tmp01_25_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006376(.in0(tmp00_52_50), .in1(tmp00_53_50), .out(tmp01_26_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006377(.in0(tmp00_54_50), .in1(tmp00_55_50), .out(tmp01_27_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006378(.in0(tmp00_56_50), .in1(tmp00_57_50), .out(tmp01_28_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006379(.in0(tmp00_58_50), .in1(tmp00_59_50), .out(tmp01_29_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006380(.in0(tmp00_60_50), .in1(tmp00_61_50), .out(tmp01_30_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006381(.in0(tmp00_62_50), .in1(tmp00_63_50), .out(tmp01_31_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006382(.in0(tmp00_64_50), .in1(tmp00_65_50), .out(tmp01_32_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006383(.in0(tmp00_66_50), .in1(tmp00_67_50), .out(tmp01_33_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006384(.in0(tmp00_68_50), .in1(tmp00_69_50), .out(tmp01_34_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006385(.in0(tmp00_70_50), .in1(tmp00_71_50), .out(tmp01_35_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006386(.in0(tmp00_72_50), .in1(tmp00_73_50), .out(tmp01_36_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006387(.in0(tmp00_74_50), .in1(tmp00_75_50), .out(tmp01_37_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006388(.in0(tmp00_76_50), .in1(tmp00_77_50), .out(tmp01_38_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006389(.in0(tmp00_78_50), .in1(tmp00_79_50), .out(tmp01_39_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006390(.in0(tmp00_80_50), .in1(tmp00_81_50), .out(tmp01_40_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006391(.in0(tmp00_82_50), .in1(tmp00_83_50), .out(tmp01_41_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006392(.in0(tmp00_84_50), .in1(tmp00_85_50), .out(tmp01_42_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006393(.in0(tmp00_86_50), .in1(tmp00_87_50), .out(tmp01_43_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006394(.in0(tmp00_88_50), .in1(tmp00_89_50), .out(tmp01_44_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006395(.in0(tmp00_90_50), .in1(tmp00_91_50), .out(tmp01_45_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006396(.in0(tmp00_92_50), .in1(tmp00_93_50), .out(tmp01_46_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006397(.in0(tmp00_94_50), .in1(tmp00_95_50), .out(tmp01_47_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006398(.in0(tmp00_96_50), .in1(tmp00_97_50), .out(tmp01_48_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006399(.in0(tmp00_98_50), .in1(tmp00_99_50), .out(tmp01_49_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006400(.in0(tmp00_100_50), .in1(tmp00_101_50), .out(tmp01_50_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006401(.in0(tmp00_102_50), .in1(tmp00_103_50), .out(tmp01_51_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006402(.in0(tmp00_104_50), .in1(tmp00_105_50), .out(tmp01_52_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006403(.in0(tmp00_106_50), .in1(tmp00_107_50), .out(tmp01_53_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006404(.in0(tmp00_108_50), .in1(tmp00_109_50), .out(tmp01_54_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006405(.in0(tmp00_110_50), .in1(tmp00_111_50), .out(tmp01_55_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006406(.in0(tmp00_112_50), .in1(tmp00_113_50), .out(tmp01_56_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006407(.in0(tmp00_114_50), .in1(tmp00_115_50), .out(tmp01_57_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006408(.in0(tmp00_116_50), .in1(tmp00_117_50), .out(tmp01_58_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006409(.in0(tmp00_118_50), .in1(tmp00_119_50), .out(tmp01_59_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006410(.in0(tmp00_120_50), .in1(tmp00_121_50), .out(tmp01_60_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006411(.in0(tmp00_122_50), .in1(tmp00_123_50), .out(tmp01_61_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006412(.in0(tmp00_124_50), .in1(tmp00_125_50), .out(tmp01_62_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006413(.in0(tmp00_126_50), .in1(tmp00_127_50), .out(tmp01_63_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006414(.in0(tmp01_0_50), .in1(tmp01_1_50), .out(tmp02_0_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006415(.in0(tmp01_2_50), .in1(tmp01_3_50), .out(tmp02_1_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006416(.in0(tmp01_4_50), .in1(tmp01_5_50), .out(tmp02_2_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006417(.in0(tmp01_6_50), .in1(tmp01_7_50), .out(tmp02_3_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006418(.in0(tmp01_8_50), .in1(tmp01_9_50), .out(tmp02_4_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006419(.in0(tmp01_10_50), .in1(tmp01_11_50), .out(tmp02_5_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006420(.in0(tmp01_12_50), .in1(tmp01_13_50), .out(tmp02_6_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006421(.in0(tmp01_14_50), .in1(tmp01_15_50), .out(tmp02_7_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006422(.in0(tmp01_16_50), .in1(tmp01_17_50), .out(tmp02_8_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006423(.in0(tmp01_18_50), .in1(tmp01_19_50), .out(tmp02_9_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006424(.in0(tmp01_20_50), .in1(tmp01_21_50), .out(tmp02_10_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006425(.in0(tmp01_22_50), .in1(tmp01_23_50), .out(tmp02_11_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006426(.in0(tmp01_24_50), .in1(tmp01_25_50), .out(tmp02_12_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006427(.in0(tmp01_26_50), .in1(tmp01_27_50), .out(tmp02_13_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006428(.in0(tmp01_28_50), .in1(tmp01_29_50), .out(tmp02_14_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006429(.in0(tmp01_30_50), .in1(tmp01_31_50), .out(tmp02_15_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006430(.in0(tmp01_32_50), .in1(tmp01_33_50), .out(tmp02_16_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006431(.in0(tmp01_34_50), .in1(tmp01_35_50), .out(tmp02_17_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006432(.in0(tmp01_36_50), .in1(tmp01_37_50), .out(tmp02_18_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006433(.in0(tmp01_38_50), .in1(tmp01_39_50), .out(tmp02_19_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006434(.in0(tmp01_40_50), .in1(tmp01_41_50), .out(tmp02_20_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006435(.in0(tmp01_42_50), .in1(tmp01_43_50), .out(tmp02_21_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006436(.in0(tmp01_44_50), .in1(tmp01_45_50), .out(tmp02_22_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006437(.in0(tmp01_46_50), .in1(tmp01_47_50), .out(tmp02_23_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006438(.in0(tmp01_48_50), .in1(tmp01_49_50), .out(tmp02_24_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006439(.in0(tmp01_50_50), .in1(tmp01_51_50), .out(tmp02_25_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006440(.in0(tmp01_52_50), .in1(tmp01_53_50), .out(tmp02_26_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006441(.in0(tmp01_54_50), .in1(tmp01_55_50), .out(tmp02_27_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006442(.in0(tmp01_56_50), .in1(tmp01_57_50), .out(tmp02_28_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006443(.in0(tmp01_58_50), .in1(tmp01_59_50), .out(tmp02_29_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006444(.in0(tmp01_60_50), .in1(tmp01_61_50), .out(tmp02_30_50));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006445(.in0(tmp01_62_50), .in1(tmp01_63_50), .out(tmp02_31_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006446(.in0(tmp02_0_50), .in1(tmp02_1_50), .out(tmp03_0_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006447(.in0(tmp02_2_50), .in1(tmp02_3_50), .out(tmp03_1_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006448(.in0(tmp02_4_50), .in1(tmp02_5_50), .out(tmp03_2_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006449(.in0(tmp02_6_50), .in1(tmp02_7_50), .out(tmp03_3_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006450(.in0(tmp02_8_50), .in1(tmp02_9_50), .out(tmp03_4_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006451(.in0(tmp02_10_50), .in1(tmp02_11_50), .out(tmp03_5_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006452(.in0(tmp02_12_50), .in1(tmp02_13_50), .out(tmp03_6_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006453(.in0(tmp02_14_50), .in1(tmp02_15_50), .out(tmp03_7_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006454(.in0(tmp02_16_50), .in1(tmp02_17_50), .out(tmp03_8_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006455(.in0(tmp02_18_50), .in1(tmp02_19_50), .out(tmp03_9_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006456(.in0(tmp02_20_50), .in1(tmp02_21_50), .out(tmp03_10_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006457(.in0(tmp02_22_50), .in1(tmp02_23_50), .out(tmp03_11_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006458(.in0(tmp02_24_50), .in1(tmp02_25_50), .out(tmp03_12_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006459(.in0(tmp02_26_50), .in1(tmp02_27_50), .out(tmp03_13_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006460(.in0(tmp02_28_50), .in1(tmp02_29_50), .out(tmp03_14_50));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006461(.in0(tmp02_30_50), .in1(tmp02_31_50), .out(tmp03_15_50));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006462(.in0(tmp03_0_50), .in1(tmp03_1_50), .out(tmp04_0_50));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006463(.in0(tmp03_2_50), .in1(tmp03_3_50), .out(tmp04_1_50));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006464(.in0(tmp03_4_50), .in1(tmp03_5_50), .out(tmp04_2_50));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006465(.in0(tmp03_6_50), .in1(tmp03_7_50), .out(tmp04_3_50));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006466(.in0(tmp03_8_50), .in1(tmp03_9_50), .out(tmp04_4_50));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006467(.in0(tmp03_10_50), .in1(tmp03_11_50), .out(tmp04_5_50));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006468(.in0(tmp03_12_50), .in1(tmp03_13_50), .out(tmp04_6_50));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006469(.in0(tmp03_14_50), .in1(tmp03_15_50), .out(tmp04_7_50));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006470(.in0(tmp04_0_50), .in1(tmp04_1_50), .out(tmp05_0_50));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006471(.in0(tmp04_2_50), .in1(tmp04_3_50), .out(tmp05_1_50));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006472(.in0(tmp04_4_50), .in1(tmp04_5_50), .out(tmp05_2_50));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006473(.in0(tmp04_6_50), .in1(tmp04_7_50), .out(tmp05_3_50));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006474(.in0(tmp05_0_50), .in1(tmp05_1_50), .out(tmp06_0_50));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006475(.in0(tmp05_2_50), .in1(tmp05_3_50), .out(tmp06_1_50));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add006476(.in0(tmp06_0_50), .in1(tmp06_1_50), .out(tmp07_0_50));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006477(.in0(tmp00_0_51), .in1(tmp00_1_51), .out(tmp01_0_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006478(.in0(tmp00_2_51), .in1(tmp00_3_51), .out(tmp01_1_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006479(.in0(tmp00_4_51), .in1(tmp00_5_51), .out(tmp01_2_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006480(.in0(tmp00_6_51), .in1(tmp00_7_51), .out(tmp01_3_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006481(.in0(tmp00_8_51), .in1(tmp00_9_51), .out(tmp01_4_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006482(.in0(tmp00_10_51), .in1(tmp00_11_51), .out(tmp01_5_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006483(.in0(tmp00_12_51), .in1(tmp00_13_51), .out(tmp01_6_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006484(.in0(tmp00_14_51), .in1(tmp00_15_51), .out(tmp01_7_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006485(.in0(tmp00_16_51), .in1(tmp00_17_51), .out(tmp01_8_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006486(.in0(tmp00_18_51), .in1(tmp00_19_51), .out(tmp01_9_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006487(.in0(tmp00_20_51), .in1(tmp00_21_51), .out(tmp01_10_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006488(.in0(tmp00_22_51), .in1(tmp00_23_51), .out(tmp01_11_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006489(.in0(tmp00_24_51), .in1(tmp00_25_51), .out(tmp01_12_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006490(.in0(tmp00_26_51), .in1(tmp00_27_51), .out(tmp01_13_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006491(.in0(tmp00_28_51), .in1(tmp00_29_51), .out(tmp01_14_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006492(.in0(tmp00_30_51), .in1(tmp00_31_51), .out(tmp01_15_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006493(.in0(tmp00_32_51), .in1(tmp00_33_51), .out(tmp01_16_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006494(.in0(tmp00_34_51), .in1(tmp00_35_51), .out(tmp01_17_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006495(.in0(tmp00_36_51), .in1(tmp00_37_51), .out(tmp01_18_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006496(.in0(tmp00_38_51), .in1(tmp00_39_51), .out(tmp01_19_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006497(.in0(tmp00_40_51), .in1(tmp00_41_51), .out(tmp01_20_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006498(.in0(tmp00_42_51), .in1(tmp00_43_51), .out(tmp01_21_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006499(.in0(tmp00_44_51), .in1(tmp00_45_51), .out(tmp01_22_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006500(.in0(tmp00_46_51), .in1(tmp00_47_51), .out(tmp01_23_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006501(.in0(tmp00_48_51), .in1(tmp00_49_51), .out(tmp01_24_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006502(.in0(tmp00_50_51), .in1(tmp00_51_51), .out(tmp01_25_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006503(.in0(tmp00_52_51), .in1(tmp00_53_51), .out(tmp01_26_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006504(.in0(tmp00_54_51), .in1(tmp00_55_51), .out(tmp01_27_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006505(.in0(tmp00_56_51), .in1(tmp00_57_51), .out(tmp01_28_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006506(.in0(tmp00_58_51), .in1(tmp00_59_51), .out(tmp01_29_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006507(.in0(tmp00_60_51), .in1(tmp00_61_51), .out(tmp01_30_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006508(.in0(tmp00_62_51), .in1(tmp00_63_51), .out(tmp01_31_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006509(.in0(tmp00_64_51), .in1(tmp00_65_51), .out(tmp01_32_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006510(.in0(tmp00_66_51), .in1(tmp00_67_51), .out(tmp01_33_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006511(.in0(tmp00_68_51), .in1(tmp00_69_51), .out(tmp01_34_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006512(.in0(tmp00_70_51), .in1(tmp00_71_51), .out(tmp01_35_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006513(.in0(tmp00_72_51), .in1(tmp00_73_51), .out(tmp01_36_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006514(.in0(tmp00_74_51), .in1(tmp00_75_51), .out(tmp01_37_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006515(.in0(tmp00_76_51), .in1(tmp00_77_51), .out(tmp01_38_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006516(.in0(tmp00_78_51), .in1(tmp00_79_51), .out(tmp01_39_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006517(.in0(tmp00_80_51), .in1(tmp00_81_51), .out(tmp01_40_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006518(.in0(tmp00_82_51), .in1(tmp00_83_51), .out(tmp01_41_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006519(.in0(tmp00_84_51), .in1(tmp00_85_51), .out(tmp01_42_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006520(.in0(tmp00_86_51), .in1(tmp00_87_51), .out(tmp01_43_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006521(.in0(tmp00_88_51), .in1(tmp00_89_51), .out(tmp01_44_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006522(.in0(tmp00_90_51), .in1(tmp00_91_51), .out(tmp01_45_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006523(.in0(tmp00_92_51), .in1(tmp00_93_51), .out(tmp01_46_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006524(.in0(tmp00_94_51), .in1(tmp00_95_51), .out(tmp01_47_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006525(.in0(tmp00_96_51), .in1(tmp00_97_51), .out(tmp01_48_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006526(.in0(tmp00_98_51), .in1(tmp00_99_51), .out(tmp01_49_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006527(.in0(tmp00_100_51), .in1(tmp00_101_51), .out(tmp01_50_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006528(.in0(tmp00_102_51), .in1(tmp00_103_51), .out(tmp01_51_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006529(.in0(tmp00_104_51), .in1(tmp00_105_51), .out(tmp01_52_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006530(.in0(tmp00_106_51), .in1(tmp00_107_51), .out(tmp01_53_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006531(.in0(tmp00_108_51), .in1(tmp00_109_51), .out(tmp01_54_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006532(.in0(tmp00_110_51), .in1(tmp00_111_51), .out(tmp01_55_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006533(.in0(tmp00_112_51), .in1(tmp00_113_51), .out(tmp01_56_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006534(.in0(tmp00_114_51), .in1(tmp00_115_51), .out(tmp01_57_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006535(.in0(tmp00_116_51), .in1(tmp00_117_51), .out(tmp01_58_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006536(.in0(tmp00_118_51), .in1(tmp00_119_51), .out(tmp01_59_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006537(.in0(tmp00_120_51), .in1(tmp00_121_51), .out(tmp01_60_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006538(.in0(tmp00_122_51), .in1(tmp00_123_51), .out(tmp01_61_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006539(.in0(tmp00_124_51), .in1(tmp00_125_51), .out(tmp01_62_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006540(.in0(tmp00_126_51), .in1(tmp00_127_51), .out(tmp01_63_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006541(.in0(tmp01_0_51), .in1(tmp01_1_51), .out(tmp02_0_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006542(.in0(tmp01_2_51), .in1(tmp01_3_51), .out(tmp02_1_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006543(.in0(tmp01_4_51), .in1(tmp01_5_51), .out(tmp02_2_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006544(.in0(tmp01_6_51), .in1(tmp01_7_51), .out(tmp02_3_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006545(.in0(tmp01_8_51), .in1(tmp01_9_51), .out(tmp02_4_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006546(.in0(tmp01_10_51), .in1(tmp01_11_51), .out(tmp02_5_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006547(.in0(tmp01_12_51), .in1(tmp01_13_51), .out(tmp02_6_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006548(.in0(tmp01_14_51), .in1(tmp01_15_51), .out(tmp02_7_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006549(.in0(tmp01_16_51), .in1(tmp01_17_51), .out(tmp02_8_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006550(.in0(tmp01_18_51), .in1(tmp01_19_51), .out(tmp02_9_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006551(.in0(tmp01_20_51), .in1(tmp01_21_51), .out(tmp02_10_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006552(.in0(tmp01_22_51), .in1(tmp01_23_51), .out(tmp02_11_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006553(.in0(tmp01_24_51), .in1(tmp01_25_51), .out(tmp02_12_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006554(.in0(tmp01_26_51), .in1(tmp01_27_51), .out(tmp02_13_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006555(.in0(tmp01_28_51), .in1(tmp01_29_51), .out(tmp02_14_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006556(.in0(tmp01_30_51), .in1(tmp01_31_51), .out(tmp02_15_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006557(.in0(tmp01_32_51), .in1(tmp01_33_51), .out(tmp02_16_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006558(.in0(tmp01_34_51), .in1(tmp01_35_51), .out(tmp02_17_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006559(.in0(tmp01_36_51), .in1(tmp01_37_51), .out(tmp02_18_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006560(.in0(tmp01_38_51), .in1(tmp01_39_51), .out(tmp02_19_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006561(.in0(tmp01_40_51), .in1(tmp01_41_51), .out(tmp02_20_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006562(.in0(tmp01_42_51), .in1(tmp01_43_51), .out(tmp02_21_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006563(.in0(tmp01_44_51), .in1(tmp01_45_51), .out(tmp02_22_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006564(.in0(tmp01_46_51), .in1(tmp01_47_51), .out(tmp02_23_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006565(.in0(tmp01_48_51), .in1(tmp01_49_51), .out(tmp02_24_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006566(.in0(tmp01_50_51), .in1(tmp01_51_51), .out(tmp02_25_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006567(.in0(tmp01_52_51), .in1(tmp01_53_51), .out(tmp02_26_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006568(.in0(tmp01_54_51), .in1(tmp01_55_51), .out(tmp02_27_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006569(.in0(tmp01_56_51), .in1(tmp01_57_51), .out(tmp02_28_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006570(.in0(tmp01_58_51), .in1(tmp01_59_51), .out(tmp02_29_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006571(.in0(tmp01_60_51), .in1(tmp01_61_51), .out(tmp02_30_51));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006572(.in0(tmp01_62_51), .in1(tmp01_63_51), .out(tmp02_31_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006573(.in0(tmp02_0_51), .in1(tmp02_1_51), .out(tmp03_0_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006574(.in0(tmp02_2_51), .in1(tmp02_3_51), .out(tmp03_1_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006575(.in0(tmp02_4_51), .in1(tmp02_5_51), .out(tmp03_2_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006576(.in0(tmp02_6_51), .in1(tmp02_7_51), .out(tmp03_3_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006577(.in0(tmp02_8_51), .in1(tmp02_9_51), .out(tmp03_4_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006578(.in0(tmp02_10_51), .in1(tmp02_11_51), .out(tmp03_5_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006579(.in0(tmp02_12_51), .in1(tmp02_13_51), .out(tmp03_6_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006580(.in0(tmp02_14_51), .in1(tmp02_15_51), .out(tmp03_7_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006581(.in0(tmp02_16_51), .in1(tmp02_17_51), .out(tmp03_8_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006582(.in0(tmp02_18_51), .in1(tmp02_19_51), .out(tmp03_9_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006583(.in0(tmp02_20_51), .in1(tmp02_21_51), .out(tmp03_10_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006584(.in0(tmp02_22_51), .in1(tmp02_23_51), .out(tmp03_11_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006585(.in0(tmp02_24_51), .in1(tmp02_25_51), .out(tmp03_12_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006586(.in0(tmp02_26_51), .in1(tmp02_27_51), .out(tmp03_13_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006587(.in0(tmp02_28_51), .in1(tmp02_29_51), .out(tmp03_14_51));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006588(.in0(tmp02_30_51), .in1(tmp02_31_51), .out(tmp03_15_51));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006589(.in0(tmp03_0_51), .in1(tmp03_1_51), .out(tmp04_0_51));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006590(.in0(tmp03_2_51), .in1(tmp03_3_51), .out(tmp04_1_51));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006591(.in0(tmp03_4_51), .in1(tmp03_5_51), .out(tmp04_2_51));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006592(.in0(tmp03_6_51), .in1(tmp03_7_51), .out(tmp04_3_51));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006593(.in0(tmp03_8_51), .in1(tmp03_9_51), .out(tmp04_4_51));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006594(.in0(tmp03_10_51), .in1(tmp03_11_51), .out(tmp04_5_51));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006595(.in0(tmp03_12_51), .in1(tmp03_13_51), .out(tmp04_6_51));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006596(.in0(tmp03_14_51), .in1(tmp03_15_51), .out(tmp04_7_51));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006597(.in0(tmp04_0_51), .in1(tmp04_1_51), .out(tmp05_0_51));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006598(.in0(tmp04_2_51), .in1(tmp04_3_51), .out(tmp05_1_51));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006599(.in0(tmp04_4_51), .in1(tmp04_5_51), .out(tmp05_2_51));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006600(.in0(tmp04_6_51), .in1(tmp04_7_51), .out(tmp05_3_51));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006601(.in0(tmp05_0_51), .in1(tmp05_1_51), .out(tmp06_0_51));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006602(.in0(tmp05_2_51), .in1(tmp05_3_51), .out(tmp06_1_51));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add006603(.in0(tmp06_0_51), .in1(tmp06_1_51), .out(tmp07_0_51));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006604(.in0(tmp00_0_52), .in1(tmp00_1_52), .out(tmp01_0_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006605(.in0(tmp00_2_52), .in1(tmp00_3_52), .out(tmp01_1_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006606(.in0(tmp00_4_52), .in1(tmp00_5_52), .out(tmp01_2_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006607(.in0(tmp00_6_52), .in1(tmp00_7_52), .out(tmp01_3_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006608(.in0(tmp00_8_52), .in1(tmp00_9_52), .out(tmp01_4_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006609(.in0(tmp00_10_52), .in1(tmp00_11_52), .out(tmp01_5_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006610(.in0(tmp00_12_52), .in1(tmp00_13_52), .out(tmp01_6_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006611(.in0(tmp00_14_52), .in1(tmp00_15_52), .out(tmp01_7_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006612(.in0(tmp00_16_52), .in1(tmp00_17_52), .out(tmp01_8_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006613(.in0(tmp00_18_52), .in1(tmp00_19_52), .out(tmp01_9_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006614(.in0(tmp00_20_52), .in1(tmp00_21_52), .out(tmp01_10_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006615(.in0(tmp00_22_52), .in1(tmp00_23_52), .out(tmp01_11_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006616(.in0(tmp00_24_52), .in1(tmp00_25_52), .out(tmp01_12_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006617(.in0(tmp00_26_52), .in1(tmp00_27_52), .out(tmp01_13_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006618(.in0(tmp00_28_52), .in1(tmp00_29_52), .out(tmp01_14_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006619(.in0(tmp00_30_52), .in1(tmp00_31_52), .out(tmp01_15_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006620(.in0(tmp00_32_52), .in1(tmp00_33_52), .out(tmp01_16_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006621(.in0(tmp00_34_52), .in1(tmp00_35_52), .out(tmp01_17_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006622(.in0(tmp00_36_52), .in1(tmp00_37_52), .out(tmp01_18_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006623(.in0(tmp00_38_52), .in1(tmp00_39_52), .out(tmp01_19_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006624(.in0(tmp00_40_52), .in1(tmp00_41_52), .out(tmp01_20_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006625(.in0(tmp00_42_52), .in1(tmp00_43_52), .out(tmp01_21_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006626(.in0(tmp00_44_52), .in1(tmp00_45_52), .out(tmp01_22_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006627(.in0(tmp00_46_52), .in1(tmp00_47_52), .out(tmp01_23_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006628(.in0(tmp00_48_52), .in1(tmp00_49_52), .out(tmp01_24_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006629(.in0(tmp00_50_52), .in1(tmp00_51_52), .out(tmp01_25_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006630(.in0(tmp00_52_52), .in1(tmp00_53_52), .out(tmp01_26_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006631(.in0(tmp00_54_52), .in1(tmp00_55_52), .out(tmp01_27_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006632(.in0(tmp00_56_52), .in1(tmp00_57_52), .out(tmp01_28_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006633(.in0(tmp00_58_52), .in1(tmp00_59_52), .out(tmp01_29_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006634(.in0(tmp00_60_52), .in1(tmp00_61_52), .out(tmp01_30_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006635(.in0(tmp00_62_52), .in1(tmp00_63_52), .out(tmp01_31_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006636(.in0(tmp00_64_52), .in1(tmp00_65_52), .out(tmp01_32_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006637(.in0(tmp00_66_52), .in1(tmp00_67_52), .out(tmp01_33_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006638(.in0(tmp00_68_52), .in1(tmp00_69_52), .out(tmp01_34_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006639(.in0(tmp00_70_52), .in1(tmp00_71_52), .out(tmp01_35_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006640(.in0(tmp00_72_52), .in1(tmp00_73_52), .out(tmp01_36_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006641(.in0(tmp00_74_52), .in1(tmp00_75_52), .out(tmp01_37_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006642(.in0(tmp00_76_52), .in1(tmp00_77_52), .out(tmp01_38_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006643(.in0(tmp00_78_52), .in1(tmp00_79_52), .out(tmp01_39_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006644(.in0(tmp00_80_52), .in1(tmp00_81_52), .out(tmp01_40_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006645(.in0(tmp00_82_52), .in1(tmp00_83_52), .out(tmp01_41_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006646(.in0(tmp00_84_52), .in1(tmp00_85_52), .out(tmp01_42_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006647(.in0(tmp00_86_52), .in1(tmp00_87_52), .out(tmp01_43_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006648(.in0(tmp00_88_52), .in1(tmp00_89_52), .out(tmp01_44_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006649(.in0(tmp00_90_52), .in1(tmp00_91_52), .out(tmp01_45_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006650(.in0(tmp00_92_52), .in1(tmp00_93_52), .out(tmp01_46_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006651(.in0(tmp00_94_52), .in1(tmp00_95_52), .out(tmp01_47_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006652(.in0(tmp00_96_52), .in1(tmp00_97_52), .out(tmp01_48_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006653(.in0(tmp00_98_52), .in1(tmp00_99_52), .out(tmp01_49_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006654(.in0(tmp00_100_52), .in1(tmp00_101_52), .out(tmp01_50_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006655(.in0(tmp00_102_52), .in1(tmp00_103_52), .out(tmp01_51_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006656(.in0(tmp00_104_52), .in1(tmp00_105_52), .out(tmp01_52_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006657(.in0(tmp00_106_52), .in1(tmp00_107_52), .out(tmp01_53_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006658(.in0(tmp00_108_52), .in1(tmp00_109_52), .out(tmp01_54_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006659(.in0(tmp00_110_52), .in1(tmp00_111_52), .out(tmp01_55_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006660(.in0(tmp00_112_52), .in1(tmp00_113_52), .out(tmp01_56_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006661(.in0(tmp00_114_52), .in1(tmp00_115_52), .out(tmp01_57_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006662(.in0(tmp00_116_52), .in1(tmp00_117_52), .out(tmp01_58_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006663(.in0(tmp00_118_52), .in1(tmp00_119_52), .out(tmp01_59_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006664(.in0(tmp00_120_52), .in1(tmp00_121_52), .out(tmp01_60_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006665(.in0(tmp00_122_52), .in1(tmp00_123_52), .out(tmp01_61_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006666(.in0(tmp00_124_52), .in1(tmp00_125_52), .out(tmp01_62_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006667(.in0(tmp00_126_52), .in1(tmp00_127_52), .out(tmp01_63_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006668(.in0(tmp01_0_52), .in1(tmp01_1_52), .out(tmp02_0_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006669(.in0(tmp01_2_52), .in1(tmp01_3_52), .out(tmp02_1_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006670(.in0(tmp01_4_52), .in1(tmp01_5_52), .out(tmp02_2_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006671(.in0(tmp01_6_52), .in1(tmp01_7_52), .out(tmp02_3_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006672(.in0(tmp01_8_52), .in1(tmp01_9_52), .out(tmp02_4_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006673(.in0(tmp01_10_52), .in1(tmp01_11_52), .out(tmp02_5_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006674(.in0(tmp01_12_52), .in1(tmp01_13_52), .out(tmp02_6_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006675(.in0(tmp01_14_52), .in1(tmp01_15_52), .out(tmp02_7_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006676(.in0(tmp01_16_52), .in1(tmp01_17_52), .out(tmp02_8_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006677(.in0(tmp01_18_52), .in1(tmp01_19_52), .out(tmp02_9_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006678(.in0(tmp01_20_52), .in1(tmp01_21_52), .out(tmp02_10_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006679(.in0(tmp01_22_52), .in1(tmp01_23_52), .out(tmp02_11_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006680(.in0(tmp01_24_52), .in1(tmp01_25_52), .out(tmp02_12_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006681(.in0(tmp01_26_52), .in1(tmp01_27_52), .out(tmp02_13_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006682(.in0(tmp01_28_52), .in1(tmp01_29_52), .out(tmp02_14_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006683(.in0(tmp01_30_52), .in1(tmp01_31_52), .out(tmp02_15_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006684(.in0(tmp01_32_52), .in1(tmp01_33_52), .out(tmp02_16_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006685(.in0(tmp01_34_52), .in1(tmp01_35_52), .out(tmp02_17_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006686(.in0(tmp01_36_52), .in1(tmp01_37_52), .out(tmp02_18_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006687(.in0(tmp01_38_52), .in1(tmp01_39_52), .out(tmp02_19_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006688(.in0(tmp01_40_52), .in1(tmp01_41_52), .out(tmp02_20_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006689(.in0(tmp01_42_52), .in1(tmp01_43_52), .out(tmp02_21_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006690(.in0(tmp01_44_52), .in1(tmp01_45_52), .out(tmp02_22_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006691(.in0(tmp01_46_52), .in1(tmp01_47_52), .out(tmp02_23_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006692(.in0(tmp01_48_52), .in1(tmp01_49_52), .out(tmp02_24_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006693(.in0(tmp01_50_52), .in1(tmp01_51_52), .out(tmp02_25_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006694(.in0(tmp01_52_52), .in1(tmp01_53_52), .out(tmp02_26_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006695(.in0(tmp01_54_52), .in1(tmp01_55_52), .out(tmp02_27_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006696(.in0(tmp01_56_52), .in1(tmp01_57_52), .out(tmp02_28_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006697(.in0(tmp01_58_52), .in1(tmp01_59_52), .out(tmp02_29_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006698(.in0(tmp01_60_52), .in1(tmp01_61_52), .out(tmp02_30_52));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006699(.in0(tmp01_62_52), .in1(tmp01_63_52), .out(tmp02_31_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006700(.in0(tmp02_0_52), .in1(tmp02_1_52), .out(tmp03_0_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006701(.in0(tmp02_2_52), .in1(tmp02_3_52), .out(tmp03_1_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006702(.in0(tmp02_4_52), .in1(tmp02_5_52), .out(tmp03_2_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006703(.in0(tmp02_6_52), .in1(tmp02_7_52), .out(tmp03_3_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006704(.in0(tmp02_8_52), .in1(tmp02_9_52), .out(tmp03_4_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006705(.in0(tmp02_10_52), .in1(tmp02_11_52), .out(tmp03_5_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006706(.in0(tmp02_12_52), .in1(tmp02_13_52), .out(tmp03_6_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006707(.in0(tmp02_14_52), .in1(tmp02_15_52), .out(tmp03_7_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006708(.in0(tmp02_16_52), .in1(tmp02_17_52), .out(tmp03_8_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006709(.in0(tmp02_18_52), .in1(tmp02_19_52), .out(tmp03_9_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006710(.in0(tmp02_20_52), .in1(tmp02_21_52), .out(tmp03_10_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006711(.in0(tmp02_22_52), .in1(tmp02_23_52), .out(tmp03_11_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006712(.in0(tmp02_24_52), .in1(tmp02_25_52), .out(tmp03_12_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006713(.in0(tmp02_26_52), .in1(tmp02_27_52), .out(tmp03_13_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006714(.in0(tmp02_28_52), .in1(tmp02_29_52), .out(tmp03_14_52));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006715(.in0(tmp02_30_52), .in1(tmp02_31_52), .out(tmp03_15_52));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006716(.in0(tmp03_0_52), .in1(tmp03_1_52), .out(tmp04_0_52));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006717(.in0(tmp03_2_52), .in1(tmp03_3_52), .out(tmp04_1_52));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006718(.in0(tmp03_4_52), .in1(tmp03_5_52), .out(tmp04_2_52));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006719(.in0(tmp03_6_52), .in1(tmp03_7_52), .out(tmp04_3_52));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006720(.in0(tmp03_8_52), .in1(tmp03_9_52), .out(tmp04_4_52));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006721(.in0(tmp03_10_52), .in1(tmp03_11_52), .out(tmp04_5_52));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006722(.in0(tmp03_12_52), .in1(tmp03_13_52), .out(tmp04_6_52));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006723(.in0(tmp03_14_52), .in1(tmp03_15_52), .out(tmp04_7_52));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006724(.in0(tmp04_0_52), .in1(tmp04_1_52), .out(tmp05_0_52));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006725(.in0(tmp04_2_52), .in1(tmp04_3_52), .out(tmp05_1_52));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006726(.in0(tmp04_4_52), .in1(tmp04_5_52), .out(tmp05_2_52));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006727(.in0(tmp04_6_52), .in1(tmp04_7_52), .out(tmp05_3_52));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006728(.in0(tmp05_0_52), .in1(tmp05_1_52), .out(tmp06_0_52));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006729(.in0(tmp05_2_52), .in1(tmp05_3_52), .out(tmp06_1_52));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add006730(.in0(tmp06_0_52), .in1(tmp06_1_52), .out(tmp07_0_52));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006731(.in0(tmp00_0_53), .in1(tmp00_1_53), .out(tmp01_0_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006732(.in0(tmp00_2_53), .in1(tmp00_3_53), .out(tmp01_1_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006733(.in0(tmp00_4_53), .in1(tmp00_5_53), .out(tmp01_2_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006734(.in0(tmp00_6_53), .in1(tmp00_7_53), .out(tmp01_3_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006735(.in0(tmp00_8_53), .in1(tmp00_9_53), .out(tmp01_4_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006736(.in0(tmp00_10_53), .in1(tmp00_11_53), .out(tmp01_5_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006737(.in0(tmp00_12_53), .in1(tmp00_13_53), .out(tmp01_6_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006738(.in0(tmp00_14_53), .in1(tmp00_15_53), .out(tmp01_7_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006739(.in0(tmp00_16_53), .in1(tmp00_17_53), .out(tmp01_8_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006740(.in0(tmp00_18_53), .in1(tmp00_19_53), .out(tmp01_9_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006741(.in0(tmp00_20_53), .in1(tmp00_21_53), .out(tmp01_10_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006742(.in0(tmp00_22_53), .in1(tmp00_23_53), .out(tmp01_11_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006743(.in0(tmp00_24_53), .in1(tmp00_25_53), .out(tmp01_12_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006744(.in0(tmp00_26_53), .in1(tmp00_27_53), .out(tmp01_13_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006745(.in0(tmp00_28_53), .in1(tmp00_29_53), .out(tmp01_14_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006746(.in0(tmp00_30_53), .in1(tmp00_31_53), .out(tmp01_15_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006747(.in0(tmp00_32_53), .in1(tmp00_33_53), .out(tmp01_16_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006748(.in0(tmp00_34_53), .in1(tmp00_35_53), .out(tmp01_17_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006749(.in0(tmp00_36_53), .in1(tmp00_37_53), .out(tmp01_18_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006750(.in0(tmp00_38_53), .in1(tmp00_39_53), .out(tmp01_19_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006751(.in0(tmp00_40_53), .in1(tmp00_41_53), .out(tmp01_20_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006752(.in0(tmp00_42_53), .in1(tmp00_43_53), .out(tmp01_21_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006753(.in0(tmp00_44_53), .in1(tmp00_45_53), .out(tmp01_22_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006754(.in0(tmp00_46_53), .in1(tmp00_47_53), .out(tmp01_23_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006755(.in0(tmp00_48_53), .in1(tmp00_49_53), .out(tmp01_24_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006756(.in0(tmp00_50_53), .in1(tmp00_51_53), .out(tmp01_25_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006757(.in0(tmp00_52_53), .in1(tmp00_53_53), .out(tmp01_26_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006758(.in0(tmp00_54_53), .in1(tmp00_55_53), .out(tmp01_27_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006759(.in0(tmp00_56_53), .in1(tmp00_57_53), .out(tmp01_28_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006760(.in0(tmp00_58_53), .in1(tmp00_59_53), .out(tmp01_29_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006761(.in0(tmp00_60_53), .in1(tmp00_61_53), .out(tmp01_30_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006762(.in0(tmp00_62_53), .in1(tmp00_63_53), .out(tmp01_31_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006763(.in0(tmp00_64_53), .in1(tmp00_65_53), .out(tmp01_32_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006764(.in0(tmp00_66_53), .in1(tmp00_67_53), .out(tmp01_33_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006765(.in0(tmp00_68_53), .in1(tmp00_69_53), .out(tmp01_34_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006766(.in0(tmp00_70_53), .in1(tmp00_71_53), .out(tmp01_35_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006767(.in0(tmp00_72_53), .in1(tmp00_73_53), .out(tmp01_36_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006768(.in0(tmp00_74_53), .in1(tmp00_75_53), .out(tmp01_37_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006769(.in0(tmp00_76_53), .in1(tmp00_77_53), .out(tmp01_38_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006770(.in0(tmp00_78_53), .in1(tmp00_79_53), .out(tmp01_39_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006771(.in0(tmp00_80_53), .in1(tmp00_81_53), .out(tmp01_40_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006772(.in0(tmp00_82_53), .in1(tmp00_83_53), .out(tmp01_41_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006773(.in0(tmp00_84_53), .in1(tmp00_85_53), .out(tmp01_42_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006774(.in0(tmp00_86_53), .in1(tmp00_87_53), .out(tmp01_43_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006775(.in0(tmp00_88_53), .in1(tmp00_89_53), .out(tmp01_44_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006776(.in0(tmp00_90_53), .in1(tmp00_91_53), .out(tmp01_45_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006777(.in0(tmp00_92_53), .in1(tmp00_93_53), .out(tmp01_46_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006778(.in0(tmp00_94_53), .in1(tmp00_95_53), .out(tmp01_47_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006779(.in0(tmp00_96_53), .in1(tmp00_97_53), .out(tmp01_48_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006780(.in0(tmp00_98_53), .in1(tmp00_99_53), .out(tmp01_49_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006781(.in0(tmp00_100_53), .in1(tmp00_101_53), .out(tmp01_50_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006782(.in0(tmp00_102_53), .in1(tmp00_103_53), .out(tmp01_51_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006783(.in0(tmp00_104_53), .in1(tmp00_105_53), .out(tmp01_52_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006784(.in0(tmp00_106_53), .in1(tmp00_107_53), .out(tmp01_53_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006785(.in0(tmp00_108_53), .in1(tmp00_109_53), .out(tmp01_54_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006786(.in0(tmp00_110_53), .in1(tmp00_111_53), .out(tmp01_55_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006787(.in0(tmp00_112_53), .in1(tmp00_113_53), .out(tmp01_56_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006788(.in0(tmp00_114_53), .in1(tmp00_115_53), .out(tmp01_57_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006789(.in0(tmp00_116_53), .in1(tmp00_117_53), .out(tmp01_58_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006790(.in0(tmp00_118_53), .in1(tmp00_119_53), .out(tmp01_59_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006791(.in0(tmp00_120_53), .in1(tmp00_121_53), .out(tmp01_60_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006792(.in0(tmp00_122_53), .in1(tmp00_123_53), .out(tmp01_61_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006793(.in0(tmp00_124_53), .in1(tmp00_125_53), .out(tmp01_62_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006794(.in0(tmp00_126_53), .in1(tmp00_127_53), .out(tmp01_63_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006795(.in0(tmp01_0_53), .in1(tmp01_1_53), .out(tmp02_0_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006796(.in0(tmp01_2_53), .in1(tmp01_3_53), .out(tmp02_1_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006797(.in0(tmp01_4_53), .in1(tmp01_5_53), .out(tmp02_2_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006798(.in0(tmp01_6_53), .in1(tmp01_7_53), .out(tmp02_3_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006799(.in0(tmp01_8_53), .in1(tmp01_9_53), .out(tmp02_4_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006800(.in0(tmp01_10_53), .in1(tmp01_11_53), .out(tmp02_5_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006801(.in0(tmp01_12_53), .in1(tmp01_13_53), .out(tmp02_6_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006802(.in0(tmp01_14_53), .in1(tmp01_15_53), .out(tmp02_7_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006803(.in0(tmp01_16_53), .in1(tmp01_17_53), .out(tmp02_8_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006804(.in0(tmp01_18_53), .in1(tmp01_19_53), .out(tmp02_9_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006805(.in0(tmp01_20_53), .in1(tmp01_21_53), .out(tmp02_10_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006806(.in0(tmp01_22_53), .in1(tmp01_23_53), .out(tmp02_11_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006807(.in0(tmp01_24_53), .in1(tmp01_25_53), .out(tmp02_12_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006808(.in0(tmp01_26_53), .in1(tmp01_27_53), .out(tmp02_13_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006809(.in0(tmp01_28_53), .in1(tmp01_29_53), .out(tmp02_14_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006810(.in0(tmp01_30_53), .in1(tmp01_31_53), .out(tmp02_15_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006811(.in0(tmp01_32_53), .in1(tmp01_33_53), .out(tmp02_16_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006812(.in0(tmp01_34_53), .in1(tmp01_35_53), .out(tmp02_17_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006813(.in0(tmp01_36_53), .in1(tmp01_37_53), .out(tmp02_18_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006814(.in0(tmp01_38_53), .in1(tmp01_39_53), .out(tmp02_19_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006815(.in0(tmp01_40_53), .in1(tmp01_41_53), .out(tmp02_20_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006816(.in0(tmp01_42_53), .in1(tmp01_43_53), .out(tmp02_21_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006817(.in0(tmp01_44_53), .in1(tmp01_45_53), .out(tmp02_22_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006818(.in0(tmp01_46_53), .in1(tmp01_47_53), .out(tmp02_23_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006819(.in0(tmp01_48_53), .in1(tmp01_49_53), .out(tmp02_24_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006820(.in0(tmp01_50_53), .in1(tmp01_51_53), .out(tmp02_25_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006821(.in0(tmp01_52_53), .in1(tmp01_53_53), .out(tmp02_26_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006822(.in0(tmp01_54_53), .in1(tmp01_55_53), .out(tmp02_27_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006823(.in0(tmp01_56_53), .in1(tmp01_57_53), .out(tmp02_28_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006824(.in0(tmp01_58_53), .in1(tmp01_59_53), .out(tmp02_29_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006825(.in0(tmp01_60_53), .in1(tmp01_61_53), .out(tmp02_30_53));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006826(.in0(tmp01_62_53), .in1(tmp01_63_53), .out(tmp02_31_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006827(.in0(tmp02_0_53), .in1(tmp02_1_53), .out(tmp03_0_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006828(.in0(tmp02_2_53), .in1(tmp02_3_53), .out(tmp03_1_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006829(.in0(tmp02_4_53), .in1(tmp02_5_53), .out(tmp03_2_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006830(.in0(tmp02_6_53), .in1(tmp02_7_53), .out(tmp03_3_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006831(.in0(tmp02_8_53), .in1(tmp02_9_53), .out(tmp03_4_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006832(.in0(tmp02_10_53), .in1(tmp02_11_53), .out(tmp03_5_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006833(.in0(tmp02_12_53), .in1(tmp02_13_53), .out(tmp03_6_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006834(.in0(tmp02_14_53), .in1(tmp02_15_53), .out(tmp03_7_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006835(.in0(tmp02_16_53), .in1(tmp02_17_53), .out(tmp03_8_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006836(.in0(tmp02_18_53), .in1(tmp02_19_53), .out(tmp03_9_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006837(.in0(tmp02_20_53), .in1(tmp02_21_53), .out(tmp03_10_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006838(.in0(tmp02_22_53), .in1(tmp02_23_53), .out(tmp03_11_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006839(.in0(tmp02_24_53), .in1(tmp02_25_53), .out(tmp03_12_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006840(.in0(tmp02_26_53), .in1(tmp02_27_53), .out(tmp03_13_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006841(.in0(tmp02_28_53), .in1(tmp02_29_53), .out(tmp03_14_53));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006842(.in0(tmp02_30_53), .in1(tmp02_31_53), .out(tmp03_15_53));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006843(.in0(tmp03_0_53), .in1(tmp03_1_53), .out(tmp04_0_53));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006844(.in0(tmp03_2_53), .in1(tmp03_3_53), .out(tmp04_1_53));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006845(.in0(tmp03_4_53), .in1(tmp03_5_53), .out(tmp04_2_53));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006846(.in0(tmp03_6_53), .in1(tmp03_7_53), .out(tmp04_3_53));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006847(.in0(tmp03_8_53), .in1(tmp03_9_53), .out(tmp04_4_53));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006848(.in0(tmp03_10_53), .in1(tmp03_11_53), .out(tmp04_5_53));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006849(.in0(tmp03_12_53), .in1(tmp03_13_53), .out(tmp04_6_53));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006850(.in0(tmp03_14_53), .in1(tmp03_15_53), .out(tmp04_7_53));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006851(.in0(tmp04_0_53), .in1(tmp04_1_53), .out(tmp05_0_53));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006852(.in0(tmp04_2_53), .in1(tmp04_3_53), .out(tmp05_1_53));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006853(.in0(tmp04_4_53), .in1(tmp04_5_53), .out(tmp05_2_53));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006854(.in0(tmp04_6_53), .in1(tmp04_7_53), .out(tmp05_3_53));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006855(.in0(tmp05_0_53), .in1(tmp05_1_53), .out(tmp06_0_53));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006856(.in0(tmp05_2_53), .in1(tmp05_3_53), .out(tmp06_1_53));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add006857(.in0(tmp06_0_53), .in1(tmp06_1_53), .out(tmp07_0_53));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006858(.in0(tmp00_0_54), .in1(tmp00_1_54), .out(tmp01_0_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006859(.in0(tmp00_2_54), .in1(tmp00_3_54), .out(tmp01_1_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006860(.in0(tmp00_4_54), .in1(tmp00_5_54), .out(tmp01_2_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006861(.in0(tmp00_6_54), .in1(tmp00_7_54), .out(tmp01_3_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006862(.in0(tmp00_8_54), .in1(tmp00_9_54), .out(tmp01_4_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006863(.in0(tmp00_10_54), .in1(tmp00_11_54), .out(tmp01_5_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006864(.in0(tmp00_12_54), .in1(tmp00_13_54), .out(tmp01_6_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006865(.in0(tmp00_14_54), .in1(tmp00_15_54), .out(tmp01_7_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006866(.in0(tmp00_16_54), .in1(tmp00_17_54), .out(tmp01_8_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006867(.in0(tmp00_18_54), .in1(tmp00_19_54), .out(tmp01_9_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006868(.in0(tmp00_20_54), .in1(tmp00_21_54), .out(tmp01_10_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006869(.in0(tmp00_22_54), .in1(tmp00_23_54), .out(tmp01_11_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006870(.in0(tmp00_24_54), .in1(tmp00_25_54), .out(tmp01_12_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006871(.in0(tmp00_26_54), .in1(tmp00_27_54), .out(tmp01_13_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006872(.in0(tmp00_28_54), .in1(tmp00_29_54), .out(tmp01_14_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006873(.in0(tmp00_30_54), .in1(tmp00_31_54), .out(tmp01_15_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006874(.in0(tmp00_32_54), .in1(tmp00_33_54), .out(tmp01_16_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006875(.in0(tmp00_34_54), .in1(tmp00_35_54), .out(tmp01_17_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006876(.in0(tmp00_36_54), .in1(tmp00_37_54), .out(tmp01_18_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006877(.in0(tmp00_38_54), .in1(tmp00_39_54), .out(tmp01_19_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006878(.in0(tmp00_40_54), .in1(tmp00_41_54), .out(tmp01_20_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006879(.in0(tmp00_42_54), .in1(tmp00_43_54), .out(tmp01_21_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006880(.in0(tmp00_44_54), .in1(tmp00_45_54), .out(tmp01_22_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006881(.in0(tmp00_46_54), .in1(tmp00_47_54), .out(tmp01_23_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006882(.in0(tmp00_48_54), .in1(tmp00_49_54), .out(tmp01_24_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006883(.in0(tmp00_50_54), .in1(tmp00_51_54), .out(tmp01_25_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006884(.in0(tmp00_52_54), .in1(tmp00_53_54), .out(tmp01_26_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006885(.in0(tmp00_54_54), .in1(tmp00_55_54), .out(tmp01_27_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006886(.in0(tmp00_56_54), .in1(tmp00_57_54), .out(tmp01_28_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006887(.in0(tmp00_58_54), .in1(tmp00_59_54), .out(tmp01_29_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006888(.in0(tmp00_60_54), .in1(tmp00_61_54), .out(tmp01_30_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006889(.in0(tmp00_62_54), .in1(tmp00_63_54), .out(tmp01_31_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006890(.in0(tmp00_64_54), .in1(tmp00_65_54), .out(tmp01_32_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006891(.in0(tmp00_66_54), .in1(tmp00_67_54), .out(tmp01_33_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006892(.in0(tmp00_68_54), .in1(tmp00_69_54), .out(tmp01_34_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006893(.in0(tmp00_70_54), .in1(tmp00_71_54), .out(tmp01_35_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006894(.in0(tmp00_72_54), .in1(tmp00_73_54), .out(tmp01_36_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006895(.in0(tmp00_74_54), .in1(tmp00_75_54), .out(tmp01_37_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006896(.in0(tmp00_76_54), .in1(tmp00_77_54), .out(tmp01_38_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006897(.in0(tmp00_78_54), .in1(tmp00_79_54), .out(tmp01_39_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006898(.in0(tmp00_80_54), .in1(tmp00_81_54), .out(tmp01_40_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006899(.in0(tmp00_82_54), .in1(tmp00_83_54), .out(tmp01_41_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006900(.in0(tmp00_84_54), .in1(tmp00_85_54), .out(tmp01_42_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006901(.in0(tmp00_86_54), .in1(tmp00_87_54), .out(tmp01_43_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006902(.in0(tmp00_88_54), .in1(tmp00_89_54), .out(tmp01_44_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006903(.in0(tmp00_90_54), .in1(tmp00_91_54), .out(tmp01_45_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006904(.in0(tmp00_92_54), .in1(tmp00_93_54), .out(tmp01_46_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006905(.in0(tmp00_94_54), .in1(tmp00_95_54), .out(tmp01_47_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006906(.in0(tmp00_96_54), .in1(tmp00_97_54), .out(tmp01_48_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006907(.in0(tmp00_98_54), .in1(tmp00_99_54), .out(tmp01_49_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006908(.in0(tmp00_100_54), .in1(tmp00_101_54), .out(tmp01_50_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006909(.in0(tmp00_102_54), .in1(tmp00_103_54), .out(tmp01_51_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006910(.in0(tmp00_104_54), .in1(tmp00_105_54), .out(tmp01_52_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006911(.in0(tmp00_106_54), .in1(tmp00_107_54), .out(tmp01_53_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006912(.in0(tmp00_108_54), .in1(tmp00_109_54), .out(tmp01_54_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006913(.in0(tmp00_110_54), .in1(tmp00_111_54), .out(tmp01_55_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006914(.in0(tmp00_112_54), .in1(tmp00_113_54), .out(tmp01_56_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006915(.in0(tmp00_114_54), .in1(tmp00_115_54), .out(tmp01_57_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006916(.in0(tmp00_116_54), .in1(tmp00_117_54), .out(tmp01_58_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006917(.in0(tmp00_118_54), .in1(tmp00_119_54), .out(tmp01_59_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006918(.in0(tmp00_120_54), .in1(tmp00_121_54), .out(tmp01_60_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006919(.in0(tmp00_122_54), .in1(tmp00_123_54), .out(tmp01_61_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006920(.in0(tmp00_124_54), .in1(tmp00_125_54), .out(tmp01_62_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006921(.in0(tmp00_126_54), .in1(tmp00_127_54), .out(tmp01_63_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006922(.in0(tmp01_0_54), .in1(tmp01_1_54), .out(tmp02_0_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006923(.in0(tmp01_2_54), .in1(tmp01_3_54), .out(tmp02_1_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006924(.in0(tmp01_4_54), .in1(tmp01_5_54), .out(tmp02_2_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006925(.in0(tmp01_6_54), .in1(tmp01_7_54), .out(tmp02_3_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006926(.in0(tmp01_8_54), .in1(tmp01_9_54), .out(tmp02_4_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006927(.in0(tmp01_10_54), .in1(tmp01_11_54), .out(tmp02_5_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006928(.in0(tmp01_12_54), .in1(tmp01_13_54), .out(tmp02_6_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006929(.in0(tmp01_14_54), .in1(tmp01_15_54), .out(tmp02_7_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006930(.in0(tmp01_16_54), .in1(tmp01_17_54), .out(tmp02_8_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006931(.in0(tmp01_18_54), .in1(tmp01_19_54), .out(tmp02_9_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006932(.in0(tmp01_20_54), .in1(tmp01_21_54), .out(tmp02_10_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006933(.in0(tmp01_22_54), .in1(tmp01_23_54), .out(tmp02_11_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006934(.in0(tmp01_24_54), .in1(tmp01_25_54), .out(tmp02_12_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006935(.in0(tmp01_26_54), .in1(tmp01_27_54), .out(tmp02_13_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006936(.in0(tmp01_28_54), .in1(tmp01_29_54), .out(tmp02_14_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006937(.in0(tmp01_30_54), .in1(tmp01_31_54), .out(tmp02_15_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006938(.in0(tmp01_32_54), .in1(tmp01_33_54), .out(tmp02_16_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006939(.in0(tmp01_34_54), .in1(tmp01_35_54), .out(tmp02_17_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006940(.in0(tmp01_36_54), .in1(tmp01_37_54), .out(tmp02_18_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006941(.in0(tmp01_38_54), .in1(tmp01_39_54), .out(tmp02_19_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006942(.in0(tmp01_40_54), .in1(tmp01_41_54), .out(tmp02_20_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006943(.in0(tmp01_42_54), .in1(tmp01_43_54), .out(tmp02_21_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006944(.in0(tmp01_44_54), .in1(tmp01_45_54), .out(tmp02_22_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006945(.in0(tmp01_46_54), .in1(tmp01_47_54), .out(tmp02_23_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006946(.in0(tmp01_48_54), .in1(tmp01_49_54), .out(tmp02_24_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006947(.in0(tmp01_50_54), .in1(tmp01_51_54), .out(tmp02_25_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006948(.in0(tmp01_52_54), .in1(tmp01_53_54), .out(tmp02_26_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006949(.in0(tmp01_54_54), .in1(tmp01_55_54), .out(tmp02_27_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006950(.in0(tmp01_56_54), .in1(tmp01_57_54), .out(tmp02_28_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006951(.in0(tmp01_58_54), .in1(tmp01_59_54), .out(tmp02_29_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006952(.in0(tmp01_60_54), .in1(tmp01_61_54), .out(tmp02_30_54));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add006953(.in0(tmp01_62_54), .in1(tmp01_63_54), .out(tmp02_31_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006954(.in0(tmp02_0_54), .in1(tmp02_1_54), .out(tmp03_0_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006955(.in0(tmp02_2_54), .in1(tmp02_3_54), .out(tmp03_1_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006956(.in0(tmp02_4_54), .in1(tmp02_5_54), .out(tmp03_2_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006957(.in0(tmp02_6_54), .in1(tmp02_7_54), .out(tmp03_3_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006958(.in0(tmp02_8_54), .in1(tmp02_9_54), .out(tmp03_4_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006959(.in0(tmp02_10_54), .in1(tmp02_11_54), .out(tmp03_5_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006960(.in0(tmp02_12_54), .in1(tmp02_13_54), .out(tmp03_6_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006961(.in0(tmp02_14_54), .in1(tmp02_15_54), .out(tmp03_7_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006962(.in0(tmp02_16_54), .in1(tmp02_17_54), .out(tmp03_8_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006963(.in0(tmp02_18_54), .in1(tmp02_19_54), .out(tmp03_9_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006964(.in0(tmp02_20_54), .in1(tmp02_21_54), .out(tmp03_10_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006965(.in0(tmp02_22_54), .in1(tmp02_23_54), .out(tmp03_11_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006966(.in0(tmp02_24_54), .in1(tmp02_25_54), .out(tmp03_12_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006967(.in0(tmp02_26_54), .in1(tmp02_27_54), .out(tmp03_13_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006968(.in0(tmp02_28_54), .in1(tmp02_29_54), .out(tmp03_14_54));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add006969(.in0(tmp02_30_54), .in1(tmp02_31_54), .out(tmp03_15_54));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006970(.in0(tmp03_0_54), .in1(tmp03_1_54), .out(tmp04_0_54));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006971(.in0(tmp03_2_54), .in1(tmp03_3_54), .out(tmp04_1_54));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006972(.in0(tmp03_4_54), .in1(tmp03_5_54), .out(tmp04_2_54));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006973(.in0(tmp03_6_54), .in1(tmp03_7_54), .out(tmp04_3_54));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006974(.in0(tmp03_8_54), .in1(tmp03_9_54), .out(tmp04_4_54));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006975(.in0(tmp03_10_54), .in1(tmp03_11_54), .out(tmp04_5_54));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006976(.in0(tmp03_12_54), .in1(tmp03_13_54), .out(tmp04_6_54));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add006977(.in0(tmp03_14_54), .in1(tmp03_15_54), .out(tmp04_7_54));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006978(.in0(tmp04_0_54), .in1(tmp04_1_54), .out(tmp05_0_54));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006979(.in0(tmp04_2_54), .in1(tmp04_3_54), .out(tmp05_1_54));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006980(.in0(tmp04_4_54), .in1(tmp04_5_54), .out(tmp05_2_54));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add006981(.in0(tmp04_6_54), .in1(tmp04_7_54), .out(tmp05_3_54));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006982(.in0(tmp05_0_54), .in1(tmp05_1_54), .out(tmp06_0_54));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add006983(.in0(tmp05_2_54), .in1(tmp05_3_54), .out(tmp06_1_54));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add006984(.in0(tmp06_0_54), .in1(tmp06_1_54), .out(tmp07_0_54));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006985(.in0(tmp00_0_55), .in1(tmp00_1_55), .out(tmp01_0_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006986(.in0(tmp00_2_55), .in1(tmp00_3_55), .out(tmp01_1_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006987(.in0(tmp00_4_55), .in1(tmp00_5_55), .out(tmp01_2_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006988(.in0(tmp00_6_55), .in1(tmp00_7_55), .out(tmp01_3_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006989(.in0(tmp00_8_55), .in1(tmp00_9_55), .out(tmp01_4_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006990(.in0(tmp00_10_55), .in1(tmp00_11_55), .out(tmp01_5_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006991(.in0(tmp00_12_55), .in1(tmp00_13_55), .out(tmp01_6_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006992(.in0(tmp00_14_55), .in1(tmp00_15_55), .out(tmp01_7_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006993(.in0(tmp00_16_55), .in1(tmp00_17_55), .out(tmp01_8_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006994(.in0(tmp00_18_55), .in1(tmp00_19_55), .out(tmp01_9_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006995(.in0(tmp00_20_55), .in1(tmp00_21_55), .out(tmp01_10_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006996(.in0(tmp00_22_55), .in1(tmp00_23_55), .out(tmp01_11_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006997(.in0(tmp00_24_55), .in1(tmp00_25_55), .out(tmp01_12_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006998(.in0(tmp00_26_55), .in1(tmp00_27_55), .out(tmp01_13_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add006999(.in0(tmp00_28_55), .in1(tmp00_29_55), .out(tmp01_14_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007000(.in0(tmp00_30_55), .in1(tmp00_31_55), .out(tmp01_15_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007001(.in0(tmp00_32_55), .in1(tmp00_33_55), .out(tmp01_16_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007002(.in0(tmp00_34_55), .in1(tmp00_35_55), .out(tmp01_17_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007003(.in0(tmp00_36_55), .in1(tmp00_37_55), .out(tmp01_18_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007004(.in0(tmp00_38_55), .in1(tmp00_39_55), .out(tmp01_19_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007005(.in0(tmp00_40_55), .in1(tmp00_41_55), .out(tmp01_20_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007006(.in0(tmp00_42_55), .in1(tmp00_43_55), .out(tmp01_21_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007007(.in0(tmp00_44_55), .in1(tmp00_45_55), .out(tmp01_22_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007008(.in0(tmp00_46_55), .in1(tmp00_47_55), .out(tmp01_23_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007009(.in0(tmp00_48_55), .in1(tmp00_49_55), .out(tmp01_24_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007010(.in0(tmp00_50_55), .in1(tmp00_51_55), .out(tmp01_25_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007011(.in0(tmp00_52_55), .in1(tmp00_53_55), .out(tmp01_26_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007012(.in0(tmp00_54_55), .in1(tmp00_55_55), .out(tmp01_27_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007013(.in0(tmp00_56_55), .in1(tmp00_57_55), .out(tmp01_28_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007014(.in0(tmp00_58_55), .in1(tmp00_59_55), .out(tmp01_29_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007015(.in0(tmp00_60_55), .in1(tmp00_61_55), .out(tmp01_30_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007016(.in0(tmp00_62_55), .in1(tmp00_63_55), .out(tmp01_31_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007017(.in0(tmp00_64_55), .in1(tmp00_65_55), .out(tmp01_32_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007018(.in0(tmp00_66_55), .in1(tmp00_67_55), .out(tmp01_33_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007019(.in0(tmp00_68_55), .in1(tmp00_69_55), .out(tmp01_34_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007020(.in0(tmp00_70_55), .in1(tmp00_71_55), .out(tmp01_35_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007021(.in0(tmp00_72_55), .in1(tmp00_73_55), .out(tmp01_36_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007022(.in0(tmp00_74_55), .in1(tmp00_75_55), .out(tmp01_37_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007023(.in0(tmp00_76_55), .in1(tmp00_77_55), .out(tmp01_38_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007024(.in0(tmp00_78_55), .in1(tmp00_79_55), .out(tmp01_39_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007025(.in0(tmp00_80_55), .in1(tmp00_81_55), .out(tmp01_40_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007026(.in0(tmp00_82_55), .in1(tmp00_83_55), .out(tmp01_41_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007027(.in0(tmp00_84_55), .in1(tmp00_85_55), .out(tmp01_42_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007028(.in0(tmp00_86_55), .in1(tmp00_87_55), .out(tmp01_43_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007029(.in0(tmp00_88_55), .in1(tmp00_89_55), .out(tmp01_44_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007030(.in0(tmp00_90_55), .in1(tmp00_91_55), .out(tmp01_45_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007031(.in0(tmp00_92_55), .in1(tmp00_93_55), .out(tmp01_46_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007032(.in0(tmp00_94_55), .in1(tmp00_95_55), .out(tmp01_47_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007033(.in0(tmp00_96_55), .in1(tmp00_97_55), .out(tmp01_48_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007034(.in0(tmp00_98_55), .in1(tmp00_99_55), .out(tmp01_49_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007035(.in0(tmp00_100_55), .in1(tmp00_101_55), .out(tmp01_50_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007036(.in0(tmp00_102_55), .in1(tmp00_103_55), .out(tmp01_51_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007037(.in0(tmp00_104_55), .in1(tmp00_105_55), .out(tmp01_52_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007038(.in0(tmp00_106_55), .in1(tmp00_107_55), .out(tmp01_53_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007039(.in0(tmp00_108_55), .in1(tmp00_109_55), .out(tmp01_54_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007040(.in0(tmp00_110_55), .in1(tmp00_111_55), .out(tmp01_55_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007041(.in0(tmp00_112_55), .in1(tmp00_113_55), .out(tmp01_56_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007042(.in0(tmp00_114_55), .in1(tmp00_115_55), .out(tmp01_57_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007043(.in0(tmp00_116_55), .in1(tmp00_117_55), .out(tmp01_58_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007044(.in0(tmp00_118_55), .in1(tmp00_119_55), .out(tmp01_59_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007045(.in0(tmp00_120_55), .in1(tmp00_121_55), .out(tmp01_60_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007046(.in0(tmp00_122_55), .in1(tmp00_123_55), .out(tmp01_61_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007047(.in0(tmp00_124_55), .in1(tmp00_125_55), .out(tmp01_62_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007048(.in0(tmp00_126_55), .in1(tmp00_127_55), .out(tmp01_63_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007049(.in0(tmp01_0_55), .in1(tmp01_1_55), .out(tmp02_0_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007050(.in0(tmp01_2_55), .in1(tmp01_3_55), .out(tmp02_1_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007051(.in0(tmp01_4_55), .in1(tmp01_5_55), .out(tmp02_2_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007052(.in0(tmp01_6_55), .in1(tmp01_7_55), .out(tmp02_3_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007053(.in0(tmp01_8_55), .in1(tmp01_9_55), .out(tmp02_4_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007054(.in0(tmp01_10_55), .in1(tmp01_11_55), .out(tmp02_5_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007055(.in0(tmp01_12_55), .in1(tmp01_13_55), .out(tmp02_6_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007056(.in0(tmp01_14_55), .in1(tmp01_15_55), .out(tmp02_7_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007057(.in0(tmp01_16_55), .in1(tmp01_17_55), .out(tmp02_8_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007058(.in0(tmp01_18_55), .in1(tmp01_19_55), .out(tmp02_9_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007059(.in0(tmp01_20_55), .in1(tmp01_21_55), .out(tmp02_10_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007060(.in0(tmp01_22_55), .in1(tmp01_23_55), .out(tmp02_11_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007061(.in0(tmp01_24_55), .in1(tmp01_25_55), .out(tmp02_12_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007062(.in0(tmp01_26_55), .in1(tmp01_27_55), .out(tmp02_13_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007063(.in0(tmp01_28_55), .in1(tmp01_29_55), .out(tmp02_14_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007064(.in0(tmp01_30_55), .in1(tmp01_31_55), .out(tmp02_15_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007065(.in0(tmp01_32_55), .in1(tmp01_33_55), .out(tmp02_16_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007066(.in0(tmp01_34_55), .in1(tmp01_35_55), .out(tmp02_17_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007067(.in0(tmp01_36_55), .in1(tmp01_37_55), .out(tmp02_18_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007068(.in0(tmp01_38_55), .in1(tmp01_39_55), .out(tmp02_19_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007069(.in0(tmp01_40_55), .in1(tmp01_41_55), .out(tmp02_20_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007070(.in0(tmp01_42_55), .in1(tmp01_43_55), .out(tmp02_21_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007071(.in0(tmp01_44_55), .in1(tmp01_45_55), .out(tmp02_22_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007072(.in0(tmp01_46_55), .in1(tmp01_47_55), .out(tmp02_23_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007073(.in0(tmp01_48_55), .in1(tmp01_49_55), .out(tmp02_24_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007074(.in0(tmp01_50_55), .in1(tmp01_51_55), .out(tmp02_25_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007075(.in0(tmp01_52_55), .in1(tmp01_53_55), .out(tmp02_26_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007076(.in0(tmp01_54_55), .in1(tmp01_55_55), .out(tmp02_27_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007077(.in0(tmp01_56_55), .in1(tmp01_57_55), .out(tmp02_28_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007078(.in0(tmp01_58_55), .in1(tmp01_59_55), .out(tmp02_29_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007079(.in0(tmp01_60_55), .in1(tmp01_61_55), .out(tmp02_30_55));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007080(.in0(tmp01_62_55), .in1(tmp01_63_55), .out(tmp02_31_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007081(.in0(tmp02_0_55), .in1(tmp02_1_55), .out(tmp03_0_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007082(.in0(tmp02_2_55), .in1(tmp02_3_55), .out(tmp03_1_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007083(.in0(tmp02_4_55), .in1(tmp02_5_55), .out(tmp03_2_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007084(.in0(tmp02_6_55), .in1(tmp02_7_55), .out(tmp03_3_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007085(.in0(tmp02_8_55), .in1(tmp02_9_55), .out(tmp03_4_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007086(.in0(tmp02_10_55), .in1(tmp02_11_55), .out(tmp03_5_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007087(.in0(tmp02_12_55), .in1(tmp02_13_55), .out(tmp03_6_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007088(.in0(tmp02_14_55), .in1(tmp02_15_55), .out(tmp03_7_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007089(.in0(tmp02_16_55), .in1(tmp02_17_55), .out(tmp03_8_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007090(.in0(tmp02_18_55), .in1(tmp02_19_55), .out(tmp03_9_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007091(.in0(tmp02_20_55), .in1(tmp02_21_55), .out(tmp03_10_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007092(.in0(tmp02_22_55), .in1(tmp02_23_55), .out(tmp03_11_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007093(.in0(tmp02_24_55), .in1(tmp02_25_55), .out(tmp03_12_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007094(.in0(tmp02_26_55), .in1(tmp02_27_55), .out(tmp03_13_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007095(.in0(tmp02_28_55), .in1(tmp02_29_55), .out(tmp03_14_55));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007096(.in0(tmp02_30_55), .in1(tmp02_31_55), .out(tmp03_15_55));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007097(.in0(tmp03_0_55), .in1(tmp03_1_55), .out(tmp04_0_55));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007098(.in0(tmp03_2_55), .in1(tmp03_3_55), .out(tmp04_1_55));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007099(.in0(tmp03_4_55), .in1(tmp03_5_55), .out(tmp04_2_55));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007100(.in0(tmp03_6_55), .in1(tmp03_7_55), .out(tmp04_3_55));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007101(.in0(tmp03_8_55), .in1(tmp03_9_55), .out(tmp04_4_55));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007102(.in0(tmp03_10_55), .in1(tmp03_11_55), .out(tmp04_5_55));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007103(.in0(tmp03_12_55), .in1(tmp03_13_55), .out(tmp04_6_55));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007104(.in0(tmp03_14_55), .in1(tmp03_15_55), .out(tmp04_7_55));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007105(.in0(tmp04_0_55), .in1(tmp04_1_55), .out(tmp05_0_55));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007106(.in0(tmp04_2_55), .in1(tmp04_3_55), .out(tmp05_1_55));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007107(.in0(tmp04_4_55), .in1(tmp04_5_55), .out(tmp05_2_55));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007108(.in0(tmp04_6_55), .in1(tmp04_7_55), .out(tmp05_3_55));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007109(.in0(tmp05_0_55), .in1(tmp05_1_55), .out(tmp06_0_55));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007110(.in0(tmp05_2_55), .in1(tmp05_3_55), .out(tmp06_1_55));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add007111(.in0(tmp06_0_55), .in1(tmp06_1_55), .out(tmp07_0_55));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007112(.in0(tmp00_0_56), .in1(tmp00_1_56), .out(tmp01_0_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007113(.in0(tmp00_2_56), .in1(tmp00_3_56), .out(tmp01_1_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007114(.in0(tmp00_4_56), .in1(tmp00_5_56), .out(tmp01_2_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007115(.in0(tmp00_6_56), .in1(tmp00_7_56), .out(tmp01_3_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007116(.in0(tmp00_8_56), .in1(tmp00_9_56), .out(tmp01_4_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007117(.in0(tmp00_10_56), .in1(tmp00_11_56), .out(tmp01_5_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007118(.in0(tmp00_12_56), .in1(tmp00_13_56), .out(tmp01_6_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007119(.in0(tmp00_14_56), .in1(tmp00_15_56), .out(tmp01_7_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007120(.in0(tmp00_16_56), .in1(tmp00_17_56), .out(tmp01_8_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007121(.in0(tmp00_18_56), .in1(tmp00_19_56), .out(tmp01_9_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007122(.in0(tmp00_20_56), .in1(tmp00_21_56), .out(tmp01_10_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007123(.in0(tmp00_22_56), .in1(tmp00_23_56), .out(tmp01_11_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007124(.in0(tmp00_24_56), .in1(tmp00_25_56), .out(tmp01_12_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007125(.in0(tmp00_26_56), .in1(tmp00_27_56), .out(tmp01_13_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007126(.in0(tmp00_28_56), .in1(tmp00_29_56), .out(tmp01_14_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007127(.in0(tmp00_30_56), .in1(tmp00_31_56), .out(tmp01_15_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007128(.in0(tmp00_32_56), .in1(tmp00_33_56), .out(tmp01_16_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007129(.in0(tmp00_34_56), .in1(tmp00_35_56), .out(tmp01_17_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007130(.in0(tmp00_36_56), .in1(tmp00_37_56), .out(tmp01_18_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007131(.in0(tmp00_38_56), .in1(tmp00_39_56), .out(tmp01_19_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007132(.in0(tmp00_40_56), .in1(tmp00_41_56), .out(tmp01_20_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007133(.in0(tmp00_42_56), .in1(tmp00_43_56), .out(tmp01_21_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007134(.in0(tmp00_44_56), .in1(tmp00_45_56), .out(tmp01_22_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007135(.in0(tmp00_46_56), .in1(tmp00_47_56), .out(tmp01_23_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007136(.in0(tmp00_48_56), .in1(tmp00_49_56), .out(tmp01_24_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007137(.in0(tmp00_50_56), .in1(tmp00_51_56), .out(tmp01_25_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007138(.in0(tmp00_52_56), .in1(tmp00_53_56), .out(tmp01_26_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007139(.in0(tmp00_54_56), .in1(tmp00_55_56), .out(tmp01_27_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007140(.in0(tmp00_56_56), .in1(tmp00_57_56), .out(tmp01_28_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007141(.in0(tmp00_58_56), .in1(tmp00_59_56), .out(tmp01_29_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007142(.in0(tmp00_60_56), .in1(tmp00_61_56), .out(tmp01_30_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007143(.in0(tmp00_62_56), .in1(tmp00_63_56), .out(tmp01_31_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007144(.in0(tmp00_64_56), .in1(tmp00_65_56), .out(tmp01_32_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007145(.in0(tmp00_66_56), .in1(tmp00_67_56), .out(tmp01_33_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007146(.in0(tmp00_68_56), .in1(tmp00_69_56), .out(tmp01_34_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007147(.in0(tmp00_70_56), .in1(tmp00_71_56), .out(tmp01_35_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007148(.in0(tmp00_72_56), .in1(tmp00_73_56), .out(tmp01_36_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007149(.in0(tmp00_74_56), .in1(tmp00_75_56), .out(tmp01_37_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007150(.in0(tmp00_76_56), .in1(tmp00_77_56), .out(tmp01_38_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007151(.in0(tmp00_78_56), .in1(tmp00_79_56), .out(tmp01_39_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007152(.in0(tmp00_80_56), .in1(tmp00_81_56), .out(tmp01_40_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007153(.in0(tmp00_82_56), .in1(tmp00_83_56), .out(tmp01_41_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007154(.in0(tmp00_84_56), .in1(tmp00_85_56), .out(tmp01_42_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007155(.in0(tmp00_86_56), .in1(tmp00_87_56), .out(tmp01_43_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007156(.in0(tmp00_88_56), .in1(tmp00_89_56), .out(tmp01_44_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007157(.in0(tmp00_90_56), .in1(tmp00_91_56), .out(tmp01_45_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007158(.in0(tmp00_92_56), .in1(tmp00_93_56), .out(tmp01_46_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007159(.in0(tmp00_94_56), .in1(tmp00_95_56), .out(tmp01_47_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007160(.in0(tmp00_96_56), .in1(tmp00_97_56), .out(tmp01_48_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007161(.in0(tmp00_98_56), .in1(tmp00_99_56), .out(tmp01_49_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007162(.in0(tmp00_100_56), .in1(tmp00_101_56), .out(tmp01_50_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007163(.in0(tmp00_102_56), .in1(tmp00_103_56), .out(tmp01_51_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007164(.in0(tmp00_104_56), .in1(tmp00_105_56), .out(tmp01_52_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007165(.in0(tmp00_106_56), .in1(tmp00_107_56), .out(tmp01_53_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007166(.in0(tmp00_108_56), .in1(tmp00_109_56), .out(tmp01_54_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007167(.in0(tmp00_110_56), .in1(tmp00_111_56), .out(tmp01_55_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007168(.in0(tmp00_112_56), .in1(tmp00_113_56), .out(tmp01_56_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007169(.in0(tmp00_114_56), .in1(tmp00_115_56), .out(tmp01_57_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007170(.in0(tmp00_116_56), .in1(tmp00_117_56), .out(tmp01_58_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007171(.in0(tmp00_118_56), .in1(tmp00_119_56), .out(tmp01_59_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007172(.in0(tmp00_120_56), .in1(tmp00_121_56), .out(tmp01_60_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007173(.in0(tmp00_122_56), .in1(tmp00_123_56), .out(tmp01_61_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007174(.in0(tmp00_124_56), .in1(tmp00_125_56), .out(tmp01_62_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007175(.in0(tmp00_126_56), .in1(tmp00_127_56), .out(tmp01_63_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007176(.in0(tmp01_0_56), .in1(tmp01_1_56), .out(tmp02_0_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007177(.in0(tmp01_2_56), .in1(tmp01_3_56), .out(tmp02_1_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007178(.in0(tmp01_4_56), .in1(tmp01_5_56), .out(tmp02_2_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007179(.in0(tmp01_6_56), .in1(tmp01_7_56), .out(tmp02_3_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007180(.in0(tmp01_8_56), .in1(tmp01_9_56), .out(tmp02_4_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007181(.in0(tmp01_10_56), .in1(tmp01_11_56), .out(tmp02_5_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007182(.in0(tmp01_12_56), .in1(tmp01_13_56), .out(tmp02_6_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007183(.in0(tmp01_14_56), .in1(tmp01_15_56), .out(tmp02_7_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007184(.in0(tmp01_16_56), .in1(tmp01_17_56), .out(tmp02_8_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007185(.in0(tmp01_18_56), .in1(tmp01_19_56), .out(tmp02_9_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007186(.in0(tmp01_20_56), .in1(tmp01_21_56), .out(tmp02_10_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007187(.in0(tmp01_22_56), .in1(tmp01_23_56), .out(tmp02_11_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007188(.in0(tmp01_24_56), .in1(tmp01_25_56), .out(tmp02_12_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007189(.in0(tmp01_26_56), .in1(tmp01_27_56), .out(tmp02_13_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007190(.in0(tmp01_28_56), .in1(tmp01_29_56), .out(tmp02_14_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007191(.in0(tmp01_30_56), .in1(tmp01_31_56), .out(tmp02_15_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007192(.in0(tmp01_32_56), .in1(tmp01_33_56), .out(tmp02_16_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007193(.in0(tmp01_34_56), .in1(tmp01_35_56), .out(tmp02_17_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007194(.in0(tmp01_36_56), .in1(tmp01_37_56), .out(tmp02_18_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007195(.in0(tmp01_38_56), .in1(tmp01_39_56), .out(tmp02_19_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007196(.in0(tmp01_40_56), .in1(tmp01_41_56), .out(tmp02_20_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007197(.in0(tmp01_42_56), .in1(tmp01_43_56), .out(tmp02_21_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007198(.in0(tmp01_44_56), .in1(tmp01_45_56), .out(tmp02_22_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007199(.in0(tmp01_46_56), .in1(tmp01_47_56), .out(tmp02_23_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007200(.in0(tmp01_48_56), .in1(tmp01_49_56), .out(tmp02_24_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007201(.in0(tmp01_50_56), .in1(tmp01_51_56), .out(tmp02_25_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007202(.in0(tmp01_52_56), .in1(tmp01_53_56), .out(tmp02_26_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007203(.in0(tmp01_54_56), .in1(tmp01_55_56), .out(tmp02_27_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007204(.in0(tmp01_56_56), .in1(tmp01_57_56), .out(tmp02_28_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007205(.in0(tmp01_58_56), .in1(tmp01_59_56), .out(tmp02_29_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007206(.in0(tmp01_60_56), .in1(tmp01_61_56), .out(tmp02_30_56));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007207(.in0(tmp01_62_56), .in1(tmp01_63_56), .out(tmp02_31_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007208(.in0(tmp02_0_56), .in1(tmp02_1_56), .out(tmp03_0_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007209(.in0(tmp02_2_56), .in1(tmp02_3_56), .out(tmp03_1_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007210(.in0(tmp02_4_56), .in1(tmp02_5_56), .out(tmp03_2_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007211(.in0(tmp02_6_56), .in1(tmp02_7_56), .out(tmp03_3_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007212(.in0(tmp02_8_56), .in1(tmp02_9_56), .out(tmp03_4_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007213(.in0(tmp02_10_56), .in1(tmp02_11_56), .out(tmp03_5_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007214(.in0(tmp02_12_56), .in1(tmp02_13_56), .out(tmp03_6_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007215(.in0(tmp02_14_56), .in1(tmp02_15_56), .out(tmp03_7_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007216(.in0(tmp02_16_56), .in1(tmp02_17_56), .out(tmp03_8_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007217(.in0(tmp02_18_56), .in1(tmp02_19_56), .out(tmp03_9_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007218(.in0(tmp02_20_56), .in1(tmp02_21_56), .out(tmp03_10_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007219(.in0(tmp02_22_56), .in1(tmp02_23_56), .out(tmp03_11_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007220(.in0(tmp02_24_56), .in1(tmp02_25_56), .out(tmp03_12_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007221(.in0(tmp02_26_56), .in1(tmp02_27_56), .out(tmp03_13_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007222(.in0(tmp02_28_56), .in1(tmp02_29_56), .out(tmp03_14_56));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007223(.in0(tmp02_30_56), .in1(tmp02_31_56), .out(tmp03_15_56));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007224(.in0(tmp03_0_56), .in1(tmp03_1_56), .out(tmp04_0_56));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007225(.in0(tmp03_2_56), .in1(tmp03_3_56), .out(tmp04_1_56));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007226(.in0(tmp03_4_56), .in1(tmp03_5_56), .out(tmp04_2_56));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007227(.in0(tmp03_6_56), .in1(tmp03_7_56), .out(tmp04_3_56));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007228(.in0(tmp03_8_56), .in1(tmp03_9_56), .out(tmp04_4_56));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007229(.in0(tmp03_10_56), .in1(tmp03_11_56), .out(tmp04_5_56));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007230(.in0(tmp03_12_56), .in1(tmp03_13_56), .out(tmp04_6_56));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007231(.in0(tmp03_14_56), .in1(tmp03_15_56), .out(tmp04_7_56));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007232(.in0(tmp04_0_56), .in1(tmp04_1_56), .out(tmp05_0_56));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007233(.in0(tmp04_2_56), .in1(tmp04_3_56), .out(tmp05_1_56));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007234(.in0(tmp04_4_56), .in1(tmp04_5_56), .out(tmp05_2_56));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007235(.in0(tmp04_6_56), .in1(tmp04_7_56), .out(tmp05_3_56));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007236(.in0(tmp05_0_56), .in1(tmp05_1_56), .out(tmp06_0_56));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007237(.in0(tmp05_2_56), .in1(tmp05_3_56), .out(tmp06_1_56));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add007238(.in0(tmp06_0_56), .in1(tmp06_1_56), .out(tmp07_0_56));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007239(.in0(tmp00_0_57), .in1(tmp00_1_57), .out(tmp01_0_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007240(.in0(tmp00_2_57), .in1(tmp00_3_57), .out(tmp01_1_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007241(.in0(tmp00_4_57), .in1(tmp00_5_57), .out(tmp01_2_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007242(.in0(tmp00_6_57), .in1(tmp00_7_57), .out(tmp01_3_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007243(.in0(tmp00_8_57), .in1(tmp00_9_57), .out(tmp01_4_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007244(.in0(tmp00_10_57), .in1(tmp00_11_57), .out(tmp01_5_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007245(.in0(tmp00_12_57), .in1(tmp00_13_57), .out(tmp01_6_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007246(.in0(tmp00_14_57), .in1(tmp00_15_57), .out(tmp01_7_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007247(.in0(tmp00_16_57), .in1(tmp00_17_57), .out(tmp01_8_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007248(.in0(tmp00_18_57), .in1(tmp00_19_57), .out(tmp01_9_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007249(.in0(tmp00_20_57), .in1(tmp00_21_57), .out(tmp01_10_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007250(.in0(tmp00_22_57), .in1(tmp00_23_57), .out(tmp01_11_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007251(.in0(tmp00_24_57), .in1(tmp00_25_57), .out(tmp01_12_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007252(.in0(tmp00_26_57), .in1(tmp00_27_57), .out(tmp01_13_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007253(.in0(tmp00_28_57), .in1(tmp00_29_57), .out(tmp01_14_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007254(.in0(tmp00_30_57), .in1(tmp00_31_57), .out(tmp01_15_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007255(.in0(tmp00_32_57), .in1(tmp00_33_57), .out(tmp01_16_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007256(.in0(tmp00_34_57), .in1(tmp00_35_57), .out(tmp01_17_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007257(.in0(tmp00_36_57), .in1(tmp00_37_57), .out(tmp01_18_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007258(.in0(tmp00_38_57), .in1(tmp00_39_57), .out(tmp01_19_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007259(.in0(tmp00_40_57), .in1(tmp00_41_57), .out(tmp01_20_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007260(.in0(tmp00_42_57), .in1(tmp00_43_57), .out(tmp01_21_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007261(.in0(tmp00_44_57), .in1(tmp00_45_57), .out(tmp01_22_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007262(.in0(tmp00_46_57), .in1(tmp00_47_57), .out(tmp01_23_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007263(.in0(tmp00_48_57), .in1(tmp00_49_57), .out(tmp01_24_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007264(.in0(tmp00_50_57), .in1(tmp00_51_57), .out(tmp01_25_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007265(.in0(tmp00_52_57), .in1(tmp00_53_57), .out(tmp01_26_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007266(.in0(tmp00_54_57), .in1(tmp00_55_57), .out(tmp01_27_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007267(.in0(tmp00_56_57), .in1(tmp00_57_57), .out(tmp01_28_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007268(.in0(tmp00_58_57), .in1(tmp00_59_57), .out(tmp01_29_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007269(.in0(tmp00_60_57), .in1(tmp00_61_57), .out(tmp01_30_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007270(.in0(tmp00_62_57), .in1(tmp00_63_57), .out(tmp01_31_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007271(.in0(tmp00_64_57), .in1(tmp00_65_57), .out(tmp01_32_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007272(.in0(tmp00_66_57), .in1(tmp00_67_57), .out(tmp01_33_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007273(.in0(tmp00_68_57), .in1(tmp00_69_57), .out(tmp01_34_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007274(.in0(tmp00_70_57), .in1(tmp00_71_57), .out(tmp01_35_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007275(.in0(tmp00_72_57), .in1(tmp00_73_57), .out(tmp01_36_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007276(.in0(tmp00_74_57), .in1(tmp00_75_57), .out(tmp01_37_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007277(.in0(tmp00_76_57), .in1(tmp00_77_57), .out(tmp01_38_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007278(.in0(tmp00_78_57), .in1(tmp00_79_57), .out(tmp01_39_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007279(.in0(tmp00_80_57), .in1(tmp00_81_57), .out(tmp01_40_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007280(.in0(tmp00_82_57), .in1(tmp00_83_57), .out(tmp01_41_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007281(.in0(tmp00_84_57), .in1(tmp00_85_57), .out(tmp01_42_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007282(.in0(tmp00_86_57), .in1(tmp00_87_57), .out(tmp01_43_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007283(.in0(tmp00_88_57), .in1(tmp00_89_57), .out(tmp01_44_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007284(.in0(tmp00_90_57), .in1(tmp00_91_57), .out(tmp01_45_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007285(.in0(tmp00_92_57), .in1(tmp00_93_57), .out(tmp01_46_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007286(.in0(tmp00_94_57), .in1(tmp00_95_57), .out(tmp01_47_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007287(.in0(tmp00_96_57), .in1(tmp00_97_57), .out(tmp01_48_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007288(.in0(tmp00_98_57), .in1(tmp00_99_57), .out(tmp01_49_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007289(.in0(tmp00_100_57), .in1(tmp00_101_57), .out(tmp01_50_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007290(.in0(tmp00_102_57), .in1(tmp00_103_57), .out(tmp01_51_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007291(.in0(tmp00_104_57), .in1(tmp00_105_57), .out(tmp01_52_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007292(.in0(tmp00_106_57), .in1(tmp00_107_57), .out(tmp01_53_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007293(.in0(tmp00_108_57), .in1(tmp00_109_57), .out(tmp01_54_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007294(.in0(tmp00_110_57), .in1(tmp00_111_57), .out(tmp01_55_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007295(.in0(tmp00_112_57), .in1(tmp00_113_57), .out(tmp01_56_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007296(.in0(tmp00_114_57), .in1(tmp00_115_57), .out(tmp01_57_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007297(.in0(tmp00_116_57), .in1(tmp00_117_57), .out(tmp01_58_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007298(.in0(tmp00_118_57), .in1(tmp00_119_57), .out(tmp01_59_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007299(.in0(tmp00_120_57), .in1(tmp00_121_57), .out(tmp01_60_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007300(.in0(tmp00_122_57), .in1(tmp00_123_57), .out(tmp01_61_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007301(.in0(tmp00_124_57), .in1(tmp00_125_57), .out(tmp01_62_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007302(.in0(tmp00_126_57), .in1(tmp00_127_57), .out(tmp01_63_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007303(.in0(tmp01_0_57), .in1(tmp01_1_57), .out(tmp02_0_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007304(.in0(tmp01_2_57), .in1(tmp01_3_57), .out(tmp02_1_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007305(.in0(tmp01_4_57), .in1(tmp01_5_57), .out(tmp02_2_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007306(.in0(tmp01_6_57), .in1(tmp01_7_57), .out(tmp02_3_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007307(.in0(tmp01_8_57), .in1(tmp01_9_57), .out(tmp02_4_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007308(.in0(tmp01_10_57), .in1(tmp01_11_57), .out(tmp02_5_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007309(.in0(tmp01_12_57), .in1(tmp01_13_57), .out(tmp02_6_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007310(.in0(tmp01_14_57), .in1(tmp01_15_57), .out(tmp02_7_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007311(.in0(tmp01_16_57), .in1(tmp01_17_57), .out(tmp02_8_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007312(.in0(tmp01_18_57), .in1(tmp01_19_57), .out(tmp02_9_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007313(.in0(tmp01_20_57), .in1(tmp01_21_57), .out(tmp02_10_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007314(.in0(tmp01_22_57), .in1(tmp01_23_57), .out(tmp02_11_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007315(.in0(tmp01_24_57), .in1(tmp01_25_57), .out(tmp02_12_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007316(.in0(tmp01_26_57), .in1(tmp01_27_57), .out(tmp02_13_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007317(.in0(tmp01_28_57), .in1(tmp01_29_57), .out(tmp02_14_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007318(.in0(tmp01_30_57), .in1(tmp01_31_57), .out(tmp02_15_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007319(.in0(tmp01_32_57), .in1(tmp01_33_57), .out(tmp02_16_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007320(.in0(tmp01_34_57), .in1(tmp01_35_57), .out(tmp02_17_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007321(.in0(tmp01_36_57), .in1(tmp01_37_57), .out(tmp02_18_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007322(.in0(tmp01_38_57), .in1(tmp01_39_57), .out(tmp02_19_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007323(.in0(tmp01_40_57), .in1(tmp01_41_57), .out(tmp02_20_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007324(.in0(tmp01_42_57), .in1(tmp01_43_57), .out(tmp02_21_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007325(.in0(tmp01_44_57), .in1(tmp01_45_57), .out(tmp02_22_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007326(.in0(tmp01_46_57), .in1(tmp01_47_57), .out(tmp02_23_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007327(.in0(tmp01_48_57), .in1(tmp01_49_57), .out(tmp02_24_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007328(.in0(tmp01_50_57), .in1(tmp01_51_57), .out(tmp02_25_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007329(.in0(tmp01_52_57), .in1(tmp01_53_57), .out(tmp02_26_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007330(.in0(tmp01_54_57), .in1(tmp01_55_57), .out(tmp02_27_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007331(.in0(tmp01_56_57), .in1(tmp01_57_57), .out(tmp02_28_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007332(.in0(tmp01_58_57), .in1(tmp01_59_57), .out(tmp02_29_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007333(.in0(tmp01_60_57), .in1(tmp01_61_57), .out(tmp02_30_57));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007334(.in0(tmp01_62_57), .in1(tmp01_63_57), .out(tmp02_31_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007335(.in0(tmp02_0_57), .in1(tmp02_1_57), .out(tmp03_0_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007336(.in0(tmp02_2_57), .in1(tmp02_3_57), .out(tmp03_1_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007337(.in0(tmp02_4_57), .in1(tmp02_5_57), .out(tmp03_2_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007338(.in0(tmp02_6_57), .in1(tmp02_7_57), .out(tmp03_3_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007339(.in0(tmp02_8_57), .in1(tmp02_9_57), .out(tmp03_4_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007340(.in0(tmp02_10_57), .in1(tmp02_11_57), .out(tmp03_5_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007341(.in0(tmp02_12_57), .in1(tmp02_13_57), .out(tmp03_6_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007342(.in0(tmp02_14_57), .in1(tmp02_15_57), .out(tmp03_7_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007343(.in0(tmp02_16_57), .in1(tmp02_17_57), .out(tmp03_8_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007344(.in0(tmp02_18_57), .in1(tmp02_19_57), .out(tmp03_9_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007345(.in0(tmp02_20_57), .in1(tmp02_21_57), .out(tmp03_10_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007346(.in0(tmp02_22_57), .in1(tmp02_23_57), .out(tmp03_11_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007347(.in0(tmp02_24_57), .in1(tmp02_25_57), .out(tmp03_12_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007348(.in0(tmp02_26_57), .in1(tmp02_27_57), .out(tmp03_13_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007349(.in0(tmp02_28_57), .in1(tmp02_29_57), .out(tmp03_14_57));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007350(.in0(tmp02_30_57), .in1(tmp02_31_57), .out(tmp03_15_57));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007351(.in0(tmp03_0_57), .in1(tmp03_1_57), .out(tmp04_0_57));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007352(.in0(tmp03_2_57), .in1(tmp03_3_57), .out(tmp04_1_57));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007353(.in0(tmp03_4_57), .in1(tmp03_5_57), .out(tmp04_2_57));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007354(.in0(tmp03_6_57), .in1(tmp03_7_57), .out(tmp04_3_57));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007355(.in0(tmp03_8_57), .in1(tmp03_9_57), .out(tmp04_4_57));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007356(.in0(tmp03_10_57), .in1(tmp03_11_57), .out(tmp04_5_57));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007357(.in0(tmp03_12_57), .in1(tmp03_13_57), .out(tmp04_6_57));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007358(.in0(tmp03_14_57), .in1(tmp03_15_57), .out(tmp04_7_57));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007359(.in0(tmp04_0_57), .in1(tmp04_1_57), .out(tmp05_0_57));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007360(.in0(tmp04_2_57), .in1(tmp04_3_57), .out(tmp05_1_57));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007361(.in0(tmp04_4_57), .in1(tmp04_5_57), .out(tmp05_2_57));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007362(.in0(tmp04_6_57), .in1(tmp04_7_57), .out(tmp05_3_57));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007363(.in0(tmp05_0_57), .in1(tmp05_1_57), .out(tmp06_0_57));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007364(.in0(tmp05_2_57), .in1(tmp05_3_57), .out(tmp06_1_57));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add007365(.in0(tmp06_0_57), .in1(tmp06_1_57), .out(tmp07_0_57));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007366(.in0(tmp00_0_58), .in1(tmp00_1_58), .out(tmp01_0_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007367(.in0(tmp00_2_58), .in1(tmp00_3_58), .out(tmp01_1_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007368(.in0(tmp00_4_58), .in1(tmp00_5_58), .out(tmp01_2_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007369(.in0(tmp00_6_58), .in1(tmp00_7_58), .out(tmp01_3_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007370(.in0(tmp00_8_58), .in1(tmp00_9_58), .out(tmp01_4_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007371(.in0(tmp00_10_58), .in1(tmp00_11_58), .out(tmp01_5_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007372(.in0(tmp00_12_58), .in1(tmp00_13_58), .out(tmp01_6_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007373(.in0(tmp00_14_58), .in1(tmp00_15_58), .out(tmp01_7_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007374(.in0(tmp00_16_58), .in1(tmp00_17_58), .out(tmp01_8_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007375(.in0(tmp00_18_58), .in1(tmp00_19_58), .out(tmp01_9_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007376(.in0(tmp00_20_58), .in1(tmp00_21_58), .out(tmp01_10_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007377(.in0(tmp00_22_58), .in1(tmp00_23_58), .out(tmp01_11_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007378(.in0(tmp00_24_58), .in1(tmp00_25_58), .out(tmp01_12_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007379(.in0(tmp00_26_58), .in1(tmp00_27_58), .out(tmp01_13_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007380(.in0(tmp00_28_58), .in1(tmp00_29_58), .out(tmp01_14_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007381(.in0(tmp00_30_58), .in1(tmp00_31_58), .out(tmp01_15_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007382(.in0(tmp00_32_58), .in1(tmp00_33_58), .out(tmp01_16_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007383(.in0(tmp00_34_58), .in1(tmp00_35_58), .out(tmp01_17_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007384(.in0(tmp00_36_58), .in1(tmp00_37_58), .out(tmp01_18_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007385(.in0(tmp00_38_58), .in1(tmp00_39_58), .out(tmp01_19_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007386(.in0(tmp00_40_58), .in1(tmp00_41_58), .out(tmp01_20_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007387(.in0(tmp00_42_58), .in1(tmp00_43_58), .out(tmp01_21_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007388(.in0(tmp00_44_58), .in1(tmp00_45_58), .out(tmp01_22_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007389(.in0(tmp00_46_58), .in1(tmp00_47_58), .out(tmp01_23_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007390(.in0(tmp00_48_58), .in1(tmp00_49_58), .out(tmp01_24_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007391(.in0(tmp00_50_58), .in1(tmp00_51_58), .out(tmp01_25_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007392(.in0(tmp00_52_58), .in1(tmp00_53_58), .out(tmp01_26_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007393(.in0(tmp00_54_58), .in1(tmp00_55_58), .out(tmp01_27_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007394(.in0(tmp00_56_58), .in1(tmp00_57_58), .out(tmp01_28_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007395(.in0(tmp00_58_58), .in1(tmp00_59_58), .out(tmp01_29_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007396(.in0(tmp00_60_58), .in1(tmp00_61_58), .out(tmp01_30_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007397(.in0(tmp00_62_58), .in1(tmp00_63_58), .out(tmp01_31_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007398(.in0(tmp00_64_58), .in1(tmp00_65_58), .out(tmp01_32_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007399(.in0(tmp00_66_58), .in1(tmp00_67_58), .out(tmp01_33_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007400(.in0(tmp00_68_58), .in1(tmp00_69_58), .out(tmp01_34_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007401(.in0(tmp00_70_58), .in1(tmp00_71_58), .out(tmp01_35_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007402(.in0(tmp00_72_58), .in1(tmp00_73_58), .out(tmp01_36_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007403(.in0(tmp00_74_58), .in1(tmp00_75_58), .out(tmp01_37_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007404(.in0(tmp00_76_58), .in1(tmp00_77_58), .out(tmp01_38_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007405(.in0(tmp00_78_58), .in1(tmp00_79_58), .out(tmp01_39_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007406(.in0(tmp00_80_58), .in1(tmp00_81_58), .out(tmp01_40_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007407(.in0(tmp00_82_58), .in1(tmp00_83_58), .out(tmp01_41_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007408(.in0(tmp00_84_58), .in1(tmp00_85_58), .out(tmp01_42_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007409(.in0(tmp00_86_58), .in1(tmp00_87_58), .out(tmp01_43_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007410(.in0(tmp00_88_58), .in1(tmp00_89_58), .out(tmp01_44_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007411(.in0(tmp00_90_58), .in1(tmp00_91_58), .out(tmp01_45_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007412(.in0(tmp00_92_58), .in1(tmp00_93_58), .out(tmp01_46_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007413(.in0(tmp00_94_58), .in1(tmp00_95_58), .out(tmp01_47_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007414(.in0(tmp00_96_58), .in1(tmp00_97_58), .out(tmp01_48_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007415(.in0(tmp00_98_58), .in1(tmp00_99_58), .out(tmp01_49_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007416(.in0(tmp00_100_58), .in1(tmp00_101_58), .out(tmp01_50_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007417(.in0(tmp00_102_58), .in1(tmp00_103_58), .out(tmp01_51_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007418(.in0(tmp00_104_58), .in1(tmp00_105_58), .out(tmp01_52_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007419(.in0(tmp00_106_58), .in1(tmp00_107_58), .out(tmp01_53_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007420(.in0(tmp00_108_58), .in1(tmp00_109_58), .out(tmp01_54_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007421(.in0(tmp00_110_58), .in1(tmp00_111_58), .out(tmp01_55_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007422(.in0(tmp00_112_58), .in1(tmp00_113_58), .out(tmp01_56_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007423(.in0(tmp00_114_58), .in1(tmp00_115_58), .out(tmp01_57_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007424(.in0(tmp00_116_58), .in1(tmp00_117_58), .out(tmp01_58_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007425(.in0(tmp00_118_58), .in1(tmp00_119_58), .out(tmp01_59_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007426(.in0(tmp00_120_58), .in1(tmp00_121_58), .out(tmp01_60_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007427(.in0(tmp00_122_58), .in1(tmp00_123_58), .out(tmp01_61_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007428(.in0(tmp00_124_58), .in1(tmp00_125_58), .out(tmp01_62_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007429(.in0(tmp00_126_58), .in1(tmp00_127_58), .out(tmp01_63_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007430(.in0(tmp01_0_58), .in1(tmp01_1_58), .out(tmp02_0_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007431(.in0(tmp01_2_58), .in1(tmp01_3_58), .out(tmp02_1_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007432(.in0(tmp01_4_58), .in1(tmp01_5_58), .out(tmp02_2_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007433(.in0(tmp01_6_58), .in1(tmp01_7_58), .out(tmp02_3_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007434(.in0(tmp01_8_58), .in1(tmp01_9_58), .out(tmp02_4_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007435(.in0(tmp01_10_58), .in1(tmp01_11_58), .out(tmp02_5_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007436(.in0(tmp01_12_58), .in1(tmp01_13_58), .out(tmp02_6_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007437(.in0(tmp01_14_58), .in1(tmp01_15_58), .out(tmp02_7_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007438(.in0(tmp01_16_58), .in1(tmp01_17_58), .out(tmp02_8_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007439(.in0(tmp01_18_58), .in1(tmp01_19_58), .out(tmp02_9_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007440(.in0(tmp01_20_58), .in1(tmp01_21_58), .out(tmp02_10_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007441(.in0(tmp01_22_58), .in1(tmp01_23_58), .out(tmp02_11_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007442(.in0(tmp01_24_58), .in1(tmp01_25_58), .out(tmp02_12_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007443(.in0(tmp01_26_58), .in1(tmp01_27_58), .out(tmp02_13_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007444(.in0(tmp01_28_58), .in1(tmp01_29_58), .out(tmp02_14_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007445(.in0(tmp01_30_58), .in1(tmp01_31_58), .out(tmp02_15_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007446(.in0(tmp01_32_58), .in1(tmp01_33_58), .out(tmp02_16_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007447(.in0(tmp01_34_58), .in1(tmp01_35_58), .out(tmp02_17_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007448(.in0(tmp01_36_58), .in1(tmp01_37_58), .out(tmp02_18_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007449(.in0(tmp01_38_58), .in1(tmp01_39_58), .out(tmp02_19_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007450(.in0(tmp01_40_58), .in1(tmp01_41_58), .out(tmp02_20_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007451(.in0(tmp01_42_58), .in1(tmp01_43_58), .out(tmp02_21_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007452(.in0(tmp01_44_58), .in1(tmp01_45_58), .out(tmp02_22_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007453(.in0(tmp01_46_58), .in1(tmp01_47_58), .out(tmp02_23_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007454(.in0(tmp01_48_58), .in1(tmp01_49_58), .out(tmp02_24_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007455(.in0(tmp01_50_58), .in1(tmp01_51_58), .out(tmp02_25_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007456(.in0(tmp01_52_58), .in1(tmp01_53_58), .out(tmp02_26_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007457(.in0(tmp01_54_58), .in1(tmp01_55_58), .out(tmp02_27_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007458(.in0(tmp01_56_58), .in1(tmp01_57_58), .out(tmp02_28_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007459(.in0(tmp01_58_58), .in1(tmp01_59_58), .out(tmp02_29_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007460(.in0(tmp01_60_58), .in1(tmp01_61_58), .out(tmp02_30_58));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007461(.in0(tmp01_62_58), .in1(tmp01_63_58), .out(tmp02_31_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007462(.in0(tmp02_0_58), .in1(tmp02_1_58), .out(tmp03_0_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007463(.in0(tmp02_2_58), .in1(tmp02_3_58), .out(tmp03_1_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007464(.in0(tmp02_4_58), .in1(tmp02_5_58), .out(tmp03_2_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007465(.in0(tmp02_6_58), .in1(tmp02_7_58), .out(tmp03_3_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007466(.in0(tmp02_8_58), .in1(tmp02_9_58), .out(tmp03_4_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007467(.in0(tmp02_10_58), .in1(tmp02_11_58), .out(tmp03_5_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007468(.in0(tmp02_12_58), .in1(tmp02_13_58), .out(tmp03_6_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007469(.in0(tmp02_14_58), .in1(tmp02_15_58), .out(tmp03_7_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007470(.in0(tmp02_16_58), .in1(tmp02_17_58), .out(tmp03_8_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007471(.in0(tmp02_18_58), .in1(tmp02_19_58), .out(tmp03_9_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007472(.in0(tmp02_20_58), .in1(tmp02_21_58), .out(tmp03_10_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007473(.in0(tmp02_22_58), .in1(tmp02_23_58), .out(tmp03_11_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007474(.in0(tmp02_24_58), .in1(tmp02_25_58), .out(tmp03_12_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007475(.in0(tmp02_26_58), .in1(tmp02_27_58), .out(tmp03_13_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007476(.in0(tmp02_28_58), .in1(tmp02_29_58), .out(tmp03_14_58));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007477(.in0(tmp02_30_58), .in1(tmp02_31_58), .out(tmp03_15_58));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007478(.in0(tmp03_0_58), .in1(tmp03_1_58), .out(tmp04_0_58));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007479(.in0(tmp03_2_58), .in1(tmp03_3_58), .out(tmp04_1_58));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007480(.in0(tmp03_4_58), .in1(tmp03_5_58), .out(tmp04_2_58));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007481(.in0(tmp03_6_58), .in1(tmp03_7_58), .out(tmp04_3_58));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007482(.in0(tmp03_8_58), .in1(tmp03_9_58), .out(tmp04_4_58));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007483(.in0(tmp03_10_58), .in1(tmp03_11_58), .out(tmp04_5_58));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007484(.in0(tmp03_12_58), .in1(tmp03_13_58), .out(tmp04_6_58));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007485(.in0(tmp03_14_58), .in1(tmp03_15_58), .out(tmp04_7_58));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007486(.in0(tmp04_0_58), .in1(tmp04_1_58), .out(tmp05_0_58));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007487(.in0(tmp04_2_58), .in1(tmp04_3_58), .out(tmp05_1_58));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007488(.in0(tmp04_4_58), .in1(tmp04_5_58), .out(tmp05_2_58));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007489(.in0(tmp04_6_58), .in1(tmp04_7_58), .out(tmp05_3_58));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007490(.in0(tmp05_0_58), .in1(tmp05_1_58), .out(tmp06_0_58));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007491(.in0(tmp05_2_58), .in1(tmp05_3_58), .out(tmp06_1_58));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add007492(.in0(tmp06_0_58), .in1(tmp06_1_58), .out(tmp07_0_58));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007493(.in0(tmp00_0_59), .in1(tmp00_1_59), .out(tmp01_0_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007494(.in0(tmp00_2_59), .in1(tmp00_3_59), .out(tmp01_1_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007495(.in0(tmp00_4_59), .in1(tmp00_5_59), .out(tmp01_2_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007496(.in0(tmp00_6_59), .in1(tmp00_7_59), .out(tmp01_3_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007497(.in0(tmp00_8_59), .in1(tmp00_9_59), .out(tmp01_4_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007498(.in0(tmp00_10_59), .in1(tmp00_11_59), .out(tmp01_5_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007499(.in0(tmp00_12_59), .in1(tmp00_13_59), .out(tmp01_6_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007500(.in0(tmp00_14_59), .in1(tmp00_15_59), .out(tmp01_7_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007501(.in0(tmp00_16_59), .in1(tmp00_17_59), .out(tmp01_8_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007502(.in0(tmp00_18_59), .in1(tmp00_19_59), .out(tmp01_9_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007503(.in0(tmp00_20_59), .in1(tmp00_21_59), .out(tmp01_10_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007504(.in0(tmp00_22_59), .in1(tmp00_23_59), .out(tmp01_11_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007505(.in0(tmp00_24_59), .in1(tmp00_25_59), .out(tmp01_12_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007506(.in0(tmp00_26_59), .in1(tmp00_27_59), .out(tmp01_13_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007507(.in0(tmp00_28_59), .in1(tmp00_29_59), .out(tmp01_14_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007508(.in0(tmp00_30_59), .in1(tmp00_31_59), .out(tmp01_15_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007509(.in0(tmp00_32_59), .in1(tmp00_33_59), .out(tmp01_16_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007510(.in0(tmp00_34_59), .in1(tmp00_35_59), .out(tmp01_17_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007511(.in0(tmp00_36_59), .in1(tmp00_37_59), .out(tmp01_18_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007512(.in0(tmp00_38_59), .in1(tmp00_39_59), .out(tmp01_19_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007513(.in0(tmp00_40_59), .in1(tmp00_41_59), .out(tmp01_20_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007514(.in0(tmp00_42_59), .in1(tmp00_43_59), .out(tmp01_21_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007515(.in0(tmp00_44_59), .in1(tmp00_45_59), .out(tmp01_22_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007516(.in0(tmp00_46_59), .in1(tmp00_47_59), .out(tmp01_23_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007517(.in0(tmp00_48_59), .in1(tmp00_49_59), .out(tmp01_24_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007518(.in0(tmp00_50_59), .in1(tmp00_51_59), .out(tmp01_25_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007519(.in0(tmp00_52_59), .in1(tmp00_53_59), .out(tmp01_26_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007520(.in0(tmp00_54_59), .in1(tmp00_55_59), .out(tmp01_27_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007521(.in0(tmp00_56_59), .in1(tmp00_57_59), .out(tmp01_28_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007522(.in0(tmp00_58_59), .in1(tmp00_59_59), .out(tmp01_29_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007523(.in0(tmp00_60_59), .in1(tmp00_61_59), .out(tmp01_30_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007524(.in0(tmp00_62_59), .in1(tmp00_63_59), .out(tmp01_31_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007525(.in0(tmp00_64_59), .in1(tmp00_65_59), .out(tmp01_32_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007526(.in0(tmp00_66_59), .in1(tmp00_67_59), .out(tmp01_33_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007527(.in0(tmp00_68_59), .in1(tmp00_69_59), .out(tmp01_34_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007528(.in0(tmp00_70_59), .in1(tmp00_71_59), .out(tmp01_35_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007529(.in0(tmp00_72_59), .in1(tmp00_73_59), .out(tmp01_36_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007530(.in0(tmp00_74_59), .in1(tmp00_75_59), .out(tmp01_37_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007531(.in0(tmp00_76_59), .in1(tmp00_77_59), .out(tmp01_38_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007532(.in0(tmp00_78_59), .in1(tmp00_79_59), .out(tmp01_39_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007533(.in0(tmp00_80_59), .in1(tmp00_81_59), .out(tmp01_40_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007534(.in0(tmp00_82_59), .in1(tmp00_83_59), .out(tmp01_41_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007535(.in0(tmp00_84_59), .in1(tmp00_85_59), .out(tmp01_42_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007536(.in0(tmp00_86_59), .in1(tmp00_87_59), .out(tmp01_43_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007537(.in0(tmp00_88_59), .in1(tmp00_89_59), .out(tmp01_44_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007538(.in0(tmp00_90_59), .in1(tmp00_91_59), .out(tmp01_45_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007539(.in0(tmp00_92_59), .in1(tmp00_93_59), .out(tmp01_46_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007540(.in0(tmp00_94_59), .in1(tmp00_95_59), .out(tmp01_47_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007541(.in0(tmp00_96_59), .in1(tmp00_97_59), .out(tmp01_48_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007542(.in0(tmp00_98_59), .in1(tmp00_99_59), .out(tmp01_49_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007543(.in0(tmp00_100_59), .in1(tmp00_101_59), .out(tmp01_50_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007544(.in0(tmp00_102_59), .in1(tmp00_103_59), .out(tmp01_51_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007545(.in0(tmp00_104_59), .in1(tmp00_105_59), .out(tmp01_52_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007546(.in0(tmp00_106_59), .in1(tmp00_107_59), .out(tmp01_53_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007547(.in0(tmp00_108_59), .in1(tmp00_109_59), .out(tmp01_54_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007548(.in0(tmp00_110_59), .in1(tmp00_111_59), .out(tmp01_55_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007549(.in0(tmp00_112_59), .in1(tmp00_113_59), .out(tmp01_56_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007550(.in0(tmp00_114_59), .in1(tmp00_115_59), .out(tmp01_57_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007551(.in0(tmp00_116_59), .in1(tmp00_117_59), .out(tmp01_58_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007552(.in0(tmp00_118_59), .in1(tmp00_119_59), .out(tmp01_59_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007553(.in0(tmp00_120_59), .in1(tmp00_121_59), .out(tmp01_60_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007554(.in0(tmp00_122_59), .in1(tmp00_123_59), .out(tmp01_61_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007555(.in0(tmp00_124_59), .in1(tmp00_125_59), .out(tmp01_62_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007556(.in0(tmp00_126_59), .in1(tmp00_127_59), .out(tmp01_63_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007557(.in0(tmp01_0_59), .in1(tmp01_1_59), .out(tmp02_0_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007558(.in0(tmp01_2_59), .in1(tmp01_3_59), .out(tmp02_1_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007559(.in0(tmp01_4_59), .in1(tmp01_5_59), .out(tmp02_2_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007560(.in0(tmp01_6_59), .in1(tmp01_7_59), .out(tmp02_3_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007561(.in0(tmp01_8_59), .in1(tmp01_9_59), .out(tmp02_4_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007562(.in0(tmp01_10_59), .in1(tmp01_11_59), .out(tmp02_5_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007563(.in0(tmp01_12_59), .in1(tmp01_13_59), .out(tmp02_6_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007564(.in0(tmp01_14_59), .in1(tmp01_15_59), .out(tmp02_7_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007565(.in0(tmp01_16_59), .in1(tmp01_17_59), .out(tmp02_8_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007566(.in0(tmp01_18_59), .in1(tmp01_19_59), .out(tmp02_9_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007567(.in0(tmp01_20_59), .in1(tmp01_21_59), .out(tmp02_10_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007568(.in0(tmp01_22_59), .in1(tmp01_23_59), .out(tmp02_11_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007569(.in0(tmp01_24_59), .in1(tmp01_25_59), .out(tmp02_12_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007570(.in0(tmp01_26_59), .in1(tmp01_27_59), .out(tmp02_13_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007571(.in0(tmp01_28_59), .in1(tmp01_29_59), .out(tmp02_14_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007572(.in0(tmp01_30_59), .in1(tmp01_31_59), .out(tmp02_15_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007573(.in0(tmp01_32_59), .in1(tmp01_33_59), .out(tmp02_16_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007574(.in0(tmp01_34_59), .in1(tmp01_35_59), .out(tmp02_17_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007575(.in0(tmp01_36_59), .in1(tmp01_37_59), .out(tmp02_18_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007576(.in0(tmp01_38_59), .in1(tmp01_39_59), .out(tmp02_19_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007577(.in0(tmp01_40_59), .in1(tmp01_41_59), .out(tmp02_20_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007578(.in0(tmp01_42_59), .in1(tmp01_43_59), .out(tmp02_21_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007579(.in0(tmp01_44_59), .in1(tmp01_45_59), .out(tmp02_22_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007580(.in0(tmp01_46_59), .in1(tmp01_47_59), .out(tmp02_23_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007581(.in0(tmp01_48_59), .in1(tmp01_49_59), .out(tmp02_24_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007582(.in0(tmp01_50_59), .in1(tmp01_51_59), .out(tmp02_25_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007583(.in0(tmp01_52_59), .in1(tmp01_53_59), .out(tmp02_26_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007584(.in0(tmp01_54_59), .in1(tmp01_55_59), .out(tmp02_27_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007585(.in0(tmp01_56_59), .in1(tmp01_57_59), .out(tmp02_28_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007586(.in0(tmp01_58_59), .in1(tmp01_59_59), .out(tmp02_29_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007587(.in0(tmp01_60_59), .in1(tmp01_61_59), .out(tmp02_30_59));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007588(.in0(tmp01_62_59), .in1(tmp01_63_59), .out(tmp02_31_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007589(.in0(tmp02_0_59), .in1(tmp02_1_59), .out(tmp03_0_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007590(.in0(tmp02_2_59), .in1(tmp02_3_59), .out(tmp03_1_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007591(.in0(tmp02_4_59), .in1(tmp02_5_59), .out(tmp03_2_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007592(.in0(tmp02_6_59), .in1(tmp02_7_59), .out(tmp03_3_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007593(.in0(tmp02_8_59), .in1(tmp02_9_59), .out(tmp03_4_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007594(.in0(tmp02_10_59), .in1(tmp02_11_59), .out(tmp03_5_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007595(.in0(tmp02_12_59), .in1(tmp02_13_59), .out(tmp03_6_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007596(.in0(tmp02_14_59), .in1(tmp02_15_59), .out(tmp03_7_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007597(.in0(tmp02_16_59), .in1(tmp02_17_59), .out(tmp03_8_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007598(.in0(tmp02_18_59), .in1(tmp02_19_59), .out(tmp03_9_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007599(.in0(tmp02_20_59), .in1(tmp02_21_59), .out(tmp03_10_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007600(.in0(tmp02_22_59), .in1(tmp02_23_59), .out(tmp03_11_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007601(.in0(tmp02_24_59), .in1(tmp02_25_59), .out(tmp03_12_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007602(.in0(tmp02_26_59), .in1(tmp02_27_59), .out(tmp03_13_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007603(.in0(tmp02_28_59), .in1(tmp02_29_59), .out(tmp03_14_59));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007604(.in0(tmp02_30_59), .in1(tmp02_31_59), .out(tmp03_15_59));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007605(.in0(tmp03_0_59), .in1(tmp03_1_59), .out(tmp04_0_59));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007606(.in0(tmp03_2_59), .in1(tmp03_3_59), .out(tmp04_1_59));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007607(.in0(tmp03_4_59), .in1(tmp03_5_59), .out(tmp04_2_59));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007608(.in0(tmp03_6_59), .in1(tmp03_7_59), .out(tmp04_3_59));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007609(.in0(tmp03_8_59), .in1(tmp03_9_59), .out(tmp04_4_59));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007610(.in0(tmp03_10_59), .in1(tmp03_11_59), .out(tmp04_5_59));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007611(.in0(tmp03_12_59), .in1(tmp03_13_59), .out(tmp04_6_59));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007612(.in0(tmp03_14_59), .in1(tmp03_15_59), .out(tmp04_7_59));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007613(.in0(tmp04_0_59), .in1(tmp04_1_59), .out(tmp05_0_59));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007614(.in0(tmp04_2_59), .in1(tmp04_3_59), .out(tmp05_1_59));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007615(.in0(tmp04_4_59), .in1(tmp04_5_59), .out(tmp05_2_59));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007616(.in0(tmp04_6_59), .in1(tmp04_7_59), .out(tmp05_3_59));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007617(.in0(tmp05_0_59), .in1(tmp05_1_59), .out(tmp06_0_59));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007618(.in0(tmp05_2_59), .in1(tmp05_3_59), .out(tmp06_1_59));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add007619(.in0(tmp06_0_59), .in1(tmp06_1_59), .out(tmp07_0_59));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007620(.in0(tmp00_0_60), .in1(tmp00_1_60), .out(tmp01_0_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007621(.in0(tmp00_2_60), .in1(tmp00_3_60), .out(tmp01_1_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007622(.in0(tmp00_4_60), .in1(tmp00_5_60), .out(tmp01_2_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007623(.in0(tmp00_6_60), .in1(tmp00_7_60), .out(tmp01_3_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007624(.in0(tmp00_8_60), .in1(tmp00_9_60), .out(tmp01_4_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007625(.in0(tmp00_10_60), .in1(tmp00_11_60), .out(tmp01_5_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007626(.in0(tmp00_12_60), .in1(tmp00_13_60), .out(tmp01_6_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007627(.in0(tmp00_14_60), .in1(tmp00_15_60), .out(tmp01_7_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007628(.in0(tmp00_16_60), .in1(tmp00_17_60), .out(tmp01_8_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007629(.in0(tmp00_18_60), .in1(tmp00_19_60), .out(tmp01_9_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007630(.in0(tmp00_20_60), .in1(tmp00_21_60), .out(tmp01_10_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007631(.in0(tmp00_22_60), .in1(tmp00_23_60), .out(tmp01_11_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007632(.in0(tmp00_24_60), .in1(tmp00_25_60), .out(tmp01_12_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007633(.in0(tmp00_26_60), .in1(tmp00_27_60), .out(tmp01_13_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007634(.in0(tmp00_28_60), .in1(tmp00_29_60), .out(tmp01_14_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007635(.in0(tmp00_30_60), .in1(tmp00_31_60), .out(tmp01_15_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007636(.in0(tmp00_32_60), .in1(tmp00_33_60), .out(tmp01_16_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007637(.in0(tmp00_34_60), .in1(tmp00_35_60), .out(tmp01_17_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007638(.in0(tmp00_36_60), .in1(tmp00_37_60), .out(tmp01_18_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007639(.in0(tmp00_38_60), .in1(tmp00_39_60), .out(tmp01_19_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007640(.in0(tmp00_40_60), .in1(tmp00_41_60), .out(tmp01_20_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007641(.in0(tmp00_42_60), .in1(tmp00_43_60), .out(tmp01_21_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007642(.in0(tmp00_44_60), .in1(tmp00_45_60), .out(tmp01_22_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007643(.in0(tmp00_46_60), .in1(tmp00_47_60), .out(tmp01_23_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007644(.in0(tmp00_48_60), .in1(tmp00_49_60), .out(tmp01_24_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007645(.in0(tmp00_50_60), .in1(tmp00_51_60), .out(tmp01_25_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007646(.in0(tmp00_52_60), .in1(tmp00_53_60), .out(tmp01_26_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007647(.in0(tmp00_54_60), .in1(tmp00_55_60), .out(tmp01_27_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007648(.in0(tmp00_56_60), .in1(tmp00_57_60), .out(tmp01_28_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007649(.in0(tmp00_58_60), .in1(tmp00_59_60), .out(tmp01_29_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007650(.in0(tmp00_60_60), .in1(tmp00_61_60), .out(tmp01_30_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007651(.in0(tmp00_62_60), .in1(tmp00_63_60), .out(tmp01_31_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007652(.in0(tmp00_64_60), .in1(tmp00_65_60), .out(tmp01_32_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007653(.in0(tmp00_66_60), .in1(tmp00_67_60), .out(tmp01_33_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007654(.in0(tmp00_68_60), .in1(tmp00_69_60), .out(tmp01_34_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007655(.in0(tmp00_70_60), .in1(tmp00_71_60), .out(tmp01_35_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007656(.in0(tmp00_72_60), .in1(tmp00_73_60), .out(tmp01_36_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007657(.in0(tmp00_74_60), .in1(tmp00_75_60), .out(tmp01_37_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007658(.in0(tmp00_76_60), .in1(tmp00_77_60), .out(tmp01_38_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007659(.in0(tmp00_78_60), .in1(tmp00_79_60), .out(tmp01_39_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007660(.in0(tmp00_80_60), .in1(tmp00_81_60), .out(tmp01_40_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007661(.in0(tmp00_82_60), .in1(tmp00_83_60), .out(tmp01_41_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007662(.in0(tmp00_84_60), .in1(tmp00_85_60), .out(tmp01_42_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007663(.in0(tmp00_86_60), .in1(tmp00_87_60), .out(tmp01_43_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007664(.in0(tmp00_88_60), .in1(tmp00_89_60), .out(tmp01_44_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007665(.in0(tmp00_90_60), .in1(tmp00_91_60), .out(tmp01_45_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007666(.in0(tmp00_92_60), .in1(tmp00_93_60), .out(tmp01_46_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007667(.in0(tmp00_94_60), .in1(tmp00_95_60), .out(tmp01_47_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007668(.in0(tmp00_96_60), .in1(tmp00_97_60), .out(tmp01_48_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007669(.in0(tmp00_98_60), .in1(tmp00_99_60), .out(tmp01_49_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007670(.in0(tmp00_100_60), .in1(tmp00_101_60), .out(tmp01_50_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007671(.in0(tmp00_102_60), .in1(tmp00_103_60), .out(tmp01_51_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007672(.in0(tmp00_104_60), .in1(tmp00_105_60), .out(tmp01_52_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007673(.in0(tmp00_106_60), .in1(tmp00_107_60), .out(tmp01_53_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007674(.in0(tmp00_108_60), .in1(tmp00_109_60), .out(tmp01_54_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007675(.in0(tmp00_110_60), .in1(tmp00_111_60), .out(tmp01_55_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007676(.in0(tmp00_112_60), .in1(tmp00_113_60), .out(tmp01_56_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007677(.in0(tmp00_114_60), .in1(tmp00_115_60), .out(tmp01_57_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007678(.in0(tmp00_116_60), .in1(tmp00_117_60), .out(tmp01_58_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007679(.in0(tmp00_118_60), .in1(tmp00_119_60), .out(tmp01_59_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007680(.in0(tmp00_120_60), .in1(tmp00_121_60), .out(tmp01_60_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007681(.in0(tmp00_122_60), .in1(tmp00_123_60), .out(tmp01_61_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007682(.in0(tmp00_124_60), .in1(tmp00_125_60), .out(tmp01_62_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007683(.in0(tmp00_126_60), .in1(tmp00_127_60), .out(tmp01_63_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007684(.in0(tmp01_0_60), .in1(tmp01_1_60), .out(tmp02_0_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007685(.in0(tmp01_2_60), .in1(tmp01_3_60), .out(tmp02_1_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007686(.in0(tmp01_4_60), .in1(tmp01_5_60), .out(tmp02_2_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007687(.in0(tmp01_6_60), .in1(tmp01_7_60), .out(tmp02_3_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007688(.in0(tmp01_8_60), .in1(tmp01_9_60), .out(tmp02_4_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007689(.in0(tmp01_10_60), .in1(tmp01_11_60), .out(tmp02_5_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007690(.in0(tmp01_12_60), .in1(tmp01_13_60), .out(tmp02_6_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007691(.in0(tmp01_14_60), .in1(tmp01_15_60), .out(tmp02_7_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007692(.in0(tmp01_16_60), .in1(tmp01_17_60), .out(tmp02_8_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007693(.in0(tmp01_18_60), .in1(tmp01_19_60), .out(tmp02_9_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007694(.in0(tmp01_20_60), .in1(tmp01_21_60), .out(tmp02_10_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007695(.in0(tmp01_22_60), .in1(tmp01_23_60), .out(tmp02_11_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007696(.in0(tmp01_24_60), .in1(tmp01_25_60), .out(tmp02_12_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007697(.in0(tmp01_26_60), .in1(tmp01_27_60), .out(tmp02_13_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007698(.in0(tmp01_28_60), .in1(tmp01_29_60), .out(tmp02_14_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007699(.in0(tmp01_30_60), .in1(tmp01_31_60), .out(tmp02_15_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007700(.in0(tmp01_32_60), .in1(tmp01_33_60), .out(tmp02_16_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007701(.in0(tmp01_34_60), .in1(tmp01_35_60), .out(tmp02_17_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007702(.in0(tmp01_36_60), .in1(tmp01_37_60), .out(tmp02_18_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007703(.in0(tmp01_38_60), .in1(tmp01_39_60), .out(tmp02_19_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007704(.in0(tmp01_40_60), .in1(tmp01_41_60), .out(tmp02_20_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007705(.in0(tmp01_42_60), .in1(tmp01_43_60), .out(tmp02_21_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007706(.in0(tmp01_44_60), .in1(tmp01_45_60), .out(tmp02_22_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007707(.in0(tmp01_46_60), .in1(tmp01_47_60), .out(tmp02_23_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007708(.in0(tmp01_48_60), .in1(tmp01_49_60), .out(tmp02_24_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007709(.in0(tmp01_50_60), .in1(tmp01_51_60), .out(tmp02_25_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007710(.in0(tmp01_52_60), .in1(tmp01_53_60), .out(tmp02_26_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007711(.in0(tmp01_54_60), .in1(tmp01_55_60), .out(tmp02_27_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007712(.in0(tmp01_56_60), .in1(tmp01_57_60), .out(tmp02_28_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007713(.in0(tmp01_58_60), .in1(tmp01_59_60), .out(tmp02_29_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007714(.in0(tmp01_60_60), .in1(tmp01_61_60), .out(tmp02_30_60));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007715(.in0(tmp01_62_60), .in1(tmp01_63_60), .out(tmp02_31_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007716(.in0(tmp02_0_60), .in1(tmp02_1_60), .out(tmp03_0_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007717(.in0(tmp02_2_60), .in1(tmp02_3_60), .out(tmp03_1_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007718(.in0(tmp02_4_60), .in1(tmp02_5_60), .out(tmp03_2_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007719(.in0(tmp02_6_60), .in1(tmp02_7_60), .out(tmp03_3_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007720(.in0(tmp02_8_60), .in1(tmp02_9_60), .out(tmp03_4_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007721(.in0(tmp02_10_60), .in1(tmp02_11_60), .out(tmp03_5_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007722(.in0(tmp02_12_60), .in1(tmp02_13_60), .out(tmp03_6_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007723(.in0(tmp02_14_60), .in1(tmp02_15_60), .out(tmp03_7_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007724(.in0(tmp02_16_60), .in1(tmp02_17_60), .out(tmp03_8_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007725(.in0(tmp02_18_60), .in1(tmp02_19_60), .out(tmp03_9_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007726(.in0(tmp02_20_60), .in1(tmp02_21_60), .out(tmp03_10_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007727(.in0(tmp02_22_60), .in1(tmp02_23_60), .out(tmp03_11_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007728(.in0(tmp02_24_60), .in1(tmp02_25_60), .out(tmp03_12_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007729(.in0(tmp02_26_60), .in1(tmp02_27_60), .out(tmp03_13_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007730(.in0(tmp02_28_60), .in1(tmp02_29_60), .out(tmp03_14_60));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007731(.in0(tmp02_30_60), .in1(tmp02_31_60), .out(tmp03_15_60));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007732(.in0(tmp03_0_60), .in1(tmp03_1_60), .out(tmp04_0_60));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007733(.in0(tmp03_2_60), .in1(tmp03_3_60), .out(tmp04_1_60));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007734(.in0(tmp03_4_60), .in1(tmp03_5_60), .out(tmp04_2_60));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007735(.in0(tmp03_6_60), .in1(tmp03_7_60), .out(tmp04_3_60));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007736(.in0(tmp03_8_60), .in1(tmp03_9_60), .out(tmp04_4_60));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007737(.in0(tmp03_10_60), .in1(tmp03_11_60), .out(tmp04_5_60));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007738(.in0(tmp03_12_60), .in1(tmp03_13_60), .out(tmp04_6_60));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007739(.in0(tmp03_14_60), .in1(tmp03_15_60), .out(tmp04_7_60));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007740(.in0(tmp04_0_60), .in1(tmp04_1_60), .out(tmp05_0_60));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007741(.in0(tmp04_2_60), .in1(tmp04_3_60), .out(tmp05_1_60));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007742(.in0(tmp04_4_60), .in1(tmp04_5_60), .out(tmp05_2_60));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007743(.in0(tmp04_6_60), .in1(tmp04_7_60), .out(tmp05_3_60));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007744(.in0(tmp05_0_60), .in1(tmp05_1_60), .out(tmp06_0_60));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007745(.in0(tmp05_2_60), .in1(tmp05_3_60), .out(tmp06_1_60));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add007746(.in0(tmp06_0_60), .in1(tmp06_1_60), .out(tmp07_0_60));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007747(.in0(tmp00_0_61), .in1(tmp00_1_61), .out(tmp01_0_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007748(.in0(tmp00_2_61), .in1(tmp00_3_61), .out(tmp01_1_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007749(.in0(tmp00_4_61), .in1(tmp00_5_61), .out(tmp01_2_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007750(.in0(tmp00_6_61), .in1(tmp00_7_61), .out(tmp01_3_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007751(.in0(tmp00_8_61), .in1(tmp00_9_61), .out(tmp01_4_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007752(.in0(tmp00_10_61), .in1(tmp00_11_61), .out(tmp01_5_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007753(.in0(tmp00_12_61), .in1(tmp00_13_61), .out(tmp01_6_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007754(.in0(tmp00_14_61), .in1(tmp00_15_61), .out(tmp01_7_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007755(.in0(tmp00_16_61), .in1(tmp00_17_61), .out(tmp01_8_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007756(.in0(tmp00_18_61), .in1(tmp00_19_61), .out(tmp01_9_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007757(.in0(tmp00_20_61), .in1(tmp00_21_61), .out(tmp01_10_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007758(.in0(tmp00_22_61), .in1(tmp00_23_61), .out(tmp01_11_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007759(.in0(tmp00_24_61), .in1(tmp00_25_61), .out(tmp01_12_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007760(.in0(tmp00_26_61), .in1(tmp00_27_61), .out(tmp01_13_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007761(.in0(tmp00_28_61), .in1(tmp00_29_61), .out(tmp01_14_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007762(.in0(tmp00_30_61), .in1(tmp00_31_61), .out(tmp01_15_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007763(.in0(tmp00_32_61), .in1(tmp00_33_61), .out(tmp01_16_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007764(.in0(tmp00_34_61), .in1(tmp00_35_61), .out(tmp01_17_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007765(.in0(tmp00_36_61), .in1(tmp00_37_61), .out(tmp01_18_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007766(.in0(tmp00_38_61), .in1(tmp00_39_61), .out(tmp01_19_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007767(.in0(tmp00_40_61), .in1(tmp00_41_61), .out(tmp01_20_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007768(.in0(tmp00_42_61), .in1(tmp00_43_61), .out(tmp01_21_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007769(.in0(tmp00_44_61), .in1(tmp00_45_61), .out(tmp01_22_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007770(.in0(tmp00_46_61), .in1(tmp00_47_61), .out(tmp01_23_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007771(.in0(tmp00_48_61), .in1(tmp00_49_61), .out(tmp01_24_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007772(.in0(tmp00_50_61), .in1(tmp00_51_61), .out(tmp01_25_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007773(.in0(tmp00_52_61), .in1(tmp00_53_61), .out(tmp01_26_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007774(.in0(tmp00_54_61), .in1(tmp00_55_61), .out(tmp01_27_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007775(.in0(tmp00_56_61), .in1(tmp00_57_61), .out(tmp01_28_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007776(.in0(tmp00_58_61), .in1(tmp00_59_61), .out(tmp01_29_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007777(.in0(tmp00_60_61), .in1(tmp00_61_61), .out(tmp01_30_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007778(.in0(tmp00_62_61), .in1(tmp00_63_61), .out(tmp01_31_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007779(.in0(tmp00_64_61), .in1(tmp00_65_61), .out(tmp01_32_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007780(.in0(tmp00_66_61), .in1(tmp00_67_61), .out(tmp01_33_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007781(.in0(tmp00_68_61), .in1(tmp00_69_61), .out(tmp01_34_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007782(.in0(tmp00_70_61), .in1(tmp00_71_61), .out(tmp01_35_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007783(.in0(tmp00_72_61), .in1(tmp00_73_61), .out(tmp01_36_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007784(.in0(tmp00_74_61), .in1(tmp00_75_61), .out(tmp01_37_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007785(.in0(tmp00_76_61), .in1(tmp00_77_61), .out(tmp01_38_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007786(.in0(tmp00_78_61), .in1(tmp00_79_61), .out(tmp01_39_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007787(.in0(tmp00_80_61), .in1(tmp00_81_61), .out(tmp01_40_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007788(.in0(tmp00_82_61), .in1(tmp00_83_61), .out(tmp01_41_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007789(.in0(tmp00_84_61), .in1(tmp00_85_61), .out(tmp01_42_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007790(.in0(tmp00_86_61), .in1(tmp00_87_61), .out(tmp01_43_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007791(.in0(tmp00_88_61), .in1(tmp00_89_61), .out(tmp01_44_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007792(.in0(tmp00_90_61), .in1(tmp00_91_61), .out(tmp01_45_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007793(.in0(tmp00_92_61), .in1(tmp00_93_61), .out(tmp01_46_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007794(.in0(tmp00_94_61), .in1(tmp00_95_61), .out(tmp01_47_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007795(.in0(tmp00_96_61), .in1(tmp00_97_61), .out(tmp01_48_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007796(.in0(tmp00_98_61), .in1(tmp00_99_61), .out(tmp01_49_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007797(.in0(tmp00_100_61), .in1(tmp00_101_61), .out(tmp01_50_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007798(.in0(tmp00_102_61), .in1(tmp00_103_61), .out(tmp01_51_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007799(.in0(tmp00_104_61), .in1(tmp00_105_61), .out(tmp01_52_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007800(.in0(tmp00_106_61), .in1(tmp00_107_61), .out(tmp01_53_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007801(.in0(tmp00_108_61), .in1(tmp00_109_61), .out(tmp01_54_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007802(.in0(tmp00_110_61), .in1(tmp00_111_61), .out(tmp01_55_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007803(.in0(tmp00_112_61), .in1(tmp00_113_61), .out(tmp01_56_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007804(.in0(tmp00_114_61), .in1(tmp00_115_61), .out(tmp01_57_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007805(.in0(tmp00_116_61), .in1(tmp00_117_61), .out(tmp01_58_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007806(.in0(tmp00_118_61), .in1(tmp00_119_61), .out(tmp01_59_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007807(.in0(tmp00_120_61), .in1(tmp00_121_61), .out(tmp01_60_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007808(.in0(tmp00_122_61), .in1(tmp00_123_61), .out(tmp01_61_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007809(.in0(tmp00_124_61), .in1(tmp00_125_61), .out(tmp01_62_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007810(.in0(tmp00_126_61), .in1(tmp00_127_61), .out(tmp01_63_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007811(.in0(tmp01_0_61), .in1(tmp01_1_61), .out(tmp02_0_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007812(.in0(tmp01_2_61), .in1(tmp01_3_61), .out(tmp02_1_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007813(.in0(tmp01_4_61), .in1(tmp01_5_61), .out(tmp02_2_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007814(.in0(tmp01_6_61), .in1(tmp01_7_61), .out(tmp02_3_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007815(.in0(tmp01_8_61), .in1(tmp01_9_61), .out(tmp02_4_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007816(.in0(tmp01_10_61), .in1(tmp01_11_61), .out(tmp02_5_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007817(.in0(tmp01_12_61), .in1(tmp01_13_61), .out(tmp02_6_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007818(.in0(tmp01_14_61), .in1(tmp01_15_61), .out(tmp02_7_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007819(.in0(tmp01_16_61), .in1(tmp01_17_61), .out(tmp02_8_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007820(.in0(tmp01_18_61), .in1(tmp01_19_61), .out(tmp02_9_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007821(.in0(tmp01_20_61), .in1(tmp01_21_61), .out(tmp02_10_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007822(.in0(tmp01_22_61), .in1(tmp01_23_61), .out(tmp02_11_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007823(.in0(tmp01_24_61), .in1(tmp01_25_61), .out(tmp02_12_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007824(.in0(tmp01_26_61), .in1(tmp01_27_61), .out(tmp02_13_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007825(.in0(tmp01_28_61), .in1(tmp01_29_61), .out(tmp02_14_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007826(.in0(tmp01_30_61), .in1(tmp01_31_61), .out(tmp02_15_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007827(.in0(tmp01_32_61), .in1(tmp01_33_61), .out(tmp02_16_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007828(.in0(tmp01_34_61), .in1(tmp01_35_61), .out(tmp02_17_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007829(.in0(tmp01_36_61), .in1(tmp01_37_61), .out(tmp02_18_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007830(.in0(tmp01_38_61), .in1(tmp01_39_61), .out(tmp02_19_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007831(.in0(tmp01_40_61), .in1(tmp01_41_61), .out(tmp02_20_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007832(.in0(tmp01_42_61), .in1(tmp01_43_61), .out(tmp02_21_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007833(.in0(tmp01_44_61), .in1(tmp01_45_61), .out(tmp02_22_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007834(.in0(tmp01_46_61), .in1(tmp01_47_61), .out(tmp02_23_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007835(.in0(tmp01_48_61), .in1(tmp01_49_61), .out(tmp02_24_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007836(.in0(tmp01_50_61), .in1(tmp01_51_61), .out(tmp02_25_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007837(.in0(tmp01_52_61), .in1(tmp01_53_61), .out(tmp02_26_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007838(.in0(tmp01_54_61), .in1(tmp01_55_61), .out(tmp02_27_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007839(.in0(tmp01_56_61), .in1(tmp01_57_61), .out(tmp02_28_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007840(.in0(tmp01_58_61), .in1(tmp01_59_61), .out(tmp02_29_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007841(.in0(tmp01_60_61), .in1(tmp01_61_61), .out(tmp02_30_61));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007842(.in0(tmp01_62_61), .in1(tmp01_63_61), .out(tmp02_31_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007843(.in0(tmp02_0_61), .in1(tmp02_1_61), .out(tmp03_0_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007844(.in0(tmp02_2_61), .in1(tmp02_3_61), .out(tmp03_1_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007845(.in0(tmp02_4_61), .in1(tmp02_5_61), .out(tmp03_2_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007846(.in0(tmp02_6_61), .in1(tmp02_7_61), .out(tmp03_3_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007847(.in0(tmp02_8_61), .in1(tmp02_9_61), .out(tmp03_4_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007848(.in0(tmp02_10_61), .in1(tmp02_11_61), .out(tmp03_5_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007849(.in0(tmp02_12_61), .in1(tmp02_13_61), .out(tmp03_6_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007850(.in0(tmp02_14_61), .in1(tmp02_15_61), .out(tmp03_7_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007851(.in0(tmp02_16_61), .in1(tmp02_17_61), .out(tmp03_8_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007852(.in0(tmp02_18_61), .in1(tmp02_19_61), .out(tmp03_9_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007853(.in0(tmp02_20_61), .in1(tmp02_21_61), .out(tmp03_10_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007854(.in0(tmp02_22_61), .in1(tmp02_23_61), .out(tmp03_11_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007855(.in0(tmp02_24_61), .in1(tmp02_25_61), .out(tmp03_12_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007856(.in0(tmp02_26_61), .in1(tmp02_27_61), .out(tmp03_13_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007857(.in0(tmp02_28_61), .in1(tmp02_29_61), .out(tmp03_14_61));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007858(.in0(tmp02_30_61), .in1(tmp02_31_61), .out(tmp03_15_61));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007859(.in0(tmp03_0_61), .in1(tmp03_1_61), .out(tmp04_0_61));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007860(.in0(tmp03_2_61), .in1(tmp03_3_61), .out(tmp04_1_61));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007861(.in0(tmp03_4_61), .in1(tmp03_5_61), .out(tmp04_2_61));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007862(.in0(tmp03_6_61), .in1(tmp03_7_61), .out(tmp04_3_61));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007863(.in0(tmp03_8_61), .in1(tmp03_9_61), .out(tmp04_4_61));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007864(.in0(tmp03_10_61), .in1(tmp03_11_61), .out(tmp04_5_61));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007865(.in0(tmp03_12_61), .in1(tmp03_13_61), .out(tmp04_6_61));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007866(.in0(tmp03_14_61), .in1(tmp03_15_61), .out(tmp04_7_61));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007867(.in0(tmp04_0_61), .in1(tmp04_1_61), .out(tmp05_0_61));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007868(.in0(tmp04_2_61), .in1(tmp04_3_61), .out(tmp05_1_61));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007869(.in0(tmp04_4_61), .in1(tmp04_5_61), .out(tmp05_2_61));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007870(.in0(tmp04_6_61), .in1(tmp04_7_61), .out(tmp05_3_61));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007871(.in0(tmp05_0_61), .in1(tmp05_1_61), .out(tmp06_0_61));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007872(.in0(tmp05_2_61), .in1(tmp05_3_61), .out(tmp06_1_61));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add007873(.in0(tmp06_0_61), .in1(tmp06_1_61), .out(tmp07_0_61));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007874(.in0(tmp00_0_62), .in1(tmp00_1_62), .out(tmp01_0_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007875(.in0(tmp00_2_62), .in1(tmp00_3_62), .out(tmp01_1_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007876(.in0(tmp00_4_62), .in1(tmp00_5_62), .out(tmp01_2_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007877(.in0(tmp00_6_62), .in1(tmp00_7_62), .out(tmp01_3_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007878(.in0(tmp00_8_62), .in1(tmp00_9_62), .out(tmp01_4_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007879(.in0(tmp00_10_62), .in1(tmp00_11_62), .out(tmp01_5_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007880(.in0(tmp00_12_62), .in1(tmp00_13_62), .out(tmp01_6_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007881(.in0(tmp00_14_62), .in1(tmp00_15_62), .out(tmp01_7_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007882(.in0(tmp00_16_62), .in1(tmp00_17_62), .out(tmp01_8_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007883(.in0(tmp00_18_62), .in1(tmp00_19_62), .out(tmp01_9_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007884(.in0(tmp00_20_62), .in1(tmp00_21_62), .out(tmp01_10_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007885(.in0(tmp00_22_62), .in1(tmp00_23_62), .out(tmp01_11_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007886(.in0(tmp00_24_62), .in1(tmp00_25_62), .out(tmp01_12_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007887(.in0(tmp00_26_62), .in1(tmp00_27_62), .out(tmp01_13_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007888(.in0(tmp00_28_62), .in1(tmp00_29_62), .out(tmp01_14_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007889(.in0(tmp00_30_62), .in1(tmp00_31_62), .out(tmp01_15_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007890(.in0(tmp00_32_62), .in1(tmp00_33_62), .out(tmp01_16_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007891(.in0(tmp00_34_62), .in1(tmp00_35_62), .out(tmp01_17_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007892(.in0(tmp00_36_62), .in1(tmp00_37_62), .out(tmp01_18_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007893(.in0(tmp00_38_62), .in1(tmp00_39_62), .out(tmp01_19_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007894(.in0(tmp00_40_62), .in1(tmp00_41_62), .out(tmp01_20_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007895(.in0(tmp00_42_62), .in1(tmp00_43_62), .out(tmp01_21_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007896(.in0(tmp00_44_62), .in1(tmp00_45_62), .out(tmp01_22_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007897(.in0(tmp00_46_62), .in1(tmp00_47_62), .out(tmp01_23_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007898(.in0(tmp00_48_62), .in1(tmp00_49_62), .out(tmp01_24_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007899(.in0(tmp00_50_62), .in1(tmp00_51_62), .out(tmp01_25_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007900(.in0(tmp00_52_62), .in1(tmp00_53_62), .out(tmp01_26_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007901(.in0(tmp00_54_62), .in1(tmp00_55_62), .out(tmp01_27_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007902(.in0(tmp00_56_62), .in1(tmp00_57_62), .out(tmp01_28_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007903(.in0(tmp00_58_62), .in1(tmp00_59_62), .out(tmp01_29_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007904(.in0(tmp00_60_62), .in1(tmp00_61_62), .out(tmp01_30_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007905(.in0(tmp00_62_62), .in1(tmp00_63_62), .out(tmp01_31_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007906(.in0(tmp00_64_62), .in1(tmp00_65_62), .out(tmp01_32_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007907(.in0(tmp00_66_62), .in1(tmp00_67_62), .out(tmp01_33_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007908(.in0(tmp00_68_62), .in1(tmp00_69_62), .out(tmp01_34_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007909(.in0(tmp00_70_62), .in1(tmp00_71_62), .out(tmp01_35_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007910(.in0(tmp00_72_62), .in1(tmp00_73_62), .out(tmp01_36_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007911(.in0(tmp00_74_62), .in1(tmp00_75_62), .out(tmp01_37_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007912(.in0(tmp00_76_62), .in1(tmp00_77_62), .out(tmp01_38_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007913(.in0(tmp00_78_62), .in1(tmp00_79_62), .out(tmp01_39_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007914(.in0(tmp00_80_62), .in1(tmp00_81_62), .out(tmp01_40_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007915(.in0(tmp00_82_62), .in1(tmp00_83_62), .out(tmp01_41_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007916(.in0(tmp00_84_62), .in1(tmp00_85_62), .out(tmp01_42_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007917(.in0(tmp00_86_62), .in1(tmp00_87_62), .out(tmp01_43_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007918(.in0(tmp00_88_62), .in1(tmp00_89_62), .out(tmp01_44_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007919(.in0(tmp00_90_62), .in1(tmp00_91_62), .out(tmp01_45_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007920(.in0(tmp00_92_62), .in1(tmp00_93_62), .out(tmp01_46_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007921(.in0(tmp00_94_62), .in1(tmp00_95_62), .out(tmp01_47_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007922(.in0(tmp00_96_62), .in1(tmp00_97_62), .out(tmp01_48_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007923(.in0(tmp00_98_62), .in1(tmp00_99_62), .out(tmp01_49_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007924(.in0(tmp00_100_62), .in1(tmp00_101_62), .out(tmp01_50_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007925(.in0(tmp00_102_62), .in1(tmp00_103_62), .out(tmp01_51_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007926(.in0(tmp00_104_62), .in1(tmp00_105_62), .out(tmp01_52_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007927(.in0(tmp00_106_62), .in1(tmp00_107_62), .out(tmp01_53_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007928(.in0(tmp00_108_62), .in1(tmp00_109_62), .out(tmp01_54_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007929(.in0(tmp00_110_62), .in1(tmp00_111_62), .out(tmp01_55_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007930(.in0(tmp00_112_62), .in1(tmp00_113_62), .out(tmp01_56_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007931(.in0(tmp00_114_62), .in1(tmp00_115_62), .out(tmp01_57_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007932(.in0(tmp00_116_62), .in1(tmp00_117_62), .out(tmp01_58_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007933(.in0(tmp00_118_62), .in1(tmp00_119_62), .out(tmp01_59_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007934(.in0(tmp00_120_62), .in1(tmp00_121_62), .out(tmp01_60_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007935(.in0(tmp00_122_62), .in1(tmp00_123_62), .out(tmp01_61_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007936(.in0(tmp00_124_62), .in1(tmp00_125_62), .out(tmp01_62_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add007937(.in0(tmp00_126_62), .in1(tmp00_127_62), .out(tmp01_63_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007938(.in0(tmp01_0_62), .in1(tmp01_1_62), .out(tmp02_0_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007939(.in0(tmp01_2_62), .in1(tmp01_3_62), .out(tmp02_1_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007940(.in0(tmp01_4_62), .in1(tmp01_5_62), .out(tmp02_2_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007941(.in0(tmp01_6_62), .in1(tmp01_7_62), .out(tmp02_3_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007942(.in0(tmp01_8_62), .in1(tmp01_9_62), .out(tmp02_4_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007943(.in0(tmp01_10_62), .in1(tmp01_11_62), .out(tmp02_5_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007944(.in0(tmp01_12_62), .in1(tmp01_13_62), .out(tmp02_6_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007945(.in0(tmp01_14_62), .in1(tmp01_15_62), .out(tmp02_7_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007946(.in0(tmp01_16_62), .in1(tmp01_17_62), .out(tmp02_8_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007947(.in0(tmp01_18_62), .in1(tmp01_19_62), .out(tmp02_9_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007948(.in0(tmp01_20_62), .in1(tmp01_21_62), .out(tmp02_10_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007949(.in0(tmp01_22_62), .in1(tmp01_23_62), .out(tmp02_11_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007950(.in0(tmp01_24_62), .in1(tmp01_25_62), .out(tmp02_12_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007951(.in0(tmp01_26_62), .in1(tmp01_27_62), .out(tmp02_13_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007952(.in0(tmp01_28_62), .in1(tmp01_29_62), .out(tmp02_14_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007953(.in0(tmp01_30_62), .in1(tmp01_31_62), .out(tmp02_15_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007954(.in0(tmp01_32_62), .in1(tmp01_33_62), .out(tmp02_16_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007955(.in0(tmp01_34_62), .in1(tmp01_35_62), .out(tmp02_17_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007956(.in0(tmp01_36_62), .in1(tmp01_37_62), .out(tmp02_18_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007957(.in0(tmp01_38_62), .in1(tmp01_39_62), .out(tmp02_19_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007958(.in0(tmp01_40_62), .in1(tmp01_41_62), .out(tmp02_20_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007959(.in0(tmp01_42_62), .in1(tmp01_43_62), .out(tmp02_21_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007960(.in0(tmp01_44_62), .in1(tmp01_45_62), .out(tmp02_22_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007961(.in0(tmp01_46_62), .in1(tmp01_47_62), .out(tmp02_23_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007962(.in0(tmp01_48_62), .in1(tmp01_49_62), .out(tmp02_24_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007963(.in0(tmp01_50_62), .in1(tmp01_51_62), .out(tmp02_25_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007964(.in0(tmp01_52_62), .in1(tmp01_53_62), .out(tmp02_26_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007965(.in0(tmp01_54_62), .in1(tmp01_55_62), .out(tmp02_27_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007966(.in0(tmp01_56_62), .in1(tmp01_57_62), .out(tmp02_28_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007967(.in0(tmp01_58_62), .in1(tmp01_59_62), .out(tmp02_29_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007968(.in0(tmp01_60_62), .in1(tmp01_61_62), .out(tmp02_30_62));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add007969(.in0(tmp01_62_62), .in1(tmp01_63_62), .out(tmp02_31_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007970(.in0(tmp02_0_62), .in1(tmp02_1_62), .out(tmp03_0_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007971(.in0(tmp02_2_62), .in1(tmp02_3_62), .out(tmp03_1_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007972(.in0(tmp02_4_62), .in1(tmp02_5_62), .out(tmp03_2_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007973(.in0(tmp02_6_62), .in1(tmp02_7_62), .out(tmp03_3_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007974(.in0(tmp02_8_62), .in1(tmp02_9_62), .out(tmp03_4_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007975(.in0(tmp02_10_62), .in1(tmp02_11_62), .out(tmp03_5_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007976(.in0(tmp02_12_62), .in1(tmp02_13_62), .out(tmp03_6_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007977(.in0(tmp02_14_62), .in1(tmp02_15_62), .out(tmp03_7_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007978(.in0(tmp02_16_62), .in1(tmp02_17_62), .out(tmp03_8_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007979(.in0(tmp02_18_62), .in1(tmp02_19_62), .out(tmp03_9_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007980(.in0(tmp02_20_62), .in1(tmp02_21_62), .out(tmp03_10_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007981(.in0(tmp02_22_62), .in1(tmp02_23_62), .out(tmp03_11_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007982(.in0(tmp02_24_62), .in1(tmp02_25_62), .out(tmp03_12_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007983(.in0(tmp02_26_62), .in1(tmp02_27_62), .out(tmp03_13_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007984(.in0(tmp02_28_62), .in1(tmp02_29_62), .out(tmp03_14_62));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add007985(.in0(tmp02_30_62), .in1(tmp02_31_62), .out(tmp03_15_62));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007986(.in0(tmp03_0_62), .in1(tmp03_1_62), .out(tmp04_0_62));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007987(.in0(tmp03_2_62), .in1(tmp03_3_62), .out(tmp04_1_62));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007988(.in0(tmp03_4_62), .in1(tmp03_5_62), .out(tmp04_2_62));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007989(.in0(tmp03_6_62), .in1(tmp03_7_62), .out(tmp04_3_62));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007990(.in0(tmp03_8_62), .in1(tmp03_9_62), .out(tmp04_4_62));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007991(.in0(tmp03_10_62), .in1(tmp03_11_62), .out(tmp04_5_62));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007992(.in0(tmp03_12_62), .in1(tmp03_13_62), .out(tmp04_6_62));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add007993(.in0(tmp03_14_62), .in1(tmp03_15_62), .out(tmp04_7_62));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007994(.in0(tmp04_0_62), .in1(tmp04_1_62), .out(tmp05_0_62));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007995(.in0(tmp04_2_62), .in1(tmp04_3_62), .out(tmp05_1_62));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007996(.in0(tmp04_4_62), .in1(tmp04_5_62), .out(tmp05_2_62));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add007997(.in0(tmp04_6_62), .in1(tmp04_7_62), .out(tmp05_3_62));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007998(.in0(tmp05_0_62), .in1(tmp05_1_62), .out(tmp06_0_62));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add007999(.in0(tmp05_2_62), .in1(tmp05_3_62), .out(tmp06_1_62));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add008000(.in0(tmp06_0_62), .in1(tmp06_1_62), .out(tmp07_0_62));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008001(.in0(tmp00_0_63), .in1(tmp00_1_63), .out(tmp01_0_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008002(.in0(tmp00_2_63), .in1(tmp00_3_63), .out(tmp01_1_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008003(.in0(tmp00_4_63), .in1(tmp00_5_63), .out(tmp01_2_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008004(.in0(tmp00_6_63), .in1(tmp00_7_63), .out(tmp01_3_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008005(.in0(tmp00_8_63), .in1(tmp00_9_63), .out(tmp01_4_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008006(.in0(tmp00_10_63), .in1(tmp00_11_63), .out(tmp01_5_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008007(.in0(tmp00_12_63), .in1(tmp00_13_63), .out(tmp01_6_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008008(.in0(tmp00_14_63), .in1(tmp00_15_63), .out(tmp01_7_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008009(.in0(tmp00_16_63), .in1(tmp00_17_63), .out(tmp01_8_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008010(.in0(tmp00_18_63), .in1(tmp00_19_63), .out(tmp01_9_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008011(.in0(tmp00_20_63), .in1(tmp00_21_63), .out(tmp01_10_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008012(.in0(tmp00_22_63), .in1(tmp00_23_63), .out(tmp01_11_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008013(.in0(tmp00_24_63), .in1(tmp00_25_63), .out(tmp01_12_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008014(.in0(tmp00_26_63), .in1(tmp00_27_63), .out(tmp01_13_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008015(.in0(tmp00_28_63), .in1(tmp00_29_63), .out(tmp01_14_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008016(.in0(tmp00_30_63), .in1(tmp00_31_63), .out(tmp01_15_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008017(.in0(tmp00_32_63), .in1(tmp00_33_63), .out(tmp01_16_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008018(.in0(tmp00_34_63), .in1(tmp00_35_63), .out(tmp01_17_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008019(.in0(tmp00_36_63), .in1(tmp00_37_63), .out(tmp01_18_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008020(.in0(tmp00_38_63), .in1(tmp00_39_63), .out(tmp01_19_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008021(.in0(tmp00_40_63), .in1(tmp00_41_63), .out(tmp01_20_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008022(.in0(tmp00_42_63), .in1(tmp00_43_63), .out(tmp01_21_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008023(.in0(tmp00_44_63), .in1(tmp00_45_63), .out(tmp01_22_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008024(.in0(tmp00_46_63), .in1(tmp00_47_63), .out(tmp01_23_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008025(.in0(tmp00_48_63), .in1(tmp00_49_63), .out(tmp01_24_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008026(.in0(tmp00_50_63), .in1(tmp00_51_63), .out(tmp01_25_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008027(.in0(tmp00_52_63), .in1(tmp00_53_63), .out(tmp01_26_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008028(.in0(tmp00_54_63), .in1(tmp00_55_63), .out(tmp01_27_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008029(.in0(tmp00_56_63), .in1(tmp00_57_63), .out(tmp01_28_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008030(.in0(tmp00_58_63), .in1(tmp00_59_63), .out(tmp01_29_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008031(.in0(tmp00_60_63), .in1(tmp00_61_63), .out(tmp01_30_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008032(.in0(tmp00_62_63), .in1(tmp00_63_63), .out(tmp01_31_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008033(.in0(tmp00_64_63), .in1(tmp00_65_63), .out(tmp01_32_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008034(.in0(tmp00_66_63), .in1(tmp00_67_63), .out(tmp01_33_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008035(.in0(tmp00_68_63), .in1(tmp00_69_63), .out(tmp01_34_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008036(.in0(tmp00_70_63), .in1(tmp00_71_63), .out(tmp01_35_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008037(.in0(tmp00_72_63), .in1(tmp00_73_63), .out(tmp01_36_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008038(.in0(tmp00_74_63), .in1(tmp00_75_63), .out(tmp01_37_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008039(.in0(tmp00_76_63), .in1(tmp00_77_63), .out(tmp01_38_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008040(.in0(tmp00_78_63), .in1(tmp00_79_63), .out(tmp01_39_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008041(.in0(tmp00_80_63), .in1(tmp00_81_63), .out(tmp01_40_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008042(.in0(tmp00_82_63), .in1(tmp00_83_63), .out(tmp01_41_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008043(.in0(tmp00_84_63), .in1(tmp00_85_63), .out(tmp01_42_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008044(.in0(tmp00_86_63), .in1(tmp00_87_63), .out(tmp01_43_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008045(.in0(tmp00_88_63), .in1(tmp00_89_63), .out(tmp01_44_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008046(.in0(tmp00_90_63), .in1(tmp00_91_63), .out(tmp01_45_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008047(.in0(tmp00_92_63), .in1(tmp00_93_63), .out(tmp01_46_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008048(.in0(tmp00_94_63), .in1(tmp00_95_63), .out(tmp01_47_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008049(.in0(tmp00_96_63), .in1(tmp00_97_63), .out(tmp01_48_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008050(.in0(tmp00_98_63), .in1(tmp00_99_63), .out(tmp01_49_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008051(.in0(tmp00_100_63), .in1(tmp00_101_63), .out(tmp01_50_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008052(.in0(tmp00_102_63), .in1(tmp00_103_63), .out(tmp01_51_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008053(.in0(tmp00_104_63), .in1(tmp00_105_63), .out(tmp01_52_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008054(.in0(tmp00_106_63), .in1(tmp00_107_63), .out(tmp01_53_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008055(.in0(tmp00_108_63), .in1(tmp00_109_63), .out(tmp01_54_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008056(.in0(tmp00_110_63), .in1(tmp00_111_63), .out(tmp01_55_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008057(.in0(tmp00_112_63), .in1(tmp00_113_63), .out(tmp01_56_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008058(.in0(tmp00_114_63), .in1(tmp00_115_63), .out(tmp01_57_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008059(.in0(tmp00_116_63), .in1(tmp00_117_63), .out(tmp01_58_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008060(.in0(tmp00_118_63), .in1(tmp00_119_63), .out(tmp01_59_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008061(.in0(tmp00_120_63), .in1(tmp00_121_63), .out(tmp01_60_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008062(.in0(tmp00_122_63), .in1(tmp00_123_63), .out(tmp01_61_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008063(.in0(tmp00_124_63), .in1(tmp00_125_63), .out(tmp01_62_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008064(.in0(tmp00_126_63), .in1(tmp00_127_63), .out(tmp01_63_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008065(.in0(tmp01_0_63), .in1(tmp01_1_63), .out(tmp02_0_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008066(.in0(tmp01_2_63), .in1(tmp01_3_63), .out(tmp02_1_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008067(.in0(tmp01_4_63), .in1(tmp01_5_63), .out(tmp02_2_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008068(.in0(tmp01_6_63), .in1(tmp01_7_63), .out(tmp02_3_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008069(.in0(tmp01_8_63), .in1(tmp01_9_63), .out(tmp02_4_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008070(.in0(tmp01_10_63), .in1(tmp01_11_63), .out(tmp02_5_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008071(.in0(tmp01_12_63), .in1(tmp01_13_63), .out(tmp02_6_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008072(.in0(tmp01_14_63), .in1(tmp01_15_63), .out(tmp02_7_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008073(.in0(tmp01_16_63), .in1(tmp01_17_63), .out(tmp02_8_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008074(.in0(tmp01_18_63), .in1(tmp01_19_63), .out(tmp02_9_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008075(.in0(tmp01_20_63), .in1(tmp01_21_63), .out(tmp02_10_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008076(.in0(tmp01_22_63), .in1(tmp01_23_63), .out(tmp02_11_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008077(.in0(tmp01_24_63), .in1(tmp01_25_63), .out(tmp02_12_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008078(.in0(tmp01_26_63), .in1(tmp01_27_63), .out(tmp02_13_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008079(.in0(tmp01_28_63), .in1(tmp01_29_63), .out(tmp02_14_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008080(.in0(tmp01_30_63), .in1(tmp01_31_63), .out(tmp02_15_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008081(.in0(tmp01_32_63), .in1(tmp01_33_63), .out(tmp02_16_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008082(.in0(tmp01_34_63), .in1(tmp01_35_63), .out(tmp02_17_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008083(.in0(tmp01_36_63), .in1(tmp01_37_63), .out(tmp02_18_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008084(.in0(tmp01_38_63), .in1(tmp01_39_63), .out(tmp02_19_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008085(.in0(tmp01_40_63), .in1(tmp01_41_63), .out(tmp02_20_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008086(.in0(tmp01_42_63), .in1(tmp01_43_63), .out(tmp02_21_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008087(.in0(tmp01_44_63), .in1(tmp01_45_63), .out(tmp02_22_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008088(.in0(tmp01_46_63), .in1(tmp01_47_63), .out(tmp02_23_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008089(.in0(tmp01_48_63), .in1(tmp01_49_63), .out(tmp02_24_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008090(.in0(tmp01_50_63), .in1(tmp01_51_63), .out(tmp02_25_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008091(.in0(tmp01_52_63), .in1(tmp01_53_63), .out(tmp02_26_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008092(.in0(tmp01_54_63), .in1(tmp01_55_63), .out(tmp02_27_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008093(.in0(tmp01_56_63), .in1(tmp01_57_63), .out(tmp02_28_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008094(.in0(tmp01_58_63), .in1(tmp01_59_63), .out(tmp02_29_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008095(.in0(tmp01_60_63), .in1(tmp01_61_63), .out(tmp02_30_63));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008096(.in0(tmp01_62_63), .in1(tmp01_63_63), .out(tmp02_31_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008097(.in0(tmp02_0_63), .in1(tmp02_1_63), .out(tmp03_0_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008098(.in0(tmp02_2_63), .in1(tmp02_3_63), .out(tmp03_1_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008099(.in0(tmp02_4_63), .in1(tmp02_5_63), .out(tmp03_2_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008100(.in0(tmp02_6_63), .in1(tmp02_7_63), .out(tmp03_3_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008101(.in0(tmp02_8_63), .in1(tmp02_9_63), .out(tmp03_4_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008102(.in0(tmp02_10_63), .in1(tmp02_11_63), .out(tmp03_5_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008103(.in0(tmp02_12_63), .in1(tmp02_13_63), .out(tmp03_6_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008104(.in0(tmp02_14_63), .in1(tmp02_15_63), .out(tmp03_7_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008105(.in0(tmp02_16_63), .in1(tmp02_17_63), .out(tmp03_8_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008106(.in0(tmp02_18_63), .in1(tmp02_19_63), .out(tmp03_9_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008107(.in0(tmp02_20_63), .in1(tmp02_21_63), .out(tmp03_10_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008108(.in0(tmp02_22_63), .in1(tmp02_23_63), .out(tmp03_11_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008109(.in0(tmp02_24_63), .in1(tmp02_25_63), .out(tmp03_12_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008110(.in0(tmp02_26_63), .in1(tmp02_27_63), .out(tmp03_13_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008111(.in0(tmp02_28_63), .in1(tmp02_29_63), .out(tmp03_14_63));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008112(.in0(tmp02_30_63), .in1(tmp02_31_63), .out(tmp03_15_63));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008113(.in0(tmp03_0_63), .in1(tmp03_1_63), .out(tmp04_0_63));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008114(.in0(tmp03_2_63), .in1(tmp03_3_63), .out(tmp04_1_63));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008115(.in0(tmp03_4_63), .in1(tmp03_5_63), .out(tmp04_2_63));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008116(.in0(tmp03_6_63), .in1(tmp03_7_63), .out(tmp04_3_63));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008117(.in0(tmp03_8_63), .in1(tmp03_9_63), .out(tmp04_4_63));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008118(.in0(tmp03_10_63), .in1(tmp03_11_63), .out(tmp04_5_63));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008119(.in0(tmp03_12_63), .in1(tmp03_13_63), .out(tmp04_6_63));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008120(.in0(tmp03_14_63), .in1(tmp03_15_63), .out(tmp04_7_63));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008121(.in0(tmp04_0_63), .in1(tmp04_1_63), .out(tmp05_0_63));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008122(.in0(tmp04_2_63), .in1(tmp04_3_63), .out(tmp05_1_63));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008123(.in0(tmp04_4_63), .in1(tmp04_5_63), .out(tmp05_2_63));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008124(.in0(tmp04_6_63), .in1(tmp04_7_63), .out(tmp05_3_63));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008125(.in0(tmp05_0_63), .in1(tmp05_1_63), .out(tmp06_0_63));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008126(.in0(tmp05_2_63), .in1(tmp05_3_63), .out(tmp06_1_63));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add008127(.in0(tmp06_0_63), .in1(tmp06_1_63), .out(tmp07_0_63));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008128(.in0(tmp00_0_64), .in1(tmp00_1_64), .out(tmp01_0_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008129(.in0(tmp00_2_64), .in1(tmp00_3_64), .out(tmp01_1_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008130(.in0(tmp00_4_64), .in1(tmp00_5_64), .out(tmp01_2_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008131(.in0(tmp00_6_64), .in1(tmp00_7_64), .out(tmp01_3_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008132(.in0(tmp00_8_64), .in1(tmp00_9_64), .out(tmp01_4_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008133(.in0(tmp00_10_64), .in1(tmp00_11_64), .out(tmp01_5_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008134(.in0(tmp00_12_64), .in1(tmp00_13_64), .out(tmp01_6_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008135(.in0(tmp00_14_64), .in1(tmp00_15_64), .out(tmp01_7_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008136(.in0(tmp00_16_64), .in1(tmp00_17_64), .out(tmp01_8_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008137(.in0(tmp00_18_64), .in1(tmp00_19_64), .out(tmp01_9_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008138(.in0(tmp00_20_64), .in1(tmp00_21_64), .out(tmp01_10_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008139(.in0(tmp00_22_64), .in1(tmp00_23_64), .out(tmp01_11_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008140(.in0(tmp00_24_64), .in1(tmp00_25_64), .out(tmp01_12_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008141(.in0(tmp00_26_64), .in1(tmp00_27_64), .out(tmp01_13_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008142(.in0(tmp00_28_64), .in1(tmp00_29_64), .out(tmp01_14_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008143(.in0(tmp00_30_64), .in1(tmp00_31_64), .out(tmp01_15_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008144(.in0(tmp00_32_64), .in1(tmp00_33_64), .out(tmp01_16_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008145(.in0(tmp00_34_64), .in1(tmp00_35_64), .out(tmp01_17_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008146(.in0(tmp00_36_64), .in1(tmp00_37_64), .out(tmp01_18_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008147(.in0(tmp00_38_64), .in1(tmp00_39_64), .out(tmp01_19_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008148(.in0(tmp00_40_64), .in1(tmp00_41_64), .out(tmp01_20_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008149(.in0(tmp00_42_64), .in1(tmp00_43_64), .out(tmp01_21_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008150(.in0(tmp00_44_64), .in1(tmp00_45_64), .out(tmp01_22_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008151(.in0(tmp00_46_64), .in1(tmp00_47_64), .out(tmp01_23_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008152(.in0(tmp00_48_64), .in1(tmp00_49_64), .out(tmp01_24_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008153(.in0(tmp00_50_64), .in1(tmp00_51_64), .out(tmp01_25_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008154(.in0(tmp00_52_64), .in1(tmp00_53_64), .out(tmp01_26_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008155(.in0(tmp00_54_64), .in1(tmp00_55_64), .out(tmp01_27_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008156(.in0(tmp00_56_64), .in1(tmp00_57_64), .out(tmp01_28_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008157(.in0(tmp00_58_64), .in1(tmp00_59_64), .out(tmp01_29_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008158(.in0(tmp00_60_64), .in1(tmp00_61_64), .out(tmp01_30_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008159(.in0(tmp00_62_64), .in1(tmp00_63_64), .out(tmp01_31_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008160(.in0(tmp00_64_64), .in1(tmp00_65_64), .out(tmp01_32_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008161(.in0(tmp00_66_64), .in1(tmp00_67_64), .out(tmp01_33_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008162(.in0(tmp00_68_64), .in1(tmp00_69_64), .out(tmp01_34_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008163(.in0(tmp00_70_64), .in1(tmp00_71_64), .out(tmp01_35_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008164(.in0(tmp00_72_64), .in1(tmp00_73_64), .out(tmp01_36_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008165(.in0(tmp00_74_64), .in1(tmp00_75_64), .out(tmp01_37_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008166(.in0(tmp00_76_64), .in1(tmp00_77_64), .out(tmp01_38_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008167(.in0(tmp00_78_64), .in1(tmp00_79_64), .out(tmp01_39_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008168(.in0(tmp00_80_64), .in1(tmp00_81_64), .out(tmp01_40_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008169(.in0(tmp00_82_64), .in1(tmp00_83_64), .out(tmp01_41_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008170(.in0(tmp00_84_64), .in1(tmp00_85_64), .out(tmp01_42_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008171(.in0(tmp00_86_64), .in1(tmp00_87_64), .out(tmp01_43_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008172(.in0(tmp00_88_64), .in1(tmp00_89_64), .out(tmp01_44_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008173(.in0(tmp00_90_64), .in1(tmp00_91_64), .out(tmp01_45_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008174(.in0(tmp00_92_64), .in1(tmp00_93_64), .out(tmp01_46_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008175(.in0(tmp00_94_64), .in1(tmp00_95_64), .out(tmp01_47_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008176(.in0(tmp00_96_64), .in1(tmp00_97_64), .out(tmp01_48_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008177(.in0(tmp00_98_64), .in1(tmp00_99_64), .out(tmp01_49_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008178(.in0(tmp00_100_64), .in1(tmp00_101_64), .out(tmp01_50_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008179(.in0(tmp00_102_64), .in1(tmp00_103_64), .out(tmp01_51_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008180(.in0(tmp00_104_64), .in1(tmp00_105_64), .out(tmp01_52_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008181(.in0(tmp00_106_64), .in1(tmp00_107_64), .out(tmp01_53_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008182(.in0(tmp00_108_64), .in1(tmp00_109_64), .out(tmp01_54_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008183(.in0(tmp00_110_64), .in1(tmp00_111_64), .out(tmp01_55_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008184(.in0(tmp00_112_64), .in1(tmp00_113_64), .out(tmp01_56_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008185(.in0(tmp00_114_64), .in1(tmp00_115_64), .out(tmp01_57_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008186(.in0(tmp00_116_64), .in1(tmp00_117_64), .out(tmp01_58_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008187(.in0(tmp00_118_64), .in1(tmp00_119_64), .out(tmp01_59_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008188(.in0(tmp00_120_64), .in1(tmp00_121_64), .out(tmp01_60_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008189(.in0(tmp00_122_64), .in1(tmp00_123_64), .out(tmp01_61_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008190(.in0(tmp00_124_64), .in1(tmp00_125_64), .out(tmp01_62_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008191(.in0(tmp00_126_64), .in1(tmp00_127_64), .out(tmp01_63_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008192(.in0(tmp01_0_64), .in1(tmp01_1_64), .out(tmp02_0_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008193(.in0(tmp01_2_64), .in1(tmp01_3_64), .out(tmp02_1_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008194(.in0(tmp01_4_64), .in1(tmp01_5_64), .out(tmp02_2_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008195(.in0(tmp01_6_64), .in1(tmp01_7_64), .out(tmp02_3_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008196(.in0(tmp01_8_64), .in1(tmp01_9_64), .out(tmp02_4_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008197(.in0(tmp01_10_64), .in1(tmp01_11_64), .out(tmp02_5_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008198(.in0(tmp01_12_64), .in1(tmp01_13_64), .out(tmp02_6_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008199(.in0(tmp01_14_64), .in1(tmp01_15_64), .out(tmp02_7_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008200(.in0(tmp01_16_64), .in1(tmp01_17_64), .out(tmp02_8_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008201(.in0(tmp01_18_64), .in1(tmp01_19_64), .out(tmp02_9_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008202(.in0(tmp01_20_64), .in1(tmp01_21_64), .out(tmp02_10_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008203(.in0(tmp01_22_64), .in1(tmp01_23_64), .out(tmp02_11_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008204(.in0(tmp01_24_64), .in1(tmp01_25_64), .out(tmp02_12_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008205(.in0(tmp01_26_64), .in1(tmp01_27_64), .out(tmp02_13_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008206(.in0(tmp01_28_64), .in1(tmp01_29_64), .out(tmp02_14_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008207(.in0(tmp01_30_64), .in1(tmp01_31_64), .out(tmp02_15_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008208(.in0(tmp01_32_64), .in1(tmp01_33_64), .out(tmp02_16_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008209(.in0(tmp01_34_64), .in1(tmp01_35_64), .out(tmp02_17_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008210(.in0(tmp01_36_64), .in1(tmp01_37_64), .out(tmp02_18_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008211(.in0(tmp01_38_64), .in1(tmp01_39_64), .out(tmp02_19_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008212(.in0(tmp01_40_64), .in1(tmp01_41_64), .out(tmp02_20_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008213(.in0(tmp01_42_64), .in1(tmp01_43_64), .out(tmp02_21_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008214(.in0(tmp01_44_64), .in1(tmp01_45_64), .out(tmp02_22_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008215(.in0(tmp01_46_64), .in1(tmp01_47_64), .out(tmp02_23_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008216(.in0(tmp01_48_64), .in1(tmp01_49_64), .out(tmp02_24_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008217(.in0(tmp01_50_64), .in1(tmp01_51_64), .out(tmp02_25_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008218(.in0(tmp01_52_64), .in1(tmp01_53_64), .out(tmp02_26_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008219(.in0(tmp01_54_64), .in1(tmp01_55_64), .out(tmp02_27_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008220(.in0(tmp01_56_64), .in1(tmp01_57_64), .out(tmp02_28_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008221(.in0(tmp01_58_64), .in1(tmp01_59_64), .out(tmp02_29_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008222(.in0(tmp01_60_64), .in1(tmp01_61_64), .out(tmp02_30_64));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008223(.in0(tmp01_62_64), .in1(tmp01_63_64), .out(tmp02_31_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008224(.in0(tmp02_0_64), .in1(tmp02_1_64), .out(tmp03_0_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008225(.in0(tmp02_2_64), .in1(tmp02_3_64), .out(tmp03_1_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008226(.in0(tmp02_4_64), .in1(tmp02_5_64), .out(tmp03_2_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008227(.in0(tmp02_6_64), .in1(tmp02_7_64), .out(tmp03_3_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008228(.in0(tmp02_8_64), .in1(tmp02_9_64), .out(tmp03_4_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008229(.in0(tmp02_10_64), .in1(tmp02_11_64), .out(tmp03_5_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008230(.in0(tmp02_12_64), .in1(tmp02_13_64), .out(tmp03_6_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008231(.in0(tmp02_14_64), .in1(tmp02_15_64), .out(tmp03_7_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008232(.in0(tmp02_16_64), .in1(tmp02_17_64), .out(tmp03_8_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008233(.in0(tmp02_18_64), .in1(tmp02_19_64), .out(tmp03_9_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008234(.in0(tmp02_20_64), .in1(tmp02_21_64), .out(tmp03_10_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008235(.in0(tmp02_22_64), .in1(tmp02_23_64), .out(tmp03_11_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008236(.in0(tmp02_24_64), .in1(tmp02_25_64), .out(tmp03_12_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008237(.in0(tmp02_26_64), .in1(tmp02_27_64), .out(tmp03_13_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008238(.in0(tmp02_28_64), .in1(tmp02_29_64), .out(tmp03_14_64));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008239(.in0(tmp02_30_64), .in1(tmp02_31_64), .out(tmp03_15_64));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008240(.in0(tmp03_0_64), .in1(tmp03_1_64), .out(tmp04_0_64));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008241(.in0(tmp03_2_64), .in1(tmp03_3_64), .out(tmp04_1_64));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008242(.in0(tmp03_4_64), .in1(tmp03_5_64), .out(tmp04_2_64));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008243(.in0(tmp03_6_64), .in1(tmp03_7_64), .out(tmp04_3_64));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008244(.in0(tmp03_8_64), .in1(tmp03_9_64), .out(tmp04_4_64));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008245(.in0(tmp03_10_64), .in1(tmp03_11_64), .out(tmp04_5_64));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008246(.in0(tmp03_12_64), .in1(tmp03_13_64), .out(tmp04_6_64));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008247(.in0(tmp03_14_64), .in1(tmp03_15_64), .out(tmp04_7_64));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008248(.in0(tmp04_0_64), .in1(tmp04_1_64), .out(tmp05_0_64));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008249(.in0(tmp04_2_64), .in1(tmp04_3_64), .out(tmp05_1_64));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008250(.in0(tmp04_4_64), .in1(tmp04_5_64), .out(tmp05_2_64));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008251(.in0(tmp04_6_64), .in1(tmp04_7_64), .out(tmp05_3_64));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008252(.in0(tmp05_0_64), .in1(tmp05_1_64), .out(tmp06_0_64));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008253(.in0(tmp05_2_64), .in1(tmp05_3_64), .out(tmp06_1_64));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add008254(.in0(tmp06_0_64), .in1(tmp06_1_64), .out(tmp07_0_64));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008255(.in0(tmp00_0_65), .in1(tmp00_1_65), .out(tmp01_0_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008256(.in0(tmp00_2_65), .in1(tmp00_3_65), .out(tmp01_1_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008257(.in0(tmp00_4_65), .in1(tmp00_5_65), .out(tmp01_2_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008258(.in0(tmp00_6_65), .in1(tmp00_7_65), .out(tmp01_3_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008259(.in0(tmp00_8_65), .in1(tmp00_9_65), .out(tmp01_4_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008260(.in0(tmp00_10_65), .in1(tmp00_11_65), .out(tmp01_5_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008261(.in0(tmp00_12_65), .in1(tmp00_13_65), .out(tmp01_6_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008262(.in0(tmp00_14_65), .in1(tmp00_15_65), .out(tmp01_7_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008263(.in0(tmp00_16_65), .in1(tmp00_17_65), .out(tmp01_8_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008264(.in0(tmp00_18_65), .in1(tmp00_19_65), .out(tmp01_9_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008265(.in0(tmp00_20_65), .in1(tmp00_21_65), .out(tmp01_10_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008266(.in0(tmp00_22_65), .in1(tmp00_23_65), .out(tmp01_11_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008267(.in0(tmp00_24_65), .in1(tmp00_25_65), .out(tmp01_12_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008268(.in0(tmp00_26_65), .in1(tmp00_27_65), .out(tmp01_13_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008269(.in0(tmp00_28_65), .in1(tmp00_29_65), .out(tmp01_14_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008270(.in0(tmp00_30_65), .in1(tmp00_31_65), .out(tmp01_15_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008271(.in0(tmp00_32_65), .in1(tmp00_33_65), .out(tmp01_16_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008272(.in0(tmp00_34_65), .in1(tmp00_35_65), .out(tmp01_17_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008273(.in0(tmp00_36_65), .in1(tmp00_37_65), .out(tmp01_18_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008274(.in0(tmp00_38_65), .in1(tmp00_39_65), .out(tmp01_19_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008275(.in0(tmp00_40_65), .in1(tmp00_41_65), .out(tmp01_20_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008276(.in0(tmp00_42_65), .in1(tmp00_43_65), .out(tmp01_21_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008277(.in0(tmp00_44_65), .in1(tmp00_45_65), .out(tmp01_22_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008278(.in0(tmp00_46_65), .in1(tmp00_47_65), .out(tmp01_23_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008279(.in0(tmp00_48_65), .in1(tmp00_49_65), .out(tmp01_24_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008280(.in0(tmp00_50_65), .in1(tmp00_51_65), .out(tmp01_25_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008281(.in0(tmp00_52_65), .in1(tmp00_53_65), .out(tmp01_26_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008282(.in0(tmp00_54_65), .in1(tmp00_55_65), .out(tmp01_27_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008283(.in0(tmp00_56_65), .in1(tmp00_57_65), .out(tmp01_28_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008284(.in0(tmp00_58_65), .in1(tmp00_59_65), .out(tmp01_29_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008285(.in0(tmp00_60_65), .in1(tmp00_61_65), .out(tmp01_30_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008286(.in0(tmp00_62_65), .in1(tmp00_63_65), .out(tmp01_31_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008287(.in0(tmp00_64_65), .in1(tmp00_65_65), .out(tmp01_32_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008288(.in0(tmp00_66_65), .in1(tmp00_67_65), .out(tmp01_33_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008289(.in0(tmp00_68_65), .in1(tmp00_69_65), .out(tmp01_34_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008290(.in0(tmp00_70_65), .in1(tmp00_71_65), .out(tmp01_35_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008291(.in0(tmp00_72_65), .in1(tmp00_73_65), .out(tmp01_36_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008292(.in0(tmp00_74_65), .in1(tmp00_75_65), .out(tmp01_37_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008293(.in0(tmp00_76_65), .in1(tmp00_77_65), .out(tmp01_38_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008294(.in0(tmp00_78_65), .in1(tmp00_79_65), .out(tmp01_39_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008295(.in0(tmp00_80_65), .in1(tmp00_81_65), .out(tmp01_40_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008296(.in0(tmp00_82_65), .in1(tmp00_83_65), .out(tmp01_41_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008297(.in0(tmp00_84_65), .in1(tmp00_85_65), .out(tmp01_42_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008298(.in0(tmp00_86_65), .in1(tmp00_87_65), .out(tmp01_43_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008299(.in0(tmp00_88_65), .in1(tmp00_89_65), .out(tmp01_44_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008300(.in0(tmp00_90_65), .in1(tmp00_91_65), .out(tmp01_45_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008301(.in0(tmp00_92_65), .in1(tmp00_93_65), .out(tmp01_46_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008302(.in0(tmp00_94_65), .in1(tmp00_95_65), .out(tmp01_47_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008303(.in0(tmp00_96_65), .in1(tmp00_97_65), .out(tmp01_48_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008304(.in0(tmp00_98_65), .in1(tmp00_99_65), .out(tmp01_49_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008305(.in0(tmp00_100_65), .in1(tmp00_101_65), .out(tmp01_50_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008306(.in0(tmp00_102_65), .in1(tmp00_103_65), .out(tmp01_51_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008307(.in0(tmp00_104_65), .in1(tmp00_105_65), .out(tmp01_52_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008308(.in0(tmp00_106_65), .in1(tmp00_107_65), .out(tmp01_53_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008309(.in0(tmp00_108_65), .in1(tmp00_109_65), .out(tmp01_54_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008310(.in0(tmp00_110_65), .in1(tmp00_111_65), .out(tmp01_55_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008311(.in0(tmp00_112_65), .in1(tmp00_113_65), .out(tmp01_56_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008312(.in0(tmp00_114_65), .in1(tmp00_115_65), .out(tmp01_57_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008313(.in0(tmp00_116_65), .in1(tmp00_117_65), .out(tmp01_58_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008314(.in0(tmp00_118_65), .in1(tmp00_119_65), .out(tmp01_59_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008315(.in0(tmp00_120_65), .in1(tmp00_121_65), .out(tmp01_60_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008316(.in0(tmp00_122_65), .in1(tmp00_123_65), .out(tmp01_61_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008317(.in0(tmp00_124_65), .in1(tmp00_125_65), .out(tmp01_62_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008318(.in0(tmp00_126_65), .in1(tmp00_127_65), .out(tmp01_63_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008319(.in0(tmp01_0_65), .in1(tmp01_1_65), .out(tmp02_0_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008320(.in0(tmp01_2_65), .in1(tmp01_3_65), .out(tmp02_1_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008321(.in0(tmp01_4_65), .in1(tmp01_5_65), .out(tmp02_2_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008322(.in0(tmp01_6_65), .in1(tmp01_7_65), .out(tmp02_3_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008323(.in0(tmp01_8_65), .in1(tmp01_9_65), .out(tmp02_4_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008324(.in0(tmp01_10_65), .in1(tmp01_11_65), .out(tmp02_5_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008325(.in0(tmp01_12_65), .in1(tmp01_13_65), .out(tmp02_6_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008326(.in0(tmp01_14_65), .in1(tmp01_15_65), .out(tmp02_7_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008327(.in0(tmp01_16_65), .in1(tmp01_17_65), .out(tmp02_8_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008328(.in0(tmp01_18_65), .in1(tmp01_19_65), .out(tmp02_9_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008329(.in0(tmp01_20_65), .in1(tmp01_21_65), .out(tmp02_10_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008330(.in0(tmp01_22_65), .in1(tmp01_23_65), .out(tmp02_11_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008331(.in0(tmp01_24_65), .in1(tmp01_25_65), .out(tmp02_12_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008332(.in0(tmp01_26_65), .in1(tmp01_27_65), .out(tmp02_13_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008333(.in0(tmp01_28_65), .in1(tmp01_29_65), .out(tmp02_14_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008334(.in0(tmp01_30_65), .in1(tmp01_31_65), .out(tmp02_15_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008335(.in0(tmp01_32_65), .in1(tmp01_33_65), .out(tmp02_16_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008336(.in0(tmp01_34_65), .in1(tmp01_35_65), .out(tmp02_17_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008337(.in0(tmp01_36_65), .in1(tmp01_37_65), .out(tmp02_18_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008338(.in0(tmp01_38_65), .in1(tmp01_39_65), .out(tmp02_19_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008339(.in0(tmp01_40_65), .in1(tmp01_41_65), .out(tmp02_20_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008340(.in0(tmp01_42_65), .in1(tmp01_43_65), .out(tmp02_21_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008341(.in0(tmp01_44_65), .in1(tmp01_45_65), .out(tmp02_22_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008342(.in0(tmp01_46_65), .in1(tmp01_47_65), .out(tmp02_23_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008343(.in0(tmp01_48_65), .in1(tmp01_49_65), .out(tmp02_24_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008344(.in0(tmp01_50_65), .in1(tmp01_51_65), .out(tmp02_25_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008345(.in0(tmp01_52_65), .in1(tmp01_53_65), .out(tmp02_26_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008346(.in0(tmp01_54_65), .in1(tmp01_55_65), .out(tmp02_27_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008347(.in0(tmp01_56_65), .in1(tmp01_57_65), .out(tmp02_28_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008348(.in0(tmp01_58_65), .in1(tmp01_59_65), .out(tmp02_29_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008349(.in0(tmp01_60_65), .in1(tmp01_61_65), .out(tmp02_30_65));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008350(.in0(tmp01_62_65), .in1(tmp01_63_65), .out(tmp02_31_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008351(.in0(tmp02_0_65), .in1(tmp02_1_65), .out(tmp03_0_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008352(.in0(tmp02_2_65), .in1(tmp02_3_65), .out(tmp03_1_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008353(.in0(tmp02_4_65), .in1(tmp02_5_65), .out(tmp03_2_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008354(.in0(tmp02_6_65), .in1(tmp02_7_65), .out(tmp03_3_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008355(.in0(tmp02_8_65), .in1(tmp02_9_65), .out(tmp03_4_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008356(.in0(tmp02_10_65), .in1(tmp02_11_65), .out(tmp03_5_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008357(.in0(tmp02_12_65), .in1(tmp02_13_65), .out(tmp03_6_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008358(.in0(tmp02_14_65), .in1(tmp02_15_65), .out(tmp03_7_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008359(.in0(tmp02_16_65), .in1(tmp02_17_65), .out(tmp03_8_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008360(.in0(tmp02_18_65), .in1(tmp02_19_65), .out(tmp03_9_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008361(.in0(tmp02_20_65), .in1(tmp02_21_65), .out(tmp03_10_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008362(.in0(tmp02_22_65), .in1(tmp02_23_65), .out(tmp03_11_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008363(.in0(tmp02_24_65), .in1(tmp02_25_65), .out(tmp03_12_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008364(.in0(tmp02_26_65), .in1(tmp02_27_65), .out(tmp03_13_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008365(.in0(tmp02_28_65), .in1(tmp02_29_65), .out(tmp03_14_65));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008366(.in0(tmp02_30_65), .in1(tmp02_31_65), .out(tmp03_15_65));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008367(.in0(tmp03_0_65), .in1(tmp03_1_65), .out(tmp04_0_65));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008368(.in0(tmp03_2_65), .in1(tmp03_3_65), .out(tmp04_1_65));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008369(.in0(tmp03_4_65), .in1(tmp03_5_65), .out(tmp04_2_65));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008370(.in0(tmp03_6_65), .in1(tmp03_7_65), .out(tmp04_3_65));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008371(.in0(tmp03_8_65), .in1(tmp03_9_65), .out(tmp04_4_65));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008372(.in0(tmp03_10_65), .in1(tmp03_11_65), .out(tmp04_5_65));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008373(.in0(tmp03_12_65), .in1(tmp03_13_65), .out(tmp04_6_65));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008374(.in0(tmp03_14_65), .in1(tmp03_15_65), .out(tmp04_7_65));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008375(.in0(tmp04_0_65), .in1(tmp04_1_65), .out(tmp05_0_65));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008376(.in0(tmp04_2_65), .in1(tmp04_3_65), .out(tmp05_1_65));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008377(.in0(tmp04_4_65), .in1(tmp04_5_65), .out(tmp05_2_65));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008378(.in0(tmp04_6_65), .in1(tmp04_7_65), .out(tmp05_3_65));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008379(.in0(tmp05_0_65), .in1(tmp05_1_65), .out(tmp06_0_65));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008380(.in0(tmp05_2_65), .in1(tmp05_3_65), .out(tmp06_1_65));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add008381(.in0(tmp06_0_65), .in1(tmp06_1_65), .out(tmp07_0_65));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008382(.in0(tmp00_0_66), .in1(tmp00_1_66), .out(tmp01_0_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008383(.in0(tmp00_2_66), .in1(tmp00_3_66), .out(tmp01_1_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008384(.in0(tmp00_4_66), .in1(tmp00_5_66), .out(tmp01_2_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008385(.in0(tmp00_6_66), .in1(tmp00_7_66), .out(tmp01_3_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008386(.in0(tmp00_8_66), .in1(tmp00_9_66), .out(tmp01_4_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008387(.in0(tmp00_10_66), .in1(tmp00_11_66), .out(tmp01_5_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008388(.in0(tmp00_12_66), .in1(tmp00_13_66), .out(tmp01_6_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008389(.in0(tmp00_14_66), .in1(tmp00_15_66), .out(tmp01_7_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008390(.in0(tmp00_16_66), .in1(tmp00_17_66), .out(tmp01_8_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008391(.in0(tmp00_18_66), .in1(tmp00_19_66), .out(tmp01_9_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008392(.in0(tmp00_20_66), .in1(tmp00_21_66), .out(tmp01_10_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008393(.in0(tmp00_22_66), .in1(tmp00_23_66), .out(tmp01_11_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008394(.in0(tmp00_24_66), .in1(tmp00_25_66), .out(tmp01_12_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008395(.in0(tmp00_26_66), .in1(tmp00_27_66), .out(tmp01_13_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008396(.in0(tmp00_28_66), .in1(tmp00_29_66), .out(tmp01_14_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008397(.in0(tmp00_30_66), .in1(tmp00_31_66), .out(tmp01_15_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008398(.in0(tmp00_32_66), .in1(tmp00_33_66), .out(tmp01_16_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008399(.in0(tmp00_34_66), .in1(tmp00_35_66), .out(tmp01_17_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008400(.in0(tmp00_36_66), .in1(tmp00_37_66), .out(tmp01_18_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008401(.in0(tmp00_38_66), .in1(tmp00_39_66), .out(tmp01_19_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008402(.in0(tmp00_40_66), .in1(tmp00_41_66), .out(tmp01_20_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008403(.in0(tmp00_42_66), .in1(tmp00_43_66), .out(tmp01_21_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008404(.in0(tmp00_44_66), .in1(tmp00_45_66), .out(tmp01_22_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008405(.in0(tmp00_46_66), .in1(tmp00_47_66), .out(tmp01_23_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008406(.in0(tmp00_48_66), .in1(tmp00_49_66), .out(tmp01_24_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008407(.in0(tmp00_50_66), .in1(tmp00_51_66), .out(tmp01_25_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008408(.in0(tmp00_52_66), .in1(tmp00_53_66), .out(tmp01_26_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008409(.in0(tmp00_54_66), .in1(tmp00_55_66), .out(tmp01_27_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008410(.in0(tmp00_56_66), .in1(tmp00_57_66), .out(tmp01_28_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008411(.in0(tmp00_58_66), .in1(tmp00_59_66), .out(tmp01_29_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008412(.in0(tmp00_60_66), .in1(tmp00_61_66), .out(tmp01_30_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008413(.in0(tmp00_62_66), .in1(tmp00_63_66), .out(tmp01_31_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008414(.in0(tmp00_64_66), .in1(tmp00_65_66), .out(tmp01_32_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008415(.in0(tmp00_66_66), .in1(tmp00_67_66), .out(tmp01_33_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008416(.in0(tmp00_68_66), .in1(tmp00_69_66), .out(tmp01_34_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008417(.in0(tmp00_70_66), .in1(tmp00_71_66), .out(tmp01_35_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008418(.in0(tmp00_72_66), .in1(tmp00_73_66), .out(tmp01_36_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008419(.in0(tmp00_74_66), .in1(tmp00_75_66), .out(tmp01_37_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008420(.in0(tmp00_76_66), .in1(tmp00_77_66), .out(tmp01_38_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008421(.in0(tmp00_78_66), .in1(tmp00_79_66), .out(tmp01_39_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008422(.in0(tmp00_80_66), .in1(tmp00_81_66), .out(tmp01_40_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008423(.in0(tmp00_82_66), .in1(tmp00_83_66), .out(tmp01_41_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008424(.in0(tmp00_84_66), .in1(tmp00_85_66), .out(tmp01_42_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008425(.in0(tmp00_86_66), .in1(tmp00_87_66), .out(tmp01_43_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008426(.in0(tmp00_88_66), .in1(tmp00_89_66), .out(tmp01_44_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008427(.in0(tmp00_90_66), .in1(tmp00_91_66), .out(tmp01_45_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008428(.in0(tmp00_92_66), .in1(tmp00_93_66), .out(tmp01_46_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008429(.in0(tmp00_94_66), .in1(tmp00_95_66), .out(tmp01_47_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008430(.in0(tmp00_96_66), .in1(tmp00_97_66), .out(tmp01_48_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008431(.in0(tmp00_98_66), .in1(tmp00_99_66), .out(tmp01_49_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008432(.in0(tmp00_100_66), .in1(tmp00_101_66), .out(tmp01_50_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008433(.in0(tmp00_102_66), .in1(tmp00_103_66), .out(tmp01_51_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008434(.in0(tmp00_104_66), .in1(tmp00_105_66), .out(tmp01_52_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008435(.in0(tmp00_106_66), .in1(tmp00_107_66), .out(tmp01_53_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008436(.in0(tmp00_108_66), .in1(tmp00_109_66), .out(tmp01_54_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008437(.in0(tmp00_110_66), .in1(tmp00_111_66), .out(tmp01_55_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008438(.in0(tmp00_112_66), .in1(tmp00_113_66), .out(tmp01_56_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008439(.in0(tmp00_114_66), .in1(tmp00_115_66), .out(tmp01_57_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008440(.in0(tmp00_116_66), .in1(tmp00_117_66), .out(tmp01_58_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008441(.in0(tmp00_118_66), .in1(tmp00_119_66), .out(tmp01_59_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008442(.in0(tmp00_120_66), .in1(tmp00_121_66), .out(tmp01_60_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008443(.in0(tmp00_122_66), .in1(tmp00_123_66), .out(tmp01_61_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008444(.in0(tmp00_124_66), .in1(tmp00_125_66), .out(tmp01_62_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008445(.in0(tmp00_126_66), .in1(tmp00_127_66), .out(tmp01_63_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008446(.in0(tmp01_0_66), .in1(tmp01_1_66), .out(tmp02_0_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008447(.in0(tmp01_2_66), .in1(tmp01_3_66), .out(tmp02_1_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008448(.in0(tmp01_4_66), .in1(tmp01_5_66), .out(tmp02_2_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008449(.in0(tmp01_6_66), .in1(tmp01_7_66), .out(tmp02_3_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008450(.in0(tmp01_8_66), .in1(tmp01_9_66), .out(tmp02_4_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008451(.in0(tmp01_10_66), .in1(tmp01_11_66), .out(tmp02_5_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008452(.in0(tmp01_12_66), .in1(tmp01_13_66), .out(tmp02_6_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008453(.in0(tmp01_14_66), .in1(tmp01_15_66), .out(tmp02_7_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008454(.in0(tmp01_16_66), .in1(tmp01_17_66), .out(tmp02_8_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008455(.in0(tmp01_18_66), .in1(tmp01_19_66), .out(tmp02_9_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008456(.in0(tmp01_20_66), .in1(tmp01_21_66), .out(tmp02_10_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008457(.in0(tmp01_22_66), .in1(tmp01_23_66), .out(tmp02_11_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008458(.in0(tmp01_24_66), .in1(tmp01_25_66), .out(tmp02_12_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008459(.in0(tmp01_26_66), .in1(tmp01_27_66), .out(tmp02_13_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008460(.in0(tmp01_28_66), .in1(tmp01_29_66), .out(tmp02_14_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008461(.in0(tmp01_30_66), .in1(tmp01_31_66), .out(tmp02_15_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008462(.in0(tmp01_32_66), .in1(tmp01_33_66), .out(tmp02_16_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008463(.in0(tmp01_34_66), .in1(tmp01_35_66), .out(tmp02_17_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008464(.in0(tmp01_36_66), .in1(tmp01_37_66), .out(tmp02_18_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008465(.in0(tmp01_38_66), .in1(tmp01_39_66), .out(tmp02_19_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008466(.in0(tmp01_40_66), .in1(tmp01_41_66), .out(tmp02_20_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008467(.in0(tmp01_42_66), .in1(tmp01_43_66), .out(tmp02_21_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008468(.in0(tmp01_44_66), .in1(tmp01_45_66), .out(tmp02_22_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008469(.in0(tmp01_46_66), .in1(tmp01_47_66), .out(tmp02_23_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008470(.in0(tmp01_48_66), .in1(tmp01_49_66), .out(tmp02_24_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008471(.in0(tmp01_50_66), .in1(tmp01_51_66), .out(tmp02_25_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008472(.in0(tmp01_52_66), .in1(tmp01_53_66), .out(tmp02_26_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008473(.in0(tmp01_54_66), .in1(tmp01_55_66), .out(tmp02_27_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008474(.in0(tmp01_56_66), .in1(tmp01_57_66), .out(tmp02_28_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008475(.in0(tmp01_58_66), .in1(tmp01_59_66), .out(tmp02_29_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008476(.in0(tmp01_60_66), .in1(tmp01_61_66), .out(tmp02_30_66));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008477(.in0(tmp01_62_66), .in1(tmp01_63_66), .out(tmp02_31_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008478(.in0(tmp02_0_66), .in1(tmp02_1_66), .out(tmp03_0_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008479(.in0(tmp02_2_66), .in1(tmp02_3_66), .out(tmp03_1_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008480(.in0(tmp02_4_66), .in1(tmp02_5_66), .out(tmp03_2_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008481(.in0(tmp02_6_66), .in1(tmp02_7_66), .out(tmp03_3_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008482(.in0(tmp02_8_66), .in1(tmp02_9_66), .out(tmp03_4_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008483(.in0(tmp02_10_66), .in1(tmp02_11_66), .out(tmp03_5_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008484(.in0(tmp02_12_66), .in1(tmp02_13_66), .out(tmp03_6_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008485(.in0(tmp02_14_66), .in1(tmp02_15_66), .out(tmp03_7_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008486(.in0(tmp02_16_66), .in1(tmp02_17_66), .out(tmp03_8_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008487(.in0(tmp02_18_66), .in1(tmp02_19_66), .out(tmp03_9_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008488(.in0(tmp02_20_66), .in1(tmp02_21_66), .out(tmp03_10_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008489(.in0(tmp02_22_66), .in1(tmp02_23_66), .out(tmp03_11_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008490(.in0(tmp02_24_66), .in1(tmp02_25_66), .out(tmp03_12_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008491(.in0(tmp02_26_66), .in1(tmp02_27_66), .out(tmp03_13_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008492(.in0(tmp02_28_66), .in1(tmp02_29_66), .out(tmp03_14_66));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008493(.in0(tmp02_30_66), .in1(tmp02_31_66), .out(tmp03_15_66));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008494(.in0(tmp03_0_66), .in1(tmp03_1_66), .out(tmp04_0_66));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008495(.in0(tmp03_2_66), .in1(tmp03_3_66), .out(tmp04_1_66));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008496(.in0(tmp03_4_66), .in1(tmp03_5_66), .out(tmp04_2_66));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008497(.in0(tmp03_6_66), .in1(tmp03_7_66), .out(tmp04_3_66));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008498(.in0(tmp03_8_66), .in1(tmp03_9_66), .out(tmp04_4_66));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008499(.in0(tmp03_10_66), .in1(tmp03_11_66), .out(tmp04_5_66));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008500(.in0(tmp03_12_66), .in1(tmp03_13_66), .out(tmp04_6_66));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008501(.in0(tmp03_14_66), .in1(tmp03_15_66), .out(tmp04_7_66));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008502(.in0(tmp04_0_66), .in1(tmp04_1_66), .out(tmp05_0_66));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008503(.in0(tmp04_2_66), .in1(tmp04_3_66), .out(tmp05_1_66));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008504(.in0(tmp04_4_66), .in1(tmp04_5_66), .out(tmp05_2_66));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008505(.in0(tmp04_6_66), .in1(tmp04_7_66), .out(tmp05_3_66));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008506(.in0(tmp05_0_66), .in1(tmp05_1_66), .out(tmp06_0_66));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008507(.in0(tmp05_2_66), .in1(tmp05_3_66), .out(tmp06_1_66));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add008508(.in0(tmp06_0_66), .in1(tmp06_1_66), .out(tmp07_0_66));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008509(.in0(tmp00_0_67), .in1(tmp00_1_67), .out(tmp01_0_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008510(.in0(tmp00_2_67), .in1(tmp00_3_67), .out(tmp01_1_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008511(.in0(tmp00_4_67), .in1(tmp00_5_67), .out(tmp01_2_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008512(.in0(tmp00_6_67), .in1(tmp00_7_67), .out(tmp01_3_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008513(.in0(tmp00_8_67), .in1(tmp00_9_67), .out(tmp01_4_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008514(.in0(tmp00_10_67), .in1(tmp00_11_67), .out(tmp01_5_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008515(.in0(tmp00_12_67), .in1(tmp00_13_67), .out(tmp01_6_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008516(.in0(tmp00_14_67), .in1(tmp00_15_67), .out(tmp01_7_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008517(.in0(tmp00_16_67), .in1(tmp00_17_67), .out(tmp01_8_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008518(.in0(tmp00_18_67), .in1(tmp00_19_67), .out(tmp01_9_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008519(.in0(tmp00_20_67), .in1(tmp00_21_67), .out(tmp01_10_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008520(.in0(tmp00_22_67), .in1(tmp00_23_67), .out(tmp01_11_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008521(.in0(tmp00_24_67), .in1(tmp00_25_67), .out(tmp01_12_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008522(.in0(tmp00_26_67), .in1(tmp00_27_67), .out(tmp01_13_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008523(.in0(tmp00_28_67), .in1(tmp00_29_67), .out(tmp01_14_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008524(.in0(tmp00_30_67), .in1(tmp00_31_67), .out(tmp01_15_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008525(.in0(tmp00_32_67), .in1(tmp00_33_67), .out(tmp01_16_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008526(.in0(tmp00_34_67), .in1(tmp00_35_67), .out(tmp01_17_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008527(.in0(tmp00_36_67), .in1(tmp00_37_67), .out(tmp01_18_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008528(.in0(tmp00_38_67), .in1(tmp00_39_67), .out(tmp01_19_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008529(.in0(tmp00_40_67), .in1(tmp00_41_67), .out(tmp01_20_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008530(.in0(tmp00_42_67), .in1(tmp00_43_67), .out(tmp01_21_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008531(.in0(tmp00_44_67), .in1(tmp00_45_67), .out(tmp01_22_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008532(.in0(tmp00_46_67), .in1(tmp00_47_67), .out(tmp01_23_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008533(.in0(tmp00_48_67), .in1(tmp00_49_67), .out(tmp01_24_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008534(.in0(tmp00_50_67), .in1(tmp00_51_67), .out(tmp01_25_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008535(.in0(tmp00_52_67), .in1(tmp00_53_67), .out(tmp01_26_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008536(.in0(tmp00_54_67), .in1(tmp00_55_67), .out(tmp01_27_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008537(.in0(tmp00_56_67), .in1(tmp00_57_67), .out(tmp01_28_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008538(.in0(tmp00_58_67), .in1(tmp00_59_67), .out(tmp01_29_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008539(.in0(tmp00_60_67), .in1(tmp00_61_67), .out(tmp01_30_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008540(.in0(tmp00_62_67), .in1(tmp00_63_67), .out(tmp01_31_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008541(.in0(tmp00_64_67), .in1(tmp00_65_67), .out(tmp01_32_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008542(.in0(tmp00_66_67), .in1(tmp00_67_67), .out(tmp01_33_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008543(.in0(tmp00_68_67), .in1(tmp00_69_67), .out(tmp01_34_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008544(.in0(tmp00_70_67), .in1(tmp00_71_67), .out(tmp01_35_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008545(.in0(tmp00_72_67), .in1(tmp00_73_67), .out(tmp01_36_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008546(.in0(tmp00_74_67), .in1(tmp00_75_67), .out(tmp01_37_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008547(.in0(tmp00_76_67), .in1(tmp00_77_67), .out(tmp01_38_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008548(.in0(tmp00_78_67), .in1(tmp00_79_67), .out(tmp01_39_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008549(.in0(tmp00_80_67), .in1(tmp00_81_67), .out(tmp01_40_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008550(.in0(tmp00_82_67), .in1(tmp00_83_67), .out(tmp01_41_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008551(.in0(tmp00_84_67), .in1(tmp00_85_67), .out(tmp01_42_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008552(.in0(tmp00_86_67), .in1(tmp00_87_67), .out(tmp01_43_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008553(.in0(tmp00_88_67), .in1(tmp00_89_67), .out(tmp01_44_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008554(.in0(tmp00_90_67), .in1(tmp00_91_67), .out(tmp01_45_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008555(.in0(tmp00_92_67), .in1(tmp00_93_67), .out(tmp01_46_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008556(.in0(tmp00_94_67), .in1(tmp00_95_67), .out(tmp01_47_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008557(.in0(tmp00_96_67), .in1(tmp00_97_67), .out(tmp01_48_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008558(.in0(tmp00_98_67), .in1(tmp00_99_67), .out(tmp01_49_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008559(.in0(tmp00_100_67), .in1(tmp00_101_67), .out(tmp01_50_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008560(.in0(tmp00_102_67), .in1(tmp00_103_67), .out(tmp01_51_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008561(.in0(tmp00_104_67), .in1(tmp00_105_67), .out(tmp01_52_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008562(.in0(tmp00_106_67), .in1(tmp00_107_67), .out(tmp01_53_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008563(.in0(tmp00_108_67), .in1(tmp00_109_67), .out(tmp01_54_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008564(.in0(tmp00_110_67), .in1(tmp00_111_67), .out(tmp01_55_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008565(.in0(tmp00_112_67), .in1(tmp00_113_67), .out(tmp01_56_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008566(.in0(tmp00_114_67), .in1(tmp00_115_67), .out(tmp01_57_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008567(.in0(tmp00_116_67), .in1(tmp00_117_67), .out(tmp01_58_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008568(.in0(tmp00_118_67), .in1(tmp00_119_67), .out(tmp01_59_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008569(.in0(tmp00_120_67), .in1(tmp00_121_67), .out(tmp01_60_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008570(.in0(tmp00_122_67), .in1(tmp00_123_67), .out(tmp01_61_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008571(.in0(tmp00_124_67), .in1(tmp00_125_67), .out(tmp01_62_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008572(.in0(tmp00_126_67), .in1(tmp00_127_67), .out(tmp01_63_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008573(.in0(tmp01_0_67), .in1(tmp01_1_67), .out(tmp02_0_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008574(.in0(tmp01_2_67), .in1(tmp01_3_67), .out(tmp02_1_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008575(.in0(tmp01_4_67), .in1(tmp01_5_67), .out(tmp02_2_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008576(.in0(tmp01_6_67), .in1(tmp01_7_67), .out(tmp02_3_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008577(.in0(tmp01_8_67), .in1(tmp01_9_67), .out(tmp02_4_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008578(.in0(tmp01_10_67), .in1(tmp01_11_67), .out(tmp02_5_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008579(.in0(tmp01_12_67), .in1(tmp01_13_67), .out(tmp02_6_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008580(.in0(tmp01_14_67), .in1(tmp01_15_67), .out(tmp02_7_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008581(.in0(tmp01_16_67), .in1(tmp01_17_67), .out(tmp02_8_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008582(.in0(tmp01_18_67), .in1(tmp01_19_67), .out(tmp02_9_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008583(.in0(tmp01_20_67), .in1(tmp01_21_67), .out(tmp02_10_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008584(.in0(tmp01_22_67), .in1(tmp01_23_67), .out(tmp02_11_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008585(.in0(tmp01_24_67), .in1(tmp01_25_67), .out(tmp02_12_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008586(.in0(tmp01_26_67), .in1(tmp01_27_67), .out(tmp02_13_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008587(.in0(tmp01_28_67), .in1(tmp01_29_67), .out(tmp02_14_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008588(.in0(tmp01_30_67), .in1(tmp01_31_67), .out(tmp02_15_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008589(.in0(tmp01_32_67), .in1(tmp01_33_67), .out(tmp02_16_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008590(.in0(tmp01_34_67), .in1(tmp01_35_67), .out(tmp02_17_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008591(.in0(tmp01_36_67), .in1(tmp01_37_67), .out(tmp02_18_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008592(.in0(tmp01_38_67), .in1(tmp01_39_67), .out(tmp02_19_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008593(.in0(tmp01_40_67), .in1(tmp01_41_67), .out(tmp02_20_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008594(.in0(tmp01_42_67), .in1(tmp01_43_67), .out(tmp02_21_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008595(.in0(tmp01_44_67), .in1(tmp01_45_67), .out(tmp02_22_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008596(.in0(tmp01_46_67), .in1(tmp01_47_67), .out(tmp02_23_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008597(.in0(tmp01_48_67), .in1(tmp01_49_67), .out(tmp02_24_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008598(.in0(tmp01_50_67), .in1(tmp01_51_67), .out(tmp02_25_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008599(.in0(tmp01_52_67), .in1(tmp01_53_67), .out(tmp02_26_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008600(.in0(tmp01_54_67), .in1(tmp01_55_67), .out(tmp02_27_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008601(.in0(tmp01_56_67), .in1(tmp01_57_67), .out(tmp02_28_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008602(.in0(tmp01_58_67), .in1(tmp01_59_67), .out(tmp02_29_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008603(.in0(tmp01_60_67), .in1(tmp01_61_67), .out(tmp02_30_67));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008604(.in0(tmp01_62_67), .in1(tmp01_63_67), .out(tmp02_31_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008605(.in0(tmp02_0_67), .in1(tmp02_1_67), .out(tmp03_0_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008606(.in0(tmp02_2_67), .in1(tmp02_3_67), .out(tmp03_1_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008607(.in0(tmp02_4_67), .in1(tmp02_5_67), .out(tmp03_2_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008608(.in0(tmp02_6_67), .in1(tmp02_7_67), .out(tmp03_3_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008609(.in0(tmp02_8_67), .in1(tmp02_9_67), .out(tmp03_4_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008610(.in0(tmp02_10_67), .in1(tmp02_11_67), .out(tmp03_5_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008611(.in0(tmp02_12_67), .in1(tmp02_13_67), .out(tmp03_6_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008612(.in0(tmp02_14_67), .in1(tmp02_15_67), .out(tmp03_7_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008613(.in0(tmp02_16_67), .in1(tmp02_17_67), .out(tmp03_8_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008614(.in0(tmp02_18_67), .in1(tmp02_19_67), .out(tmp03_9_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008615(.in0(tmp02_20_67), .in1(tmp02_21_67), .out(tmp03_10_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008616(.in0(tmp02_22_67), .in1(tmp02_23_67), .out(tmp03_11_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008617(.in0(tmp02_24_67), .in1(tmp02_25_67), .out(tmp03_12_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008618(.in0(tmp02_26_67), .in1(tmp02_27_67), .out(tmp03_13_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008619(.in0(tmp02_28_67), .in1(tmp02_29_67), .out(tmp03_14_67));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008620(.in0(tmp02_30_67), .in1(tmp02_31_67), .out(tmp03_15_67));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008621(.in0(tmp03_0_67), .in1(tmp03_1_67), .out(tmp04_0_67));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008622(.in0(tmp03_2_67), .in1(tmp03_3_67), .out(tmp04_1_67));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008623(.in0(tmp03_4_67), .in1(tmp03_5_67), .out(tmp04_2_67));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008624(.in0(tmp03_6_67), .in1(tmp03_7_67), .out(tmp04_3_67));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008625(.in0(tmp03_8_67), .in1(tmp03_9_67), .out(tmp04_4_67));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008626(.in0(tmp03_10_67), .in1(tmp03_11_67), .out(tmp04_5_67));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008627(.in0(tmp03_12_67), .in1(tmp03_13_67), .out(tmp04_6_67));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008628(.in0(tmp03_14_67), .in1(tmp03_15_67), .out(tmp04_7_67));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008629(.in0(tmp04_0_67), .in1(tmp04_1_67), .out(tmp05_0_67));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008630(.in0(tmp04_2_67), .in1(tmp04_3_67), .out(tmp05_1_67));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008631(.in0(tmp04_4_67), .in1(tmp04_5_67), .out(tmp05_2_67));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008632(.in0(tmp04_6_67), .in1(tmp04_7_67), .out(tmp05_3_67));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008633(.in0(tmp05_0_67), .in1(tmp05_1_67), .out(tmp06_0_67));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008634(.in0(tmp05_2_67), .in1(tmp05_3_67), .out(tmp06_1_67));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add008635(.in0(tmp06_0_67), .in1(tmp06_1_67), .out(tmp07_0_67));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008636(.in0(tmp00_0_68), .in1(tmp00_1_68), .out(tmp01_0_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008637(.in0(tmp00_2_68), .in1(tmp00_3_68), .out(tmp01_1_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008638(.in0(tmp00_4_68), .in1(tmp00_5_68), .out(tmp01_2_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008639(.in0(tmp00_6_68), .in1(tmp00_7_68), .out(tmp01_3_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008640(.in0(tmp00_8_68), .in1(tmp00_9_68), .out(tmp01_4_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008641(.in0(tmp00_10_68), .in1(tmp00_11_68), .out(tmp01_5_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008642(.in0(tmp00_12_68), .in1(tmp00_13_68), .out(tmp01_6_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008643(.in0(tmp00_14_68), .in1(tmp00_15_68), .out(tmp01_7_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008644(.in0(tmp00_16_68), .in1(tmp00_17_68), .out(tmp01_8_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008645(.in0(tmp00_18_68), .in1(tmp00_19_68), .out(tmp01_9_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008646(.in0(tmp00_20_68), .in1(tmp00_21_68), .out(tmp01_10_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008647(.in0(tmp00_22_68), .in1(tmp00_23_68), .out(tmp01_11_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008648(.in0(tmp00_24_68), .in1(tmp00_25_68), .out(tmp01_12_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008649(.in0(tmp00_26_68), .in1(tmp00_27_68), .out(tmp01_13_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008650(.in0(tmp00_28_68), .in1(tmp00_29_68), .out(tmp01_14_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008651(.in0(tmp00_30_68), .in1(tmp00_31_68), .out(tmp01_15_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008652(.in0(tmp00_32_68), .in1(tmp00_33_68), .out(tmp01_16_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008653(.in0(tmp00_34_68), .in1(tmp00_35_68), .out(tmp01_17_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008654(.in0(tmp00_36_68), .in1(tmp00_37_68), .out(tmp01_18_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008655(.in0(tmp00_38_68), .in1(tmp00_39_68), .out(tmp01_19_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008656(.in0(tmp00_40_68), .in1(tmp00_41_68), .out(tmp01_20_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008657(.in0(tmp00_42_68), .in1(tmp00_43_68), .out(tmp01_21_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008658(.in0(tmp00_44_68), .in1(tmp00_45_68), .out(tmp01_22_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008659(.in0(tmp00_46_68), .in1(tmp00_47_68), .out(tmp01_23_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008660(.in0(tmp00_48_68), .in1(tmp00_49_68), .out(tmp01_24_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008661(.in0(tmp00_50_68), .in1(tmp00_51_68), .out(tmp01_25_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008662(.in0(tmp00_52_68), .in1(tmp00_53_68), .out(tmp01_26_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008663(.in0(tmp00_54_68), .in1(tmp00_55_68), .out(tmp01_27_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008664(.in0(tmp00_56_68), .in1(tmp00_57_68), .out(tmp01_28_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008665(.in0(tmp00_58_68), .in1(tmp00_59_68), .out(tmp01_29_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008666(.in0(tmp00_60_68), .in1(tmp00_61_68), .out(tmp01_30_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008667(.in0(tmp00_62_68), .in1(tmp00_63_68), .out(tmp01_31_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008668(.in0(tmp00_64_68), .in1(tmp00_65_68), .out(tmp01_32_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008669(.in0(tmp00_66_68), .in1(tmp00_67_68), .out(tmp01_33_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008670(.in0(tmp00_68_68), .in1(tmp00_69_68), .out(tmp01_34_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008671(.in0(tmp00_70_68), .in1(tmp00_71_68), .out(tmp01_35_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008672(.in0(tmp00_72_68), .in1(tmp00_73_68), .out(tmp01_36_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008673(.in0(tmp00_74_68), .in1(tmp00_75_68), .out(tmp01_37_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008674(.in0(tmp00_76_68), .in1(tmp00_77_68), .out(tmp01_38_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008675(.in0(tmp00_78_68), .in1(tmp00_79_68), .out(tmp01_39_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008676(.in0(tmp00_80_68), .in1(tmp00_81_68), .out(tmp01_40_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008677(.in0(tmp00_82_68), .in1(tmp00_83_68), .out(tmp01_41_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008678(.in0(tmp00_84_68), .in1(tmp00_85_68), .out(tmp01_42_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008679(.in0(tmp00_86_68), .in1(tmp00_87_68), .out(tmp01_43_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008680(.in0(tmp00_88_68), .in1(tmp00_89_68), .out(tmp01_44_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008681(.in0(tmp00_90_68), .in1(tmp00_91_68), .out(tmp01_45_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008682(.in0(tmp00_92_68), .in1(tmp00_93_68), .out(tmp01_46_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008683(.in0(tmp00_94_68), .in1(tmp00_95_68), .out(tmp01_47_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008684(.in0(tmp00_96_68), .in1(tmp00_97_68), .out(tmp01_48_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008685(.in0(tmp00_98_68), .in1(tmp00_99_68), .out(tmp01_49_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008686(.in0(tmp00_100_68), .in1(tmp00_101_68), .out(tmp01_50_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008687(.in0(tmp00_102_68), .in1(tmp00_103_68), .out(tmp01_51_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008688(.in0(tmp00_104_68), .in1(tmp00_105_68), .out(tmp01_52_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008689(.in0(tmp00_106_68), .in1(tmp00_107_68), .out(tmp01_53_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008690(.in0(tmp00_108_68), .in1(tmp00_109_68), .out(tmp01_54_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008691(.in0(tmp00_110_68), .in1(tmp00_111_68), .out(tmp01_55_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008692(.in0(tmp00_112_68), .in1(tmp00_113_68), .out(tmp01_56_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008693(.in0(tmp00_114_68), .in1(tmp00_115_68), .out(tmp01_57_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008694(.in0(tmp00_116_68), .in1(tmp00_117_68), .out(tmp01_58_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008695(.in0(tmp00_118_68), .in1(tmp00_119_68), .out(tmp01_59_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008696(.in0(tmp00_120_68), .in1(tmp00_121_68), .out(tmp01_60_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008697(.in0(tmp00_122_68), .in1(tmp00_123_68), .out(tmp01_61_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008698(.in0(tmp00_124_68), .in1(tmp00_125_68), .out(tmp01_62_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008699(.in0(tmp00_126_68), .in1(tmp00_127_68), .out(tmp01_63_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008700(.in0(tmp01_0_68), .in1(tmp01_1_68), .out(tmp02_0_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008701(.in0(tmp01_2_68), .in1(tmp01_3_68), .out(tmp02_1_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008702(.in0(tmp01_4_68), .in1(tmp01_5_68), .out(tmp02_2_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008703(.in0(tmp01_6_68), .in1(tmp01_7_68), .out(tmp02_3_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008704(.in0(tmp01_8_68), .in1(tmp01_9_68), .out(tmp02_4_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008705(.in0(tmp01_10_68), .in1(tmp01_11_68), .out(tmp02_5_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008706(.in0(tmp01_12_68), .in1(tmp01_13_68), .out(tmp02_6_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008707(.in0(tmp01_14_68), .in1(tmp01_15_68), .out(tmp02_7_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008708(.in0(tmp01_16_68), .in1(tmp01_17_68), .out(tmp02_8_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008709(.in0(tmp01_18_68), .in1(tmp01_19_68), .out(tmp02_9_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008710(.in0(tmp01_20_68), .in1(tmp01_21_68), .out(tmp02_10_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008711(.in0(tmp01_22_68), .in1(tmp01_23_68), .out(tmp02_11_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008712(.in0(tmp01_24_68), .in1(tmp01_25_68), .out(tmp02_12_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008713(.in0(tmp01_26_68), .in1(tmp01_27_68), .out(tmp02_13_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008714(.in0(tmp01_28_68), .in1(tmp01_29_68), .out(tmp02_14_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008715(.in0(tmp01_30_68), .in1(tmp01_31_68), .out(tmp02_15_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008716(.in0(tmp01_32_68), .in1(tmp01_33_68), .out(tmp02_16_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008717(.in0(tmp01_34_68), .in1(tmp01_35_68), .out(tmp02_17_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008718(.in0(tmp01_36_68), .in1(tmp01_37_68), .out(tmp02_18_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008719(.in0(tmp01_38_68), .in1(tmp01_39_68), .out(tmp02_19_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008720(.in0(tmp01_40_68), .in1(tmp01_41_68), .out(tmp02_20_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008721(.in0(tmp01_42_68), .in1(tmp01_43_68), .out(tmp02_21_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008722(.in0(tmp01_44_68), .in1(tmp01_45_68), .out(tmp02_22_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008723(.in0(tmp01_46_68), .in1(tmp01_47_68), .out(tmp02_23_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008724(.in0(tmp01_48_68), .in1(tmp01_49_68), .out(tmp02_24_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008725(.in0(tmp01_50_68), .in1(tmp01_51_68), .out(tmp02_25_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008726(.in0(tmp01_52_68), .in1(tmp01_53_68), .out(tmp02_26_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008727(.in0(tmp01_54_68), .in1(tmp01_55_68), .out(tmp02_27_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008728(.in0(tmp01_56_68), .in1(tmp01_57_68), .out(tmp02_28_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008729(.in0(tmp01_58_68), .in1(tmp01_59_68), .out(tmp02_29_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008730(.in0(tmp01_60_68), .in1(tmp01_61_68), .out(tmp02_30_68));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008731(.in0(tmp01_62_68), .in1(tmp01_63_68), .out(tmp02_31_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008732(.in0(tmp02_0_68), .in1(tmp02_1_68), .out(tmp03_0_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008733(.in0(tmp02_2_68), .in1(tmp02_3_68), .out(tmp03_1_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008734(.in0(tmp02_4_68), .in1(tmp02_5_68), .out(tmp03_2_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008735(.in0(tmp02_6_68), .in1(tmp02_7_68), .out(tmp03_3_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008736(.in0(tmp02_8_68), .in1(tmp02_9_68), .out(tmp03_4_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008737(.in0(tmp02_10_68), .in1(tmp02_11_68), .out(tmp03_5_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008738(.in0(tmp02_12_68), .in1(tmp02_13_68), .out(tmp03_6_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008739(.in0(tmp02_14_68), .in1(tmp02_15_68), .out(tmp03_7_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008740(.in0(tmp02_16_68), .in1(tmp02_17_68), .out(tmp03_8_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008741(.in0(tmp02_18_68), .in1(tmp02_19_68), .out(tmp03_9_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008742(.in0(tmp02_20_68), .in1(tmp02_21_68), .out(tmp03_10_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008743(.in0(tmp02_22_68), .in1(tmp02_23_68), .out(tmp03_11_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008744(.in0(tmp02_24_68), .in1(tmp02_25_68), .out(tmp03_12_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008745(.in0(tmp02_26_68), .in1(tmp02_27_68), .out(tmp03_13_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008746(.in0(tmp02_28_68), .in1(tmp02_29_68), .out(tmp03_14_68));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008747(.in0(tmp02_30_68), .in1(tmp02_31_68), .out(tmp03_15_68));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008748(.in0(tmp03_0_68), .in1(tmp03_1_68), .out(tmp04_0_68));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008749(.in0(tmp03_2_68), .in1(tmp03_3_68), .out(tmp04_1_68));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008750(.in0(tmp03_4_68), .in1(tmp03_5_68), .out(tmp04_2_68));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008751(.in0(tmp03_6_68), .in1(tmp03_7_68), .out(tmp04_3_68));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008752(.in0(tmp03_8_68), .in1(tmp03_9_68), .out(tmp04_4_68));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008753(.in0(tmp03_10_68), .in1(tmp03_11_68), .out(tmp04_5_68));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008754(.in0(tmp03_12_68), .in1(tmp03_13_68), .out(tmp04_6_68));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008755(.in0(tmp03_14_68), .in1(tmp03_15_68), .out(tmp04_7_68));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008756(.in0(tmp04_0_68), .in1(tmp04_1_68), .out(tmp05_0_68));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008757(.in0(tmp04_2_68), .in1(tmp04_3_68), .out(tmp05_1_68));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008758(.in0(tmp04_4_68), .in1(tmp04_5_68), .out(tmp05_2_68));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008759(.in0(tmp04_6_68), .in1(tmp04_7_68), .out(tmp05_3_68));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008760(.in0(tmp05_0_68), .in1(tmp05_1_68), .out(tmp06_0_68));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008761(.in0(tmp05_2_68), .in1(tmp05_3_68), .out(tmp06_1_68));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add008762(.in0(tmp06_0_68), .in1(tmp06_1_68), .out(tmp07_0_68));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008763(.in0(tmp00_0_69), .in1(tmp00_1_69), .out(tmp01_0_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008764(.in0(tmp00_2_69), .in1(tmp00_3_69), .out(tmp01_1_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008765(.in0(tmp00_4_69), .in1(tmp00_5_69), .out(tmp01_2_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008766(.in0(tmp00_6_69), .in1(tmp00_7_69), .out(tmp01_3_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008767(.in0(tmp00_8_69), .in1(tmp00_9_69), .out(tmp01_4_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008768(.in0(tmp00_10_69), .in1(tmp00_11_69), .out(tmp01_5_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008769(.in0(tmp00_12_69), .in1(tmp00_13_69), .out(tmp01_6_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008770(.in0(tmp00_14_69), .in1(tmp00_15_69), .out(tmp01_7_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008771(.in0(tmp00_16_69), .in1(tmp00_17_69), .out(tmp01_8_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008772(.in0(tmp00_18_69), .in1(tmp00_19_69), .out(tmp01_9_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008773(.in0(tmp00_20_69), .in1(tmp00_21_69), .out(tmp01_10_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008774(.in0(tmp00_22_69), .in1(tmp00_23_69), .out(tmp01_11_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008775(.in0(tmp00_24_69), .in1(tmp00_25_69), .out(tmp01_12_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008776(.in0(tmp00_26_69), .in1(tmp00_27_69), .out(tmp01_13_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008777(.in0(tmp00_28_69), .in1(tmp00_29_69), .out(tmp01_14_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008778(.in0(tmp00_30_69), .in1(tmp00_31_69), .out(tmp01_15_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008779(.in0(tmp00_32_69), .in1(tmp00_33_69), .out(tmp01_16_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008780(.in0(tmp00_34_69), .in1(tmp00_35_69), .out(tmp01_17_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008781(.in0(tmp00_36_69), .in1(tmp00_37_69), .out(tmp01_18_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008782(.in0(tmp00_38_69), .in1(tmp00_39_69), .out(tmp01_19_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008783(.in0(tmp00_40_69), .in1(tmp00_41_69), .out(tmp01_20_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008784(.in0(tmp00_42_69), .in1(tmp00_43_69), .out(tmp01_21_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008785(.in0(tmp00_44_69), .in1(tmp00_45_69), .out(tmp01_22_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008786(.in0(tmp00_46_69), .in1(tmp00_47_69), .out(tmp01_23_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008787(.in0(tmp00_48_69), .in1(tmp00_49_69), .out(tmp01_24_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008788(.in0(tmp00_50_69), .in1(tmp00_51_69), .out(tmp01_25_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008789(.in0(tmp00_52_69), .in1(tmp00_53_69), .out(tmp01_26_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008790(.in0(tmp00_54_69), .in1(tmp00_55_69), .out(tmp01_27_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008791(.in0(tmp00_56_69), .in1(tmp00_57_69), .out(tmp01_28_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008792(.in0(tmp00_58_69), .in1(tmp00_59_69), .out(tmp01_29_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008793(.in0(tmp00_60_69), .in1(tmp00_61_69), .out(tmp01_30_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008794(.in0(tmp00_62_69), .in1(tmp00_63_69), .out(tmp01_31_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008795(.in0(tmp00_64_69), .in1(tmp00_65_69), .out(tmp01_32_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008796(.in0(tmp00_66_69), .in1(tmp00_67_69), .out(tmp01_33_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008797(.in0(tmp00_68_69), .in1(tmp00_69_69), .out(tmp01_34_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008798(.in0(tmp00_70_69), .in1(tmp00_71_69), .out(tmp01_35_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008799(.in0(tmp00_72_69), .in1(tmp00_73_69), .out(tmp01_36_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008800(.in0(tmp00_74_69), .in1(tmp00_75_69), .out(tmp01_37_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008801(.in0(tmp00_76_69), .in1(tmp00_77_69), .out(tmp01_38_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008802(.in0(tmp00_78_69), .in1(tmp00_79_69), .out(tmp01_39_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008803(.in0(tmp00_80_69), .in1(tmp00_81_69), .out(tmp01_40_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008804(.in0(tmp00_82_69), .in1(tmp00_83_69), .out(tmp01_41_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008805(.in0(tmp00_84_69), .in1(tmp00_85_69), .out(tmp01_42_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008806(.in0(tmp00_86_69), .in1(tmp00_87_69), .out(tmp01_43_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008807(.in0(tmp00_88_69), .in1(tmp00_89_69), .out(tmp01_44_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008808(.in0(tmp00_90_69), .in1(tmp00_91_69), .out(tmp01_45_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008809(.in0(tmp00_92_69), .in1(tmp00_93_69), .out(tmp01_46_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008810(.in0(tmp00_94_69), .in1(tmp00_95_69), .out(tmp01_47_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008811(.in0(tmp00_96_69), .in1(tmp00_97_69), .out(tmp01_48_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008812(.in0(tmp00_98_69), .in1(tmp00_99_69), .out(tmp01_49_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008813(.in0(tmp00_100_69), .in1(tmp00_101_69), .out(tmp01_50_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008814(.in0(tmp00_102_69), .in1(tmp00_103_69), .out(tmp01_51_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008815(.in0(tmp00_104_69), .in1(tmp00_105_69), .out(tmp01_52_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008816(.in0(tmp00_106_69), .in1(tmp00_107_69), .out(tmp01_53_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008817(.in0(tmp00_108_69), .in1(tmp00_109_69), .out(tmp01_54_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008818(.in0(tmp00_110_69), .in1(tmp00_111_69), .out(tmp01_55_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008819(.in0(tmp00_112_69), .in1(tmp00_113_69), .out(tmp01_56_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008820(.in0(tmp00_114_69), .in1(tmp00_115_69), .out(tmp01_57_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008821(.in0(tmp00_116_69), .in1(tmp00_117_69), .out(tmp01_58_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008822(.in0(tmp00_118_69), .in1(tmp00_119_69), .out(tmp01_59_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008823(.in0(tmp00_120_69), .in1(tmp00_121_69), .out(tmp01_60_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008824(.in0(tmp00_122_69), .in1(tmp00_123_69), .out(tmp01_61_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008825(.in0(tmp00_124_69), .in1(tmp00_125_69), .out(tmp01_62_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008826(.in0(tmp00_126_69), .in1(tmp00_127_69), .out(tmp01_63_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008827(.in0(tmp01_0_69), .in1(tmp01_1_69), .out(tmp02_0_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008828(.in0(tmp01_2_69), .in1(tmp01_3_69), .out(tmp02_1_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008829(.in0(tmp01_4_69), .in1(tmp01_5_69), .out(tmp02_2_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008830(.in0(tmp01_6_69), .in1(tmp01_7_69), .out(tmp02_3_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008831(.in0(tmp01_8_69), .in1(tmp01_9_69), .out(tmp02_4_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008832(.in0(tmp01_10_69), .in1(tmp01_11_69), .out(tmp02_5_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008833(.in0(tmp01_12_69), .in1(tmp01_13_69), .out(tmp02_6_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008834(.in0(tmp01_14_69), .in1(tmp01_15_69), .out(tmp02_7_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008835(.in0(tmp01_16_69), .in1(tmp01_17_69), .out(tmp02_8_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008836(.in0(tmp01_18_69), .in1(tmp01_19_69), .out(tmp02_9_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008837(.in0(tmp01_20_69), .in1(tmp01_21_69), .out(tmp02_10_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008838(.in0(tmp01_22_69), .in1(tmp01_23_69), .out(tmp02_11_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008839(.in0(tmp01_24_69), .in1(tmp01_25_69), .out(tmp02_12_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008840(.in0(tmp01_26_69), .in1(tmp01_27_69), .out(tmp02_13_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008841(.in0(tmp01_28_69), .in1(tmp01_29_69), .out(tmp02_14_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008842(.in0(tmp01_30_69), .in1(tmp01_31_69), .out(tmp02_15_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008843(.in0(tmp01_32_69), .in1(tmp01_33_69), .out(tmp02_16_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008844(.in0(tmp01_34_69), .in1(tmp01_35_69), .out(tmp02_17_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008845(.in0(tmp01_36_69), .in1(tmp01_37_69), .out(tmp02_18_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008846(.in0(tmp01_38_69), .in1(tmp01_39_69), .out(tmp02_19_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008847(.in0(tmp01_40_69), .in1(tmp01_41_69), .out(tmp02_20_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008848(.in0(tmp01_42_69), .in1(tmp01_43_69), .out(tmp02_21_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008849(.in0(tmp01_44_69), .in1(tmp01_45_69), .out(tmp02_22_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008850(.in0(tmp01_46_69), .in1(tmp01_47_69), .out(tmp02_23_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008851(.in0(tmp01_48_69), .in1(tmp01_49_69), .out(tmp02_24_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008852(.in0(tmp01_50_69), .in1(tmp01_51_69), .out(tmp02_25_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008853(.in0(tmp01_52_69), .in1(tmp01_53_69), .out(tmp02_26_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008854(.in0(tmp01_54_69), .in1(tmp01_55_69), .out(tmp02_27_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008855(.in0(tmp01_56_69), .in1(tmp01_57_69), .out(tmp02_28_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008856(.in0(tmp01_58_69), .in1(tmp01_59_69), .out(tmp02_29_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008857(.in0(tmp01_60_69), .in1(tmp01_61_69), .out(tmp02_30_69));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008858(.in0(tmp01_62_69), .in1(tmp01_63_69), .out(tmp02_31_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008859(.in0(tmp02_0_69), .in1(tmp02_1_69), .out(tmp03_0_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008860(.in0(tmp02_2_69), .in1(tmp02_3_69), .out(tmp03_1_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008861(.in0(tmp02_4_69), .in1(tmp02_5_69), .out(tmp03_2_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008862(.in0(tmp02_6_69), .in1(tmp02_7_69), .out(tmp03_3_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008863(.in0(tmp02_8_69), .in1(tmp02_9_69), .out(tmp03_4_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008864(.in0(tmp02_10_69), .in1(tmp02_11_69), .out(tmp03_5_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008865(.in0(tmp02_12_69), .in1(tmp02_13_69), .out(tmp03_6_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008866(.in0(tmp02_14_69), .in1(tmp02_15_69), .out(tmp03_7_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008867(.in0(tmp02_16_69), .in1(tmp02_17_69), .out(tmp03_8_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008868(.in0(tmp02_18_69), .in1(tmp02_19_69), .out(tmp03_9_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008869(.in0(tmp02_20_69), .in1(tmp02_21_69), .out(tmp03_10_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008870(.in0(tmp02_22_69), .in1(tmp02_23_69), .out(tmp03_11_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008871(.in0(tmp02_24_69), .in1(tmp02_25_69), .out(tmp03_12_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008872(.in0(tmp02_26_69), .in1(tmp02_27_69), .out(tmp03_13_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008873(.in0(tmp02_28_69), .in1(tmp02_29_69), .out(tmp03_14_69));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008874(.in0(tmp02_30_69), .in1(tmp02_31_69), .out(tmp03_15_69));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008875(.in0(tmp03_0_69), .in1(tmp03_1_69), .out(tmp04_0_69));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008876(.in0(tmp03_2_69), .in1(tmp03_3_69), .out(tmp04_1_69));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008877(.in0(tmp03_4_69), .in1(tmp03_5_69), .out(tmp04_2_69));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008878(.in0(tmp03_6_69), .in1(tmp03_7_69), .out(tmp04_3_69));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008879(.in0(tmp03_8_69), .in1(tmp03_9_69), .out(tmp04_4_69));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008880(.in0(tmp03_10_69), .in1(tmp03_11_69), .out(tmp04_5_69));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008881(.in0(tmp03_12_69), .in1(tmp03_13_69), .out(tmp04_6_69));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add008882(.in0(tmp03_14_69), .in1(tmp03_15_69), .out(tmp04_7_69));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008883(.in0(tmp04_0_69), .in1(tmp04_1_69), .out(tmp05_0_69));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008884(.in0(tmp04_2_69), .in1(tmp04_3_69), .out(tmp05_1_69));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008885(.in0(tmp04_4_69), .in1(tmp04_5_69), .out(tmp05_2_69));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add008886(.in0(tmp04_6_69), .in1(tmp04_7_69), .out(tmp05_3_69));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008887(.in0(tmp05_0_69), .in1(tmp05_1_69), .out(tmp06_0_69));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add008888(.in0(tmp05_2_69), .in1(tmp05_3_69), .out(tmp06_1_69));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add008889(.in0(tmp06_0_69), .in1(tmp06_1_69), .out(tmp07_0_69));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008890(.in0(tmp00_0_70), .in1(tmp00_1_70), .out(tmp01_0_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008891(.in0(tmp00_2_70), .in1(tmp00_3_70), .out(tmp01_1_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008892(.in0(tmp00_4_70), .in1(tmp00_5_70), .out(tmp01_2_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008893(.in0(tmp00_6_70), .in1(tmp00_7_70), .out(tmp01_3_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008894(.in0(tmp00_8_70), .in1(tmp00_9_70), .out(tmp01_4_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008895(.in0(tmp00_10_70), .in1(tmp00_11_70), .out(tmp01_5_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008896(.in0(tmp00_12_70), .in1(tmp00_13_70), .out(tmp01_6_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008897(.in0(tmp00_14_70), .in1(tmp00_15_70), .out(tmp01_7_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008898(.in0(tmp00_16_70), .in1(tmp00_17_70), .out(tmp01_8_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008899(.in0(tmp00_18_70), .in1(tmp00_19_70), .out(tmp01_9_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008900(.in0(tmp00_20_70), .in1(tmp00_21_70), .out(tmp01_10_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008901(.in0(tmp00_22_70), .in1(tmp00_23_70), .out(tmp01_11_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008902(.in0(tmp00_24_70), .in1(tmp00_25_70), .out(tmp01_12_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008903(.in0(tmp00_26_70), .in1(tmp00_27_70), .out(tmp01_13_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008904(.in0(tmp00_28_70), .in1(tmp00_29_70), .out(tmp01_14_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008905(.in0(tmp00_30_70), .in1(tmp00_31_70), .out(tmp01_15_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008906(.in0(tmp00_32_70), .in1(tmp00_33_70), .out(tmp01_16_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008907(.in0(tmp00_34_70), .in1(tmp00_35_70), .out(tmp01_17_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008908(.in0(tmp00_36_70), .in1(tmp00_37_70), .out(tmp01_18_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008909(.in0(tmp00_38_70), .in1(tmp00_39_70), .out(tmp01_19_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008910(.in0(tmp00_40_70), .in1(tmp00_41_70), .out(tmp01_20_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008911(.in0(tmp00_42_70), .in1(tmp00_43_70), .out(tmp01_21_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008912(.in0(tmp00_44_70), .in1(tmp00_45_70), .out(tmp01_22_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008913(.in0(tmp00_46_70), .in1(tmp00_47_70), .out(tmp01_23_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008914(.in0(tmp00_48_70), .in1(tmp00_49_70), .out(tmp01_24_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008915(.in0(tmp00_50_70), .in1(tmp00_51_70), .out(tmp01_25_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008916(.in0(tmp00_52_70), .in1(tmp00_53_70), .out(tmp01_26_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008917(.in0(tmp00_54_70), .in1(tmp00_55_70), .out(tmp01_27_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008918(.in0(tmp00_56_70), .in1(tmp00_57_70), .out(tmp01_28_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008919(.in0(tmp00_58_70), .in1(tmp00_59_70), .out(tmp01_29_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008920(.in0(tmp00_60_70), .in1(tmp00_61_70), .out(tmp01_30_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008921(.in0(tmp00_62_70), .in1(tmp00_63_70), .out(tmp01_31_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008922(.in0(tmp00_64_70), .in1(tmp00_65_70), .out(tmp01_32_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008923(.in0(tmp00_66_70), .in1(tmp00_67_70), .out(tmp01_33_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008924(.in0(tmp00_68_70), .in1(tmp00_69_70), .out(tmp01_34_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008925(.in0(tmp00_70_70), .in1(tmp00_71_70), .out(tmp01_35_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008926(.in0(tmp00_72_70), .in1(tmp00_73_70), .out(tmp01_36_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008927(.in0(tmp00_74_70), .in1(tmp00_75_70), .out(tmp01_37_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008928(.in0(tmp00_76_70), .in1(tmp00_77_70), .out(tmp01_38_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008929(.in0(tmp00_78_70), .in1(tmp00_79_70), .out(tmp01_39_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008930(.in0(tmp00_80_70), .in1(tmp00_81_70), .out(tmp01_40_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008931(.in0(tmp00_82_70), .in1(tmp00_83_70), .out(tmp01_41_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008932(.in0(tmp00_84_70), .in1(tmp00_85_70), .out(tmp01_42_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008933(.in0(tmp00_86_70), .in1(tmp00_87_70), .out(tmp01_43_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008934(.in0(tmp00_88_70), .in1(tmp00_89_70), .out(tmp01_44_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008935(.in0(tmp00_90_70), .in1(tmp00_91_70), .out(tmp01_45_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008936(.in0(tmp00_92_70), .in1(tmp00_93_70), .out(tmp01_46_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008937(.in0(tmp00_94_70), .in1(tmp00_95_70), .out(tmp01_47_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008938(.in0(tmp00_96_70), .in1(tmp00_97_70), .out(tmp01_48_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008939(.in0(tmp00_98_70), .in1(tmp00_99_70), .out(tmp01_49_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008940(.in0(tmp00_100_70), .in1(tmp00_101_70), .out(tmp01_50_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008941(.in0(tmp00_102_70), .in1(tmp00_103_70), .out(tmp01_51_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008942(.in0(tmp00_104_70), .in1(tmp00_105_70), .out(tmp01_52_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008943(.in0(tmp00_106_70), .in1(tmp00_107_70), .out(tmp01_53_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008944(.in0(tmp00_108_70), .in1(tmp00_109_70), .out(tmp01_54_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008945(.in0(tmp00_110_70), .in1(tmp00_111_70), .out(tmp01_55_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008946(.in0(tmp00_112_70), .in1(tmp00_113_70), .out(tmp01_56_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008947(.in0(tmp00_114_70), .in1(tmp00_115_70), .out(tmp01_57_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008948(.in0(tmp00_116_70), .in1(tmp00_117_70), .out(tmp01_58_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008949(.in0(tmp00_118_70), .in1(tmp00_119_70), .out(tmp01_59_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008950(.in0(tmp00_120_70), .in1(tmp00_121_70), .out(tmp01_60_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008951(.in0(tmp00_122_70), .in1(tmp00_123_70), .out(tmp01_61_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008952(.in0(tmp00_124_70), .in1(tmp00_125_70), .out(tmp01_62_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add008953(.in0(tmp00_126_70), .in1(tmp00_127_70), .out(tmp01_63_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008954(.in0(tmp01_0_70), .in1(tmp01_1_70), .out(tmp02_0_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008955(.in0(tmp01_2_70), .in1(tmp01_3_70), .out(tmp02_1_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008956(.in0(tmp01_4_70), .in1(tmp01_5_70), .out(tmp02_2_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008957(.in0(tmp01_6_70), .in1(tmp01_7_70), .out(tmp02_3_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008958(.in0(tmp01_8_70), .in1(tmp01_9_70), .out(tmp02_4_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008959(.in0(tmp01_10_70), .in1(tmp01_11_70), .out(tmp02_5_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008960(.in0(tmp01_12_70), .in1(tmp01_13_70), .out(tmp02_6_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008961(.in0(tmp01_14_70), .in1(tmp01_15_70), .out(tmp02_7_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008962(.in0(tmp01_16_70), .in1(tmp01_17_70), .out(tmp02_8_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008963(.in0(tmp01_18_70), .in1(tmp01_19_70), .out(tmp02_9_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008964(.in0(tmp01_20_70), .in1(tmp01_21_70), .out(tmp02_10_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008965(.in0(tmp01_22_70), .in1(tmp01_23_70), .out(tmp02_11_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008966(.in0(tmp01_24_70), .in1(tmp01_25_70), .out(tmp02_12_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008967(.in0(tmp01_26_70), .in1(tmp01_27_70), .out(tmp02_13_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008968(.in0(tmp01_28_70), .in1(tmp01_29_70), .out(tmp02_14_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008969(.in0(tmp01_30_70), .in1(tmp01_31_70), .out(tmp02_15_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008970(.in0(tmp01_32_70), .in1(tmp01_33_70), .out(tmp02_16_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008971(.in0(tmp01_34_70), .in1(tmp01_35_70), .out(tmp02_17_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008972(.in0(tmp01_36_70), .in1(tmp01_37_70), .out(tmp02_18_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008973(.in0(tmp01_38_70), .in1(tmp01_39_70), .out(tmp02_19_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008974(.in0(tmp01_40_70), .in1(tmp01_41_70), .out(tmp02_20_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008975(.in0(tmp01_42_70), .in1(tmp01_43_70), .out(tmp02_21_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008976(.in0(tmp01_44_70), .in1(tmp01_45_70), .out(tmp02_22_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008977(.in0(tmp01_46_70), .in1(tmp01_47_70), .out(tmp02_23_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008978(.in0(tmp01_48_70), .in1(tmp01_49_70), .out(tmp02_24_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008979(.in0(tmp01_50_70), .in1(tmp01_51_70), .out(tmp02_25_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008980(.in0(tmp01_52_70), .in1(tmp01_53_70), .out(tmp02_26_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008981(.in0(tmp01_54_70), .in1(tmp01_55_70), .out(tmp02_27_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008982(.in0(tmp01_56_70), .in1(tmp01_57_70), .out(tmp02_28_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008983(.in0(tmp01_58_70), .in1(tmp01_59_70), .out(tmp02_29_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008984(.in0(tmp01_60_70), .in1(tmp01_61_70), .out(tmp02_30_70));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add008985(.in0(tmp01_62_70), .in1(tmp01_63_70), .out(tmp02_31_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008986(.in0(tmp02_0_70), .in1(tmp02_1_70), .out(tmp03_0_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008987(.in0(tmp02_2_70), .in1(tmp02_3_70), .out(tmp03_1_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008988(.in0(tmp02_4_70), .in1(tmp02_5_70), .out(tmp03_2_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008989(.in0(tmp02_6_70), .in1(tmp02_7_70), .out(tmp03_3_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008990(.in0(tmp02_8_70), .in1(tmp02_9_70), .out(tmp03_4_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008991(.in0(tmp02_10_70), .in1(tmp02_11_70), .out(tmp03_5_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008992(.in0(tmp02_12_70), .in1(tmp02_13_70), .out(tmp03_6_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008993(.in0(tmp02_14_70), .in1(tmp02_15_70), .out(tmp03_7_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008994(.in0(tmp02_16_70), .in1(tmp02_17_70), .out(tmp03_8_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008995(.in0(tmp02_18_70), .in1(tmp02_19_70), .out(tmp03_9_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008996(.in0(tmp02_20_70), .in1(tmp02_21_70), .out(tmp03_10_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008997(.in0(tmp02_22_70), .in1(tmp02_23_70), .out(tmp03_11_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008998(.in0(tmp02_24_70), .in1(tmp02_25_70), .out(tmp03_12_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add008999(.in0(tmp02_26_70), .in1(tmp02_27_70), .out(tmp03_13_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009000(.in0(tmp02_28_70), .in1(tmp02_29_70), .out(tmp03_14_70));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009001(.in0(tmp02_30_70), .in1(tmp02_31_70), .out(tmp03_15_70));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009002(.in0(tmp03_0_70), .in1(tmp03_1_70), .out(tmp04_0_70));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009003(.in0(tmp03_2_70), .in1(tmp03_3_70), .out(tmp04_1_70));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009004(.in0(tmp03_4_70), .in1(tmp03_5_70), .out(tmp04_2_70));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009005(.in0(tmp03_6_70), .in1(tmp03_7_70), .out(tmp04_3_70));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009006(.in0(tmp03_8_70), .in1(tmp03_9_70), .out(tmp04_4_70));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009007(.in0(tmp03_10_70), .in1(tmp03_11_70), .out(tmp04_5_70));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009008(.in0(tmp03_12_70), .in1(tmp03_13_70), .out(tmp04_6_70));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009009(.in0(tmp03_14_70), .in1(tmp03_15_70), .out(tmp04_7_70));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009010(.in0(tmp04_0_70), .in1(tmp04_1_70), .out(tmp05_0_70));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009011(.in0(tmp04_2_70), .in1(tmp04_3_70), .out(tmp05_1_70));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009012(.in0(tmp04_4_70), .in1(tmp04_5_70), .out(tmp05_2_70));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009013(.in0(tmp04_6_70), .in1(tmp04_7_70), .out(tmp05_3_70));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009014(.in0(tmp05_0_70), .in1(tmp05_1_70), .out(tmp06_0_70));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009015(.in0(tmp05_2_70), .in1(tmp05_3_70), .out(tmp06_1_70));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add009016(.in0(tmp06_0_70), .in1(tmp06_1_70), .out(tmp07_0_70));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009017(.in0(tmp00_0_71), .in1(tmp00_1_71), .out(tmp01_0_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009018(.in0(tmp00_2_71), .in1(tmp00_3_71), .out(tmp01_1_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009019(.in0(tmp00_4_71), .in1(tmp00_5_71), .out(tmp01_2_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009020(.in0(tmp00_6_71), .in1(tmp00_7_71), .out(tmp01_3_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009021(.in0(tmp00_8_71), .in1(tmp00_9_71), .out(tmp01_4_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009022(.in0(tmp00_10_71), .in1(tmp00_11_71), .out(tmp01_5_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009023(.in0(tmp00_12_71), .in1(tmp00_13_71), .out(tmp01_6_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009024(.in0(tmp00_14_71), .in1(tmp00_15_71), .out(tmp01_7_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009025(.in0(tmp00_16_71), .in1(tmp00_17_71), .out(tmp01_8_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009026(.in0(tmp00_18_71), .in1(tmp00_19_71), .out(tmp01_9_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009027(.in0(tmp00_20_71), .in1(tmp00_21_71), .out(tmp01_10_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009028(.in0(tmp00_22_71), .in1(tmp00_23_71), .out(tmp01_11_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009029(.in0(tmp00_24_71), .in1(tmp00_25_71), .out(tmp01_12_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009030(.in0(tmp00_26_71), .in1(tmp00_27_71), .out(tmp01_13_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009031(.in0(tmp00_28_71), .in1(tmp00_29_71), .out(tmp01_14_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009032(.in0(tmp00_30_71), .in1(tmp00_31_71), .out(tmp01_15_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009033(.in0(tmp00_32_71), .in1(tmp00_33_71), .out(tmp01_16_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009034(.in0(tmp00_34_71), .in1(tmp00_35_71), .out(tmp01_17_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009035(.in0(tmp00_36_71), .in1(tmp00_37_71), .out(tmp01_18_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009036(.in0(tmp00_38_71), .in1(tmp00_39_71), .out(tmp01_19_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009037(.in0(tmp00_40_71), .in1(tmp00_41_71), .out(tmp01_20_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009038(.in0(tmp00_42_71), .in1(tmp00_43_71), .out(tmp01_21_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009039(.in0(tmp00_44_71), .in1(tmp00_45_71), .out(tmp01_22_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009040(.in0(tmp00_46_71), .in1(tmp00_47_71), .out(tmp01_23_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009041(.in0(tmp00_48_71), .in1(tmp00_49_71), .out(tmp01_24_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009042(.in0(tmp00_50_71), .in1(tmp00_51_71), .out(tmp01_25_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009043(.in0(tmp00_52_71), .in1(tmp00_53_71), .out(tmp01_26_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009044(.in0(tmp00_54_71), .in1(tmp00_55_71), .out(tmp01_27_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009045(.in0(tmp00_56_71), .in1(tmp00_57_71), .out(tmp01_28_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009046(.in0(tmp00_58_71), .in1(tmp00_59_71), .out(tmp01_29_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009047(.in0(tmp00_60_71), .in1(tmp00_61_71), .out(tmp01_30_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009048(.in0(tmp00_62_71), .in1(tmp00_63_71), .out(tmp01_31_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009049(.in0(tmp00_64_71), .in1(tmp00_65_71), .out(tmp01_32_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009050(.in0(tmp00_66_71), .in1(tmp00_67_71), .out(tmp01_33_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009051(.in0(tmp00_68_71), .in1(tmp00_69_71), .out(tmp01_34_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009052(.in0(tmp00_70_71), .in1(tmp00_71_71), .out(tmp01_35_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009053(.in0(tmp00_72_71), .in1(tmp00_73_71), .out(tmp01_36_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009054(.in0(tmp00_74_71), .in1(tmp00_75_71), .out(tmp01_37_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009055(.in0(tmp00_76_71), .in1(tmp00_77_71), .out(tmp01_38_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009056(.in0(tmp00_78_71), .in1(tmp00_79_71), .out(tmp01_39_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009057(.in0(tmp00_80_71), .in1(tmp00_81_71), .out(tmp01_40_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009058(.in0(tmp00_82_71), .in1(tmp00_83_71), .out(tmp01_41_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009059(.in0(tmp00_84_71), .in1(tmp00_85_71), .out(tmp01_42_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009060(.in0(tmp00_86_71), .in1(tmp00_87_71), .out(tmp01_43_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009061(.in0(tmp00_88_71), .in1(tmp00_89_71), .out(tmp01_44_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009062(.in0(tmp00_90_71), .in1(tmp00_91_71), .out(tmp01_45_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009063(.in0(tmp00_92_71), .in1(tmp00_93_71), .out(tmp01_46_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009064(.in0(tmp00_94_71), .in1(tmp00_95_71), .out(tmp01_47_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009065(.in0(tmp00_96_71), .in1(tmp00_97_71), .out(tmp01_48_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009066(.in0(tmp00_98_71), .in1(tmp00_99_71), .out(tmp01_49_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009067(.in0(tmp00_100_71), .in1(tmp00_101_71), .out(tmp01_50_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009068(.in0(tmp00_102_71), .in1(tmp00_103_71), .out(tmp01_51_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009069(.in0(tmp00_104_71), .in1(tmp00_105_71), .out(tmp01_52_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009070(.in0(tmp00_106_71), .in1(tmp00_107_71), .out(tmp01_53_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009071(.in0(tmp00_108_71), .in1(tmp00_109_71), .out(tmp01_54_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009072(.in0(tmp00_110_71), .in1(tmp00_111_71), .out(tmp01_55_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009073(.in0(tmp00_112_71), .in1(tmp00_113_71), .out(tmp01_56_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009074(.in0(tmp00_114_71), .in1(tmp00_115_71), .out(tmp01_57_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009075(.in0(tmp00_116_71), .in1(tmp00_117_71), .out(tmp01_58_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009076(.in0(tmp00_118_71), .in1(tmp00_119_71), .out(tmp01_59_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009077(.in0(tmp00_120_71), .in1(tmp00_121_71), .out(tmp01_60_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009078(.in0(tmp00_122_71), .in1(tmp00_123_71), .out(tmp01_61_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009079(.in0(tmp00_124_71), .in1(tmp00_125_71), .out(tmp01_62_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009080(.in0(tmp00_126_71), .in1(tmp00_127_71), .out(tmp01_63_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009081(.in0(tmp01_0_71), .in1(tmp01_1_71), .out(tmp02_0_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009082(.in0(tmp01_2_71), .in1(tmp01_3_71), .out(tmp02_1_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009083(.in0(tmp01_4_71), .in1(tmp01_5_71), .out(tmp02_2_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009084(.in0(tmp01_6_71), .in1(tmp01_7_71), .out(tmp02_3_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009085(.in0(tmp01_8_71), .in1(tmp01_9_71), .out(tmp02_4_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009086(.in0(tmp01_10_71), .in1(tmp01_11_71), .out(tmp02_5_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009087(.in0(tmp01_12_71), .in1(tmp01_13_71), .out(tmp02_6_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009088(.in0(tmp01_14_71), .in1(tmp01_15_71), .out(tmp02_7_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009089(.in0(tmp01_16_71), .in1(tmp01_17_71), .out(tmp02_8_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009090(.in0(tmp01_18_71), .in1(tmp01_19_71), .out(tmp02_9_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009091(.in0(tmp01_20_71), .in1(tmp01_21_71), .out(tmp02_10_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009092(.in0(tmp01_22_71), .in1(tmp01_23_71), .out(tmp02_11_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009093(.in0(tmp01_24_71), .in1(tmp01_25_71), .out(tmp02_12_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009094(.in0(tmp01_26_71), .in1(tmp01_27_71), .out(tmp02_13_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009095(.in0(tmp01_28_71), .in1(tmp01_29_71), .out(tmp02_14_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009096(.in0(tmp01_30_71), .in1(tmp01_31_71), .out(tmp02_15_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009097(.in0(tmp01_32_71), .in1(tmp01_33_71), .out(tmp02_16_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009098(.in0(tmp01_34_71), .in1(tmp01_35_71), .out(tmp02_17_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009099(.in0(tmp01_36_71), .in1(tmp01_37_71), .out(tmp02_18_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009100(.in0(tmp01_38_71), .in1(tmp01_39_71), .out(tmp02_19_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009101(.in0(tmp01_40_71), .in1(tmp01_41_71), .out(tmp02_20_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009102(.in0(tmp01_42_71), .in1(tmp01_43_71), .out(tmp02_21_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009103(.in0(tmp01_44_71), .in1(tmp01_45_71), .out(tmp02_22_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009104(.in0(tmp01_46_71), .in1(tmp01_47_71), .out(tmp02_23_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009105(.in0(tmp01_48_71), .in1(tmp01_49_71), .out(tmp02_24_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009106(.in0(tmp01_50_71), .in1(tmp01_51_71), .out(tmp02_25_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009107(.in0(tmp01_52_71), .in1(tmp01_53_71), .out(tmp02_26_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009108(.in0(tmp01_54_71), .in1(tmp01_55_71), .out(tmp02_27_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009109(.in0(tmp01_56_71), .in1(tmp01_57_71), .out(tmp02_28_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009110(.in0(tmp01_58_71), .in1(tmp01_59_71), .out(tmp02_29_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009111(.in0(tmp01_60_71), .in1(tmp01_61_71), .out(tmp02_30_71));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009112(.in0(tmp01_62_71), .in1(tmp01_63_71), .out(tmp02_31_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009113(.in0(tmp02_0_71), .in1(tmp02_1_71), .out(tmp03_0_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009114(.in0(tmp02_2_71), .in1(tmp02_3_71), .out(tmp03_1_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009115(.in0(tmp02_4_71), .in1(tmp02_5_71), .out(tmp03_2_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009116(.in0(tmp02_6_71), .in1(tmp02_7_71), .out(tmp03_3_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009117(.in0(tmp02_8_71), .in1(tmp02_9_71), .out(tmp03_4_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009118(.in0(tmp02_10_71), .in1(tmp02_11_71), .out(tmp03_5_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009119(.in0(tmp02_12_71), .in1(tmp02_13_71), .out(tmp03_6_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009120(.in0(tmp02_14_71), .in1(tmp02_15_71), .out(tmp03_7_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009121(.in0(tmp02_16_71), .in1(tmp02_17_71), .out(tmp03_8_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009122(.in0(tmp02_18_71), .in1(tmp02_19_71), .out(tmp03_9_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009123(.in0(tmp02_20_71), .in1(tmp02_21_71), .out(tmp03_10_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009124(.in0(tmp02_22_71), .in1(tmp02_23_71), .out(tmp03_11_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009125(.in0(tmp02_24_71), .in1(tmp02_25_71), .out(tmp03_12_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009126(.in0(tmp02_26_71), .in1(tmp02_27_71), .out(tmp03_13_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009127(.in0(tmp02_28_71), .in1(tmp02_29_71), .out(tmp03_14_71));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009128(.in0(tmp02_30_71), .in1(tmp02_31_71), .out(tmp03_15_71));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009129(.in0(tmp03_0_71), .in1(tmp03_1_71), .out(tmp04_0_71));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009130(.in0(tmp03_2_71), .in1(tmp03_3_71), .out(tmp04_1_71));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009131(.in0(tmp03_4_71), .in1(tmp03_5_71), .out(tmp04_2_71));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009132(.in0(tmp03_6_71), .in1(tmp03_7_71), .out(tmp04_3_71));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009133(.in0(tmp03_8_71), .in1(tmp03_9_71), .out(tmp04_4_71));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009134(.in0(tmp03_10_71), .in1(tmp03_11_71), .out(tmp04_5_71));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009135(.in0(tmp03_12_71), .in1(tmp03_13_71), .out(tmp04_6_71));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009136(.in0(tmp03_14_71), .in1(tmp03_15_71), .out(tmp04_7_71));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009137(.in0(tmp04_0_71), .in1(tmp04_1_71), .out(tmp05_0_71));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009138(.in0(tmp04_2_71), .in1(tmp04_3_71), .out(tmp05_1_71));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009139(.in0(tmp04_4_71), .in1(tmp04_5_71), .out(tmp05_2_71));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009140(.in0(tmp04_6_71), .in1(tmp04_7_71), .out(tmp05_3_71));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009141(.in0(tmp05_0_71), .in1(tmp05_1_71), .out(tmp06_0_71));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009142(.in0(tmp05_2_71), .in1(tmp05_3_71), .out(tmp06_1_71));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add009143(.in0(tmp06_0_71), .in1(tmp06_1_71), .out(tmp07_0_71));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009144(.in0(tmp00_0_72), .in1(tmp00_1_72), .out(tmp01_0_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009145(.in0(tmp00_2_72), .in1(tmp00_3_72), .out(tmp01_1_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009146(.in0(tmp00_4_72), .in1(tmp00_5_72), .out(tmp01_2_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009147(.in0(tmp00_6_72), .in1(tmp00_7_72), .out(tmp01_3_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009148(.in0(tmp00_8_72), .in1(tmp00_9_72), .out(tmp01_4_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009149(.in0(tmp00_10_72), .in1(tmp00_11_72), .out(tmp01_5_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009150(.in0(tmp00_12_72), .in1(tmp00_13_72), .out(tmp01_6_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009151(.in0(tmp00_14_72), .in1(tmp00_15_72), .out(tmp01_7_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009152(.in0(tmp00_16_72), .in1(tmp00_17_72), .out(tmp01_8_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009153(.in0(tmp00_18_72), .in1(tmp00_19_72), .out(tmp01_9_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009154(.in0(tmp00_20_72), .in1(tmp00_21_72), .out(tmp01_10_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009155(.in0(tmp00_22_72), .in1(tmp00_23_72), .out(tmp01_11_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009156(.in0(tmp00_24_72), .in1(tmp00_25_72), .out(tmp01_12_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009157(.in0(tmp00_26_72), .in1(tmp00_27_72), .out(tmp01_13_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009158(.in0(tmp00_28_72), .in1(tmp00_29_72), .out(tmp01_14_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009159(.in0(tmp00_30_72), .in1(tmp00_31_72), .out(tmp01_15_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009160(.in0(tmp00_32_72), .in1(tmp00_33_72), .out(tmp01_16_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009161(.in0(tmp00_34_72), .in1(tmp00_35_72), .out(tmp01_17_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009162(.in0(tmp00_36_72), .in1(tmp00_37_72), .out(tmp01_18_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009163(.in0(tmp00_38_72), .in1(tmp00_39_72), .out(tmp01_19_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009164(.in0(tmp00_40_72), .in1(tmp00_41_72), .out(tmp01_20_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009165(.in0(tmp00_42_72), .in1(tmp00_43_72), .out(tmp01_21_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009166(.in0(tmp00_44_72), .in1(tmp00_45_72), .out(tmp01_22_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009167(.in0(tmp00_46_72), .in1(tmp00_47_72), .out(tmp01_23_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009168(.in0(tmp00_48_72), .in1(tmp00_49_72), .out(tmp01_24_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009169(.in0(tmp00_50_72), .in1(tmp00_51_72), .out(tmp01_25_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009170(.in0(tmp00_52_72), .in1(tmp00_53_72), .out(tmp01_26_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009171(.in0(tmp00_54_72), .in1(tmp00_55_72), .out(tmp01_27_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009172(.in0(tmp00_56_72), .in1(tmp00_57_72), .out(tmp01_28_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009173(.in0(tmp00_58_72), .in1(tmp00_59_72), .out(tmp01_29_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009174(.in0(tmp00_60_72), .in1(tmp00_61_72), .out(tmp01_30_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009175(.in0(tmp00_62_72), .in1(tmp00_63_72), .out(tmp01_31_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009176(.in0(tmp00_64_72), .in1(tmp00_65_72), .out(tmp01_32_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009177(.in0(tmp00_66_72), .in1(tmp00_67_72), .out(tmp01_33_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009178(.in0(tmp00_68_72), .in1(tmp00_69_72), .out(tmp01_34_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009179(.in0(tmp00_70_72), .in1(tmp00_71_72), .out(tmp01_35_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009180(.in0(tmp00_72_72), .in1(tmp00_73_72), .out(tmp01_36_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009181(.in0(tmp00_74_72), .in1(tmp00_75_72), .out(tmp01_37_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009182(.in0(tmp00_76_72), .in1(tmp00_77_72), .out(tmp01_38_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009183(.in0(tmp00_78_72), .in1(tmp00_79_72), .out(tmp01_39_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009184(.in0(tmp00_80_72), .in1(tmp00_81_72), .out(tmp01_40_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009185(.in0(tmp00_82_72), .in1(tmp00_83_72), .out(tmp01_41_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009186(.in0(tmp00_84_72), .in1(tmp00_85_72), .out(tmp01_42_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009187(.in0(tmp00_86_72), .in1(tmp00_87_72), .out(tmp01_43_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009188(.in0(tmp00_88_72), .in1(tmp00_89_72), .out(tmp01_44_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009189(.in0(tmp00_90_72), .in1(tmp00_91_72), .out(tmp01_45_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009190(.in0(tmp00_92_72), .in1(tmp00_93_72), .out(tmp01_46_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009191(.in0(tmp00_94_72), .in1(tmp00_95_72), .out(tmp01_47_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009192(.in0(tmp00_96_72), .in1(tmp00_97_72), .out(tmp01_48_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009193(.in0(tmp00_98_72), .in1(tmp00_99_72), .out(tmp01_49_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009194(.in0(tmp00_100_72), .in1(tmp00_101_72), .out(tmp01_50_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009195(.in0(tmp00_102_72), .in1(tmp00_103_72), .out(tmp01_51_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009196(.in0(tmp00_104_72), .in1(tmp00_105_72), .out(tmp01_52_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009197(.in0(tmp00_106_72), .in1(tmp00_107_72), .out(tmp01_53_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009198(.in0(tmp00_108_72), .in1(tmp00_109_72), .out(tmp01_54_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009199(.in0(tmp00_110_72), .in1(tmp00_111_72), .out(tmp01_55_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009200(.in0(tmp00_112_72), .in1(tmp00_113_72), .out(tmp01_56_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009201(.in0(tmp00_114_72), .in1(tmp00_115_72), .out(tmp01_57_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009202(.in0(tmp00_116_72), .in1(tmp00_117_72), .out(tmp01_58_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009203(.in0(tmp00_118_72), .in1(tmp00_119_72), .out(tmp01_59_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009204(.in0(tmp00_120_72), .in1(tmp00_121_72), .out(tmp01_60_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009205(.in0(tmp00_122_72), .in1(tmp00_123_72), .out(tmp01_61_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009206(.in0(tmp00_124_72), .in1(tmp00_125_72), .out(tmp01_62_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009207(.in0(tmp00_126_72), .in1(tmp00_127_72), .out(tmp01_63_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009208(.in0(tmp01_0_72), .in1(tmp01_1_72), .out(tmp02_0_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009209(.in0(tmp01_2_72), .in1(tmp01_3_72), .out(tmp02_1_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009210(.in0(tmp01_4_72), .in1(tmp01_5_72), .out(tmp02_2_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009211(.in0(tmp01_6_72), .in1(tmp01_7_72), .out(tmp02_3_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009212(.in0(tmp01_8_72), .in1(tmp01_9_72), .out(tmp02_4_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009213(.in0(tmp01_10_72), .in1(tmp01_11_72), .out(tmp02_5_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009214(.in0(tmp01_12_72), .in1(tmp01_13_72), .out(tmp02_6_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009215(.in0(tmp01_14_72), .in1(tmp01_15_72), .out(tmp02_7_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009216(.in0(tmp01_16_72), .in1(tmp01_17_72), .out(tmp02_8_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009217(.in0(tmp01_18_72), .in1(tmp01_19_72), .out(tmp02_9_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009218(.in0(tmp01_20_72), .in1(tmp01_21_72), .out(tmp02_10_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009219(.in0(tmp01_22_72), .in1(tmp01_23_72), .out(tmp02_11_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009220(.in0(tmp01_24_72), .in1(tmp01_25_72), .out(tmp02_12_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009221(.in0(tmp01_26_72), .in1(tmp01_27_72), .out(tmp02_13_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009222(.in0(tmp01_28_72), .in1(tmp01_29_72), .out(tmp02_14_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009223(.in0(tmp01_30_72), .in1(tmp01_31_72), .out(tmp02_15_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009224(.in0(tmp01_32_72), .in1(tmp01_33_72), .out(tmp02_16_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009225(.in0(tmp01_34_72), .in1(tmp01_35_72), .out(tmp02_17_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009226(.in0(tmp01_36_72), .in1(tmp01_37_72), .out(tmp02_18_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009227(.in0(tmp01_38_72), .in1(tmp01_39_72), .out(tmp02_19_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009228(.in0(tmp01_40_72), .in1(tmp01_41_72), .out(tmp02_20_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009229(.in0(tmp01_42_72), .in1(tmp01_43_72), .out(tmp02_21_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009230(.in0(tmp01_44_72), .in1(tmp01_45_72), .out(tmp02_22_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009231(.in0(tmp01_46_72), .in1(tmp01_47_72), .out(tmp02_23_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009232(.in0(tmp01_48_72), .in1(tmp01_49_72), .out(tmp02_24_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009233(.in0(tmp01_50_72), .in1(tmp01_51_72), .out(tmp02_25_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009234(.in0(tmp01_52_72), .in1(tmp01_53_72), .out(tmp02_26_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009235(.in0(tmp01_54_72), .in1(tmp01_55_72), .out(tmp02_27_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009236(.in0(tmp01_56_72), .in1(tmp01_57_72), .out(tmp02_28_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009237(.in0(tmp01_58_72), .in1(tmp01_59_72), .out(tmp02_29_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009238(.in0(tmp01_60_72), .in1(tmp01_61_72), .out(tmp02_30_72));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009239(.in0(tmp01_62_72), .in1(tmp01_63_72), .out(tmp02_31_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009240(.in0(tmp02_0_72), .in1(tmp02_1_72), .out(tmp03_0_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009241(.in0(tmp02_2_72), .in1(tmp02_3_72), .out(tmp03_1_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009242(.in0(tmp02_4_72), .in1(tmp02_5_72), .out(tmp03_2_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009243(.in0(tmp02_6_72), .in1(tmp02_7_72), .out(tmp03_3_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009244(.in0(tmp02_8_72), .in1(tmp02_9_72), .out(tmp03_4_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009245(.in0(tmp02_10_72), .in1(tmp02_11_72), .out(tmp03_5_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009246(.in0(tmp02_12_72), .in1(tmp02_13_72), .out(tmp03_6_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009247(.in0(tmp02_14_72), .in1(tmp02_15_72), .out(tmp03_7_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009248(.in0(tmp02_16_72), .in1(tmp02_17_72), .out(tmp03_8_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009249(.in0(tmp02_18_72), .in1(tmp02_19_72), .out(tmp03_9_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009250(.in0(tmp02_20_72), .in1(tmp02_21_72), .out(tmp03_10_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009251(.in0(tmp02_22_72), .in1(tmp02_23_72), .out(tmp03_11_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009252(.in0(tmp02_24_72), .in1(tmp02_25_72), .out(tmp03_12_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009253(.in0(tmp02_26_72), .in1(tmp02_27_72), .out(tmp03_13_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009254(.in0(tmp02_28_72), .in1(tmp02_29_72), .out(tmp03_14_72));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009255(.in0(tmp02_30_72), .in1(tmp02_31_72), .out(tmp03_15_72));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009256(.in0(tmp03_0_72), .in1(tmp03_1_72), .out(tmp04_0_72));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009257(.in0(tmp03_2_72), .in1(tmp03_3_72), .out(tmp04_1_72));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009258(.in0(tmp03_4_72), .in1(tmp03_5_72), .out(tmp04_2_72));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009259(.in0(tmp03_6_72), .in1(tmp03_7_72), .out(tmp04_3_72));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009260(.in0(tmp03_8_72), .in1(tmp03_9_72), .out(tmp04_4_72));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009261(.in0(tmp03_10_72), .in1(tmp03_11_72), .out(tmp04_5_72));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009262(.in0(tmp03_12_72), .in1(tmp03_13_72), .out(tmp04_6_72));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009263(.in0(tmp03_14_72), .in1(tmp03_15_72), .out(tmp04_7_72));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009264(.in0(tmp04_0_72), .in1(tmp04_1_72), .out(tmp05_0_72));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009265(.in0(tmp04_2_72), .in1(tmp04_3_72), .out(tmp05_1_72));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009266(.in0(tmp04_4_72), .in1(tmp04_5_72), .out(tmp05_2_72));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009267(.in0(tmp04_6_72), .in1(tmp04_7_72), .out(tmp05_3_72));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009268(.in0(tmp05_0_72), .in1(tmp05_1_72), .out(tmp06_0_72));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009269(.in0(tmp05_2_72), .in1(tmp05_3_72), .out(tmp06_1_72));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add009270(.in0(tmp06_0_72), .in1(tmp06_1_72), .out(tmp07_0_72));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009271(.in0(tmp00_0_73), .in1(tmp00_1_73), .out(tmp01_0_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009272(.in0(tmp00_2_73), .in1(tmp00_3_73), .out(tmp01_1_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009273(.in0(tmp00_4_73), .in1(tmp00_5_73), .out(tmp01_2_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009274(.in0(tmp00_6_73), .in1(tmp00_7_73), .out(tmp01_3_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009275(.in0(tmp00_8_73), .in1(tmp00_9_73), .out(tmp01_4_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009276(.in0(tmp00_10_73), .in1(tmp00_11_73), .out(tmp01_5_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009277(.in0(tmp00_12_73), .in1(tmp00_13_73), .out(tmp01_6_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009278(.in0(tmp00_14_73), .in1(tmp00_15_73), .out(tmp01_7_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009279(.in0(tmp00_16_73), .in1(tmp00_17_73), .out(tmp01_8_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009280(.in0(tmp00_18_73), .in1(tmp00_19_73), .out(tmp01_9_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009281(.in0(tmp00_20_73), .in1(tmp00_21_73), .out(tmp01_10_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009282(.in0(tmp00_22_73), .in1(tmp00_23_73), .out(tmp01_11_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009283(.in0(tmp00_24_73), .in1(tmp00_25_73), .out(tmp01_12_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009284(.in0(tmp00_26_73), .in1(tmp00_27_73), .out(tmp01_13_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009285(.in0(tmp00_28_73), .in1(tmp00_29_73), .out(tmp01_14_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009286(.in0(tmp00_30_73), .in1(tmp00_31_73), .out(tmp01_15_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009287(.in0(tmp00_32_73), .in1(tmp00_33_73), .out(tmp01_16_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009288(.in0(tmp00_34_73), .in1(tmp00_35_73), .out(tmp01_17_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009289(.in0(tmp00_36_73), .in1(tmp00_37_73), .out(tmp01_18_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009290(.in0(tmp00_38_73), .in1(tmp00_39_73), .out(tmp01_19_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009291(.in0(tmp00_40_73), .in1(tmp00_41_73), .out(tmp01_20_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009292(.in0(tmp00_42_73), .in1(tmp00_43_73), .out(tmp01_21_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009293(.in0(tmp00_44_73), .in1(tmp00_45_73), .out(tmp01_22_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009294(.in0(tmp00_46_73), .in1(tmp00_47_73), .out(tmp01_23_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009295(.in0(tmp00_48_73), .in1(tmp00_49_73), .out(tmp01_24_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009296(.in0(tmp00_50_73), .in1(tmp00_51_73), .out(tmp01_25_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009297(.in0(tmp00_52_73), .in1(tmp00_53_73), .out(tmp01_26_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009298(.in0(tmp00_54_73), .in1(tmp00_55_73), .out(tmp01_27_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009299(.in0(tmp00_56_73), .in1(tmp00_57_73), .out(tmp01_28_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009300(.in0(tmp00_58_73), .in1(tmp00_59_73), .out(tmp01_29_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009301(.in0(tmp00_60_73), .in1(tmp00_61_73), .out(tmp01_30_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009302(.in0(tmp00_62_73), .in1(tmp00_63_73), .out(tmp01_31_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009303(.in0(tmp00_64_73), .in1(tmp00_65_73), .out(tmp01_32_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009304(.in0(tmp00_66_73), .in1(tmp00_67_73), .out(tmp01_33_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009305(.in0(tmp00_68_73), .in1(tmp00_69_73), .out(tmp01_34_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009306(.in0(tmp00_70_73), .in1(tmp00_71_73), .out(tmp01_35_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009307(.in0(tmp00_72_73), .in1(tmp00_73_73), .out(tmp01_36_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009308(.in0(tmp00_74_73), .in1(tmp00_75_73), .out(tmp01_37_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009309(.in0(tmp00_76_73), .in1(tmp00_77_73), .out(tmp01_38_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009310(.in0(tmp00_78_73), .in1(tmp00_79_73), .out(tmp01_39_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009311(.in0(tmp00_80_73), .in1(tmp00_81_73), .out(tmp01_40_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009312(.in0(tmp00_82_73), .in1(tmp00_83_73), .out(tmp01_41_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009313(.in0(tmp00_84_73), .in1(tmp00_85_73), .out(tmp01_42_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009314(.in0(tmp00_86_73), .in1(tmp00_87_73), .out(tmp01_43_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009315(.in0(tmp00_88_73), .in1(tmp00_89_73), .out(tmp01_44_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009316(.in0(tmp00_90_73), .in1(tmp00_91_73), .out(tmp01_45_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009317(.in0(tmp00_92_73), .in1(tmp00_93_73), .out(tmp01_46_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009318(.in0(tmp00_94_73), .in1(tmp00_95_73), .out(tmp01_47_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009319(.in0(tmp00_96_73), .in1(tmp00_97_73), .out(tmp01_48_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009320(.in0(tmp00_98_73), .in1(tmp00_99_73), .out(tmp01_49_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009321(.in0(tmp00_100_73), .in1(tmp00_101_73), .out(tmp01_50_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009322(.in0(tmp00_102_73), .in1(tmp00_103_73), .out(tmp01_51_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009323(.in0(tmp00_104_73), .in1(tmp00_105_73), .out(tmp01_52_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009324(.in0(tmp00_106_73), .in1(tmp00_107_73), .out(tmp01_53_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009325(.in0(tmp00_108_73), .in1(tmp00_109_73), .out(tmp01_54_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009326(.in0(tmp00_110_73), .in1(tmp00_111_73), .out(tmp01_55_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009327(.in0(tmp00_112_73), .in1(tmp00_113_73), .out(tmp01_56_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009328(.in0(tmp00_114_73), .in1(tmp00_115_73), .out(tmp01_57_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009329(.in0(tmp00_116_73), .in1(tmp00_117_73), .out(tmp01_58_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009330(.in0(tmp00_118_73), .in1(tmp00_119_73), .out(tmp01_59_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009331(.in0(tmp00_120_73), .in1(tmp00_121_73), .out(tmp01_60_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009332(.in0(tmp00_122_73), .in1(tmp00_123_73), .out(tmp01_61_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009333(.in0(tmp00_124_73), .in1(tmp00_125_73), .out(tmp01_62_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009334(.in0(tmp00_126_73), .in1(tmp00_127_73), .out(tmp01_63_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009335(.in0(tmp01_0_73), .in1(tmp01_1_73), .out(tmp02_0_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009336(.in0(tmp01_2_73), .in1(tmp01_3_73), .out(tmp02_1_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009337(.in0(tmp01_4_73), .in1(tmp01_5_73), .out(tmp02_2_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009338(.in0(tmp01_6_73), .in1(tmp01_7_73), .out(tmp02_3_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009339(.in0(tmp01_8_73), .in1(tmp01_9_73), .out(tmp02_4_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009340(.in0(tmp01_10_73), .in1(tmp01_11_73), .out(tmp02_5_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009341(.in0(tmp01_12_73), .in1(tmp01_13_73), .out(tmp02_6_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009342(.in0(tmp01_14_73), .in1(tmp01_15_73), .out(tmp02_7_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009343(.in0(tmp01_16_73), .in1(tmp01_17_73), .out(tmp02_8_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009344(.in0(tmp01_18_73), .in1(tmp01_19_73), .out(tmp02_9_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009345(.in0(tmp01_20_73), .in1(tmp01_21_73), .out(tmp02_10_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009346(.in0(tmp01_22_73), .in1(tmp01_23_73), .out(tmp02_11_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009347(.in0(tmp01_24_73), .in1(tmp01_25_73), .out(tmp02_12_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009348(.in0(tmp01_26_73), .in1(tmp01_27_73), .out(tmp02_13_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009349(.in0(tmp01_28_73), .in1(tmp01_29_73), .out(tmp02_14_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009350(.in0(tmp01_30_73), .in1(tmp01_31_73), .out(tmp02_15_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009351(.in0(tmp01_32_73), .in1(tmp01_33_73), .out(tmp02_16_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009352(.in0(tmp01_34_73), .in1(tmp01_35_73), .out(tmp02_17_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009353(.in0(tmp01_36_73), .in1(tmp01_37_73), .out(tmp02_18_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009354(.in0(tmp01_38_73), .in1(tmp01_39_73), .out(tmp02_19_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009355(.in0(tmp01_40_73), .in1(tmp01_41_73), .out(tmp02_20_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009356(.in0(tmp01_42_73), .in1(tmp01_43_73), .out(tmp02_21_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009357(.in0(tmp01_44_73), .in1(tmp01_45_73), .out(tmp02_22_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009358(.in0(tmp01_46_73), .in1(tmp01_47_73), .out(tmp02_23_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009359(.in0(tmp01_48_73), .in1(tmp01_49_73), .out(tmp02_24_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009360(.in0(tmp01_50_73), .in1(tmp01_51_73), .out(tmp02_25_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009361(.in0(tmp01_52_73), .in1(tmp01_53_73), .out(tmp02_26_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009362(.in0(tmp01_54_73), .in1(tmp01_55_73), .out(tmp02_27_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009363(.in0(tmp01_56_73), .in1(tmp01_57_73), .out(tmp02_28_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009364(.in0(tmp01_58_73), .in1(tmp01_59_73), .out(tmp02_29_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009365(.in0(tmp01_60_73), .in1(tmp01_61_73), .out(tmp02_30_73));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009366(.in0(tmp01_62_73), .in1(tmp01_63_73), .out(tmp02_31_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009367(.in0(tmp02_0_73), .in1(tmp02_1_73), .out(tmp03_0_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009368(.in0(tmp02_2_73), .in1(tmp02_3_73), .out(tmp03_1_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009369(.in0(tmp02_4_73), .in1(tmp02_5_73), .out(tmp03_2_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009370(.in0(tmp02_6_73), .in1(tmp02_7_73), .out(tmp03_3_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009371(.in0(tmp02_8_73), .in1(tmp02_9_73), .out(tmp03_4_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009372(.in0(tmp02_10_73), .in1(tmp02_11_73), .out(tmp03_5_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009373(.in0(tmp02_12_73), .in1(tmp02_13_73), .out(tmp03_6_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009374(.in0(tmp02_14_73), .in1(tmp02_15_73), .out(tmp03_7_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009375(.in0(tmp02_16_73), .in1(tmp02_17_73), .out(tmp03_8_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009376(.in0(tmp02_18_73), .in1(tmp02_19_73), .out(tmp03_9_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009377(.in0(tmp02_20_73), .in1(tmp02_21_73), .out(tmp03_10_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009378(.in0(tmp02_22_73), .in1(tmp02_23_73), .out(tmp03_11_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009379(.in0(tmp02_24_73), .in1(tmp02_25_73), .out(tmp03_12_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009380(.in0(tmp02_26_73), .in1(tmp02_27_73), .out(tmp03_13_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009381(.in0(tmp02_28_73), .in1(tmp02_29_73), .out(tmp03_14_73));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009382(.in0(tmp02_30_73), .in1(tmp02_31_73), .out(tmp03_15_73));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009383(.in0(tmp03_0_73), .in1(tmp03_1_73), .out(tmp04_0_73));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009384(.in0(tmp03_2_73), .in1(tmp03_3_73), .out(tmp04_1_73));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009385(.in0(tmp03_4_73), .in1(tmp03_5_73), .out(tmp04_2_73));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009386(.in0(tmp03_6_73), .in1(tmp03_7_73), .out(tmp04_3_73));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009387(.in0(tmp03_8_73), .in1(tmp03_9_73), .out(tmp04_4_73));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009388(.in0(tmp03_10_73), .in1(tmp03_11_73), .out(tmp04_5_73));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009389(.in0(tmp03_12_73), .in1(tmp03_13_73), .out(tmp04_6_73));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009390(.in0(tmp03_14_73), .in1(tmp03_15_73), .out(tmp04_7_73));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009391(.in0(tmp04_0_73), .in1(tmp04_1_73), .out(tmp05_0_73));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009392(.in0(tmp04_2_73), .in1(tmp04_3_73), .out(tmp05_1_73));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009393(.in0(tmp04_4_73), .in1(tmp04_5_73), .out(tmp05_2_73));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009394(.in0(tmp04_6_73), .in1(tmp04_7_73), .out(tmp05_3_73));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009395(.in0(tmp05_0_73), .in1(tmp05_1_73), .out(tmp06_0_73));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009396(.in0(tmp05_2_73), .in1(tmp05_3_73), .out(tmp06_1_73));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add009397(.in0(tmp06_0_73), .in1(tmp06_1_73), .out(tmp07_0_73));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009398(.in0(tmp00_0_74), .in1(tmp00_1_74), .out(tmp01_0_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009399(.in0(tmp00_2_74), .in1(tmp00_3_74), .out(tmp01_1_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009400(.in0(tmp00_4_74), .in1(tmp00_5_74), .out(tmp01_2_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009401(.in0(tmp00_6_74), .in1(tmp00_7_74), .out(tmp01_3_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009402(.in0(tmp00_8_74), .in1(tmp00_9_74), .out(tmp01_4_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009403(.in0(tmp00_10_74), .in1(tmp00_11_74), .out(tmp01_5_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009404(.in0(tmp00_12_74), .in1(tmp00_13_74), .out(tmp01_6_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009405(.in0(tmp00_14_74), .in1(tmp00_15_74), .out(tmp01_7_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009406(.in0(tmp00_16_74), .in1(tmp00_17_74), .out(tmp01_8_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009407(.in0(tmp00_18_74), .in1(tmp00_19_74), .out(tmp01_9_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009408(.in0(tmp00_20_74), .in1(tmp00_21_74), .out(tmp01_10_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009409(.in0(tmp00_22_74), .in1(tmp00_23_74), .out(tmp01_11_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009410(.in0(tmp00_24_74), .in1(tmp00_25_74), .out(tmp01_12_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009411(.in0(tmp00_26_74), .in1(tmp00_27_74), .out(tmp01_13_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009412(.in0(tmp00_28_74), .in1(tmp00_29_74), .out(tmp01_14_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009413(.in0(tmp00_30_74), .in1(tmp00_31_74), .out(tmp01_15_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009414(.in0(tmp00_32_74), .in1(tmp00_33_74), .out(tmp01_16_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009415(.in0(tmp00_34_74), .in1(tmp00_35_74), .out(tmp01_17_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009416(.in0(tmp00_36_74), .in1(tmp00_37_74), .out(tmp01_18_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009417(.in0(tmp00_38_74), .in1(tmp00_39_74), .out(tmp01_19_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009418(.in0(tmp00_40_74), .in1(tmp00_41_74), .out(tmp01_20_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009419(.in0(tmp00_42_74), .in1(tmp00_43_74), .out(tmp01_21_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009420(.in0(tmp00_44_74), .in1(tmp00_45_74), .out(tmp01_22_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009421(.in0(tmp00_46_74), .in1(tmp00_47_74), .out(tmp01_23_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009422(.in0(tmp00_48_74), .in1(tmp00_49_74), .out(tmp01_24_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009423(.in0(tmp00_50_74), .in1(tmp00_51_74), .out(tmp01_25_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009424(.in0(tmp00_52_74), .in1(tmp00_53_74), .out(tmp01_26_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009425(.in0(tmp00_54_74), .in1(tmp00_55_74), .out(tmp01_27_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009426(.in0(tmp00_56_74), .in1(tmp00_57_74), .out(tmp01_28_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009427(.in0(tmp00_58_74), .in1(tmp00_59_74), .out(tmp01_29_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009428(.in0(tmp00_60_74), .in1(tmp00_61_74), .out(tmp01_30_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009429(.in0(tmp00_62_74), .in1(tmp00_63_74), .out(tmp01_31_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009430(.in0(tmp00_64_74), .in1(tmp00_65_74), .out(tmp01_32_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009431(.in0(tmp00_66_74), .in1(tmp00_67_74), .out(tmp01_33_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009432(.in0(tmp00_68_74), .in1(tmp00_69_74), .out(tmp01_34_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009433(.in0(tmp00_70_74), .in1(tmp00_71_74), .out(tmp01_35_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009434(.in0(tmp00_72_74), .in1(tmp00_73_74), .out(tmp01_36_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009435(.in0(tmp00_74_74), .in1(tmp00_75_74), .out(tmp01_37_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009436(.in0(tmp00_76_74), .in1(tmp00_77_74), .out(tmp01_38_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009437(.in0(tmp00_78_74), .in1(tmp00_79_74), .out(tmp01_39_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009438(.in0(tmp00_80_74), .in1(tmp00_81_74), .out(tmp01_40_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009439(.in0(tmp00_82_74), .in1(tmp00_83_74), .out(tmp01_41_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009440(.in0(tmp00_84_74), .in1(tmp00_85_74), .out(tmp01_42_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009441(.in0(tmp00_86_74), .in1(tmp00_87_74), .out(tmp01_43_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009442(.in0(tmp00_88_74), .in1(tmp00_89_74), .out(tmp01_44_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009443(.in0(tmp00_90_74), .in1(tmp00_91_74), .out(tmp01_45_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009444(.in0(tmp00_92_74), .in1(tmp00_93_74), .out(tmp01_46_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009445(.in0(tmp00_94_74), .in1(tmp00_95_74), .out(tmp01_47_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009446(.in0(tmp00_96_74), .in1(tmp00_97_74), .out(tmp01_48_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009447(.in0(tmp00_98_74), .in1(tmp00_99_74), .out(tmp01_49_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009448(.in0(tmp00_100_74), .in1(tmp00_101_74), .out(tmp01_50_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009449(.in0(tmp00_102_74), .in1(tmp00_103_74), .out(tmp01_51_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009450(.in0(tmp00_104_74), .in1(tmp00_105_74), .out(tmp01_52_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009451(.in0(tmp00_106_74), .in1(tmp00_107_74), .out(tmp01_53_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009452(.in0(tmp00_108_74), .in1(tmp00_109_74), .out(tmp01_54_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009453(.in0(tmp00_110_74), .in1(tmp00_111_74), .out(tmp01_55_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009454(.in0(tmp00_112_74), .in1(tmp00_113_74), .out(tmp01_56_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009455(.in0(tmp00_114_74), .in1(tmp00_115_74), .out(tmp01_57_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009456(.in0(tmp00_116_74), .in1(tmp00_117_74), .out(tmp01_58_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009457(.in0(tmp00_118_74), .in1(tmp00_119_74), .out(tmp01_59_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009458(.in0(tmp00_120_74), .in1(tmp00_121_74), .out(tmp01_60_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009459(.in0(tmp00_122_74), .in1(tmp00_123_74), .out(tmp01_61_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009460(.in0(tmp00_124_74), .in1(tmp00_125_74), .out(tmp01_62_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009461(.in0(tmp00_126_74), .in1(tmp00_127_74), .out(tmp01_63_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009462(.in0(tmp01_0_74), .in1(tmp01_1_74), .out(tmp02_0_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009463(.in0(tmp01_2_74), .in1(tmp01_3_74), .out(tmp02_1_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009464(.in0(tmp01_4_74), .in1(tmp01_5_74), .out(tmp02_2_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009465(.in0(tmp01_6_74), .in1(tmp01_7_74), .out(tmp02_3_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009466(.in0(tmp01_8_74), .in1(tmp01_9_74), .out(tmp02_4_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009467(.in0(tmp01_10_74), .in1(tmp01_11_74), .out(tmp02_5_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009468(.in0(tmp01_12_74), .in1(tmp01_13_74), .out(tmp02_6_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009469(.in0(tmp01_14_74), .in1(tmp01_15_74), .out(tmp02_7_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009470(.in0(tmp01_16_74), .in1(tmp01_17_74), .out(tmp02_8_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009471(.in0(tmp01_18_74), .in1(tmp01_19_74), .out(tmp02_9_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009472(.in0(tmp01_20_74), .in1(tmp01_21_74), .out(tmp02_10_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009473(.in0(tmp01_22_74), .in1(tmp01_23_74), .out(tmp02_11_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009474(.in0(tmp01_24_74), .in1(tmp01_25_74), .out(tmp02_12_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009475(.in0(tmp01_26_74), .in1(tmp01_27_74), .out(tmp02_13_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009476(.in0(tmp01_28_74), .in1(tmp01_29_74), .out(tmp02_14_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009477(.in0(tmp01_30_74), .in1(tmp01_31_74), .out(tmp02_15_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009478(.in0(tmp01_32_74), .in1(tmp01_33_74), .out(tmp02_16_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009479(.in0(tmp01_34_74), .in1(tmp01_35_74), .out(tmp02_17_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009480(.in0(tmp01_36_74), .in1(tmp01_37_74), .out(tmp02_18_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009481(.in0(tmp01_38_74), .in1(tmp01_39_74), .out(tmp02_19_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009482(.in0(tmp01_40_74), .in1(tmp01_41_74), .out(tmp02_20_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009483(.in0(tmp01_42_74), .in1(tmp01_43_74), .out(tmp02_21_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009484(.in0(tmp01_44_74), .in1(tmp01_45_74), .out(tmp02_22_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009485(.in0(tmp01_46_74), .in1(tmp01_47_74), .out(tmp02_23_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009486(.in0(tmp01_48_74), .in1(tmp01_49_74), .out(tmp02_24_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009487(.in0(tmp01_50_74), .in1(tmp01_51_74), .out(tmp02_25_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009488(.in0(tmp01_52_74), .in1(tmp01_53_74), .out(tmp02_26_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009489(.in0(tmp01_54_74), .in1(tmp01_55_74), .out(tmp02_27_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009490(.in0(tmp01_56_74), .in1(tmp01_57_74), .out(tmp02_28_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009491(.in0(tmp01_58_74), .in1(tmp01_59_74), .out(tmp02_29_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009492(.in0(tmp01_60_74), .in1(tmp01_61_74), .out(tmp02_30_74));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009493(.in0(tmp01_62_74), .in1(tmp01_63_74), .out(tmp02_31_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009494(.in0(tmp02_0_74), .in1(tmp02_1_74), .out(tmp03_0_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009495(.in0(tmp02_2_74), .in1(tmp02_3_74), .out(tmp03_1_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009496(.in0(tmp02_4_74), .in1(tmp02_5_74), .out(tmp03_2_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009497(.in0(tmp02_6_74), .in1(tmp02_7_74), .out(tmp03_3_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009498(.in0(tmp02_8_74), .in1(tmp02_9_74), .out(tmp03_4_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009499(.in0(tmp02_10_74), .in1(tmp02_11_74), .out(tmp03_5_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009500(.in0(tmp02_12_74), .in1(tmp02_13_74), .out(tmp03_6_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009501(.in0(tmp02_14_74), .in1(tmp02_15_74), .out(tmp03_7_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009502(.in0(tmp02_16_74), .in1(tmp02_17_74), .out(tmp03_8_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009503(.in0(tmp02_18_74), .in1(tmp02_19_74), .out(tmp03_9_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009504(.in0(tmp02_20_74), .in1(tmp02_21_74), .out(tmp03_10_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009505(.in0(tmp02_22_74), .in1(tmp02_23_74), .out(tmp03_11_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009506(.in0(tmp02_24_74), .in1(tmp02_25_74), .out(tmp03_12_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009507(.in0(tmp02_26_74), .in1(tmp02_27_74), .out(tmp03_13_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009508(.in0(tmp02_28_74), .in1(tmp02_29_74), .out(tmp03_14_74));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009509(.in0(tmp02_30_74), .in1(tmp02_31_74), .out(tmp03_15_74));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009510(.in0(tmp03_0_74), .in1(tmp03_1_74), .out(tmp04_0_74));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009511(.in0(tmp03_2_74), .in1(tmp03_3_74), .out(tmp04_1_74));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009512(.in0(tmp03_4_74), .in1(tmp03_5_74), .out(tmp04_2_74));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009513(.in0(tmp03_6_74), .in1(tmp03_7_74), .out(tmp04_3_74));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009514(.in0(tmp03_8_74), .in1(tmp03_9_74), .out(tmp04_4_74));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009515(.in0(tmp03_10_74), .in1(tmp03_11_74), .out(tmp04_5_74));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009516(.in0(tmp03_12_74), .in1(tmp03_13_74), .out(tmp04_6_74));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009517(.in0(tmp03_14_74), .in1(tmp03_15_74), .out(tmp04_7_74));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009518(.in0(tmp04_0_74), .in1(tmp04_1_74), .out(tmp05_0_74));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009519(.in0(tmp04_2_74), .in1(tmp04_3_74), .out(tmp05_1_74));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009520(.in0(tmp04_4_74), .in1(tmp04_5_74), .out(tmp05_2_74));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009521(.in0(tmp04_6_74), .in1(tmp04_7_74), .out(tmp05_3_74));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009522(.in0(tmp05_0_74), .in1(tmp05_1_74), .out(tmp06_0_74));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009523(.in0(tmp05_2_74), .in1(tmp05_3_74), .out(tmp06_1_74));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add009524(.in0(tmp06_0_74), .in1(tmp06_1_74), .out(tmp07_0_74));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009525(.in0(tmp00_0_75), .in1(tmp00_1_75), .out(tmp01_0_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009526(.in0(tmp00_2_75), .in1(tmp00_3_75), .out(tmp01_1_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009527(.in0(tmp00_4_75), .in1(tmp00_5_75), .out(tmp01_2_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009528(.in0(tmp00_6_75), .in1(tmp00_7_75), .out(tmp01_3_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009529(.in0(tmp00_8_75), .in1(tmp00_9_75), .out(tmp01_4_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009530(.in0(tmp00_10_75), .in1(tmp00_11_75), .out(tmp01_5_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009531(.in0(tmp00_12_75), .in1(tmp00_13_75), .out(tmp01_6_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009532(.in0(tmp00_14_75), .in1(tmp00_15_75), .out(tmp01_7_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009533(.in0(tmp00_16_75), .in1(tmp00_17_75), .out(tmp01_8_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009534(.in0(tmp00_18_75), .in1(tmp00_19_75), .out(tmp01_9_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009535(.in0(tmp00_20_75), .in1(tmp00_21_75), .out(tmp01_10_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009536(.in0(tmp00_22_75), .in1(tmp00_23_75), .out(tmp01_11_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009537(.in0(tmp00_24_75), .in1(tmp00_25_75), .out(tmp01_12_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009538(.in0(tmp00_26_75), .in1(tmp00_27_75), .out(tmp01_13_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009539(.in0(tmp00_28_75), .in1(tmp00_29_75), .out(tmp01_14_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009540(.in0(tmp00_30_75), .in1(tmp00_31_75), .out(tmp01_15_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009541(.in0(tmp00_32_75), .in1(tmp00_33_75), .out(tmp01_16_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009542(.in0(tmp00_34_75), .in1(tmp00_35_75), .out(tmp01_17_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009543(.in0(tmp00_36_75), .in1(tmp00_37_75), .out(tmp01_18_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009544(.in0(tmp00_38_75), .in1(tmp00_39_75), .out(tmp01_19_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009545(.in0(tmp00_40_75), .in1(tmp00_41_75), .out(tmp01_20_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009546(.in0(tmp00_42_75), .in1(tmp00_43_75), .out(tmp01_21_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009547(.in0(tmp00_44_75), .in1(tmp00_45_75), .out(tmp01_22_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009548(.in0(tmp00_46_75), .in1(tmp00_47_75), .out(tmp01_23_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009549(.in0(tmp00_48_75), .in1(tmp00_49_75), .out(tmp01_24_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009550(.in0(tmp00_50_75), .in1(tmp00_51_75), .out(tmp01_25_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009551(.in0(tmp00_52_75), .in1(tmp00_53_75), .out(tmp01_26_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009552(.in0(tmp00_54_75), .in1(tmp00_55_75), .out(tmp01_27_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009553(.in0(tmp00_56_75), .in1(tmp00_57_75), .out(tmp01_28_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009554(.in0(tmp00_58_75), .in1(tmp00_59_75), .out(tmp01_29_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009555(.in0(tmp00_60_75), .in1(tmp00_61_75), .out(tmp01_30_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009556(.in0(tmp00_62_75), .in1(tmp00_63_75), .out(tmp01_31_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009557(.in0(tmp00_64_75), .in1(tmp00_65_75), .out(tmp01_32_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009558(.in0(tmp00_66_75), .in1(tmp00_67_75), .out(tmp01_33_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009559(.in0(tmp00_68_75), .in1(tmp00_69_75), .out(tmp01_34_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009560(.in0(tmp00_70_75), .in1(tmp00_71_75), .out(tmp01_35_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009561(.in0(tmp00_72_75), .in1(tmp00_73_75), .out(tmp01_36_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009562(.in0(tmp00_74_75), .in1(tmp00_75_75), .out(tmp01_37_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009563(.in0(tmp00_76_75), .in1(tmp00_77_75), .out(tmp01_38_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009564(.in0(tmp00_78_75), .in1(tmp00_79_75), .out(tmp01_39_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009565(.in0(tmp00_80_75), .in1(tmp00_81_75), .out(tmp01_40_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009566(.in0(tmp00_82_75), .in1(tmp00_83_75), .out(tmp01_41_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009567(.in0(tmp00_84_75), .in1(tmp00_85_75), .out(tmp01_42_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009568(.in0(tmp00_86_75), .in1(tmp00_87_75), .out(tmp01_43_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009569(.in0(tmp00_88_75), .in1(tmp00_89_75), .out(tmp01_44_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009570(.in0(tmp00_90_75), .in1(tmp00_91_75), .out(tmp01_45_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009571(.in0(tmp00_92_75), .in1(tmp00_93_75), .out(tmp01_46_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009572(.in0(tmp00_94_75), .in1(tmp00_95_75), .out(tmp01_47_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009573(.in0(tmp00_96_75), .in1(tmp00_97_75), .out(tmp01_48_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009574(.in0(tmp00_98_75), .in1(tmp00_99_75), .out(tmp01_49_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009575(.in0(tmp00_100_75), .in1(tmp00_101_75), .out(tmp01_50_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009576(.in0(tmp00_102_75), .in1(tmp00_103_75), .out(tmp01_51_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009577(.in0(tmp00_104_75), .in1(tmp00_105_75), .out(tmp01_52_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009578(.in0(tmp00_106_75), .in1(tmp00_107_75), .out(tmp01_53_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009579(.in0(tmp00_108_75), .in1(tmp00_109_75), .out(tmp01_54_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009580(.in0(tmp00_110_75), .in1(tmp00_111_75), .out(tmp01_55_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009581(.in0(tmp00_112_75), .in1(tmp00_113_75), .out(tmp01_56_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009582(.in0(tmp00_114_75), .in1(tmp00_115_75), .out(tmp01_57_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009583(.in0(tmp00_116_75), .in1(tmp00_117_75), .out(tmp01_58_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009584(.in0(tmp00_118_75), .in1(tmp00_119_75), .out(tmp01_59_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009585(.in0(tmp00_120_75), .in1(tmp00_121_75), .out(tmp01_60_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009586(.in0(tmp00_122_75), .in1(tmp00_123_75), .out(tmp01_61_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009587(.in0(tmp00_124_75), .in1(tmp00_125_75), .out(tmp01_62_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009588(.in0(tmp00_126_75), .in1(tmp00_127_75), .out(tmp01_63_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009589(.in0(tmp01_0_75), .in1(tmp01_1_75), .out(tmp02_0_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009590(.in0(tmp01_2_75), .in1(tmp01_3_75), .out(tmp02_1_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009591(.in0(tmp01_4_75), .in1(tmp01_5_75), .out(tmp02_2_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009592(.in0(tmp01_6_75), .in1(tmp01_7_75), .out(tmp02_3_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009593(.in0(tmp01_8_75), .in1(tmp01_9_75), .out(tmp02_4_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009594(.in0(tmp01_10_75), .in1(tmp01_11_75), .out(tmp02_5_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009595(.in0(tmp01_12_75), .in1(tmp01_13_75), .out(tmp02_6_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009596(.in0(tmp01_14_75), .in1(tmp01_15_75), .out(tmp02_7_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009597(.in0(tmp01_16_75), .in1(tmp01_17_75), .out(tmp02_8_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009598(.in0(tmp01_18_75), .in1(tmp01_19_75), .out(tmp02_9_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009599(.in0(tmp01_20_75), .in1(tmp01_21_75), .out(tmp02_10_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009600(.in0(tmp01_22_75), .in1(tmp01_23_75), .out(tmp02_11_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009601(.in0(tmp01_24_75), .in1(tmp01_25_75), .out(tmp02_12_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009602(.in0(tmp01_26_75), .in1(tmp01_27_75), .out(tmp02_13_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009603(.in0(tmp01_28_75), .in1(tmp01_29_75), .out(tmp02_14_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009604(.in0(tmp01_30_75), .in1(tmp01_31_75), .out(tmp02_15_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009605(.in0(tmp01_32_75), .in1(tmp01_33_75), .out(tmp02_16_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009606(.in0(tmp01_34_75), .in1(tmp01_35_75), .out(tmp02_17_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009607(.in0(tmp01_36_75), .in1(tmp01_37_75), .out(tmp02_18_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009608(.in0(tmp01_38_75), .in1(tmp01_39_75), .out(tmp02_19_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009609(.in0(tmp01_40_75), .in1(tmp01_41_75), .out(tmp02_20_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009610(.in0(tmp01_42_75), .in1(tmp01_43_75), .out(tmp02_21_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009611(.in0(tmp01_44_75), .in1(tmp01_45_75), .out(tmp02_22_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009612(.in0(tmp01_46_75), .in1(tmp01_47_75), .out(tmp02_23_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009613(.in0(tmp01_48_75), .in1(tmp01_49_75), .out(tmp02_24_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009614(.in0(tmp01_50_75), .in1(tmp01_51_75), .out(tmp02_25_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009615(.in0(tmp01_52_75), .in1(tmp01_53_75), .out(tmp02_26_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009616(.in0(tmp01_54_75), .in1(tmp01_55_75), .out(tmp02_27_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009617(.in0(tmp01_56_75), .in1(tmp01_57_75), .out(tmp02_28_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009618(.in0(tmp01_58_75), .in1(tmp01_59_75), .out(tmp02_29_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009619(.in0(tmp01_60_75), .in1(tmp01_61_75), .out(tmp02_30_75));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009620(.in0(tmp01_62_75), .in1(tmp01_63_75), .out(tmp02_31_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009621(.in0(tmp02_0_75), .in1(tmp02_1_75), .out(tmp03_0_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009622(.in0(tmp02_2_75), .in1(tmp02_3_75), .out(tmp03_1_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009623(.in0(tmp02_4_75), .in1(tmp02_5_75), .out(tmp03_2_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009624(.in0(tmp02_6_75), .in1(tmp02_7_75), .out(tmp03_3_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009625(.in0(tmp02_8_75), .in1(tmp02_9_75), .out(tmp03_4_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009626(.in0(tmp02_10_75), .in1(tmp02_11_75), .out(tmp03_5_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009627(.in0(tmp02_12_75), .in1(tmp02_13_75), .out(tmp03_6_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009628(.in0(tmp02_14_75), .in1(tmp02_15_75), .out(tmp03_7_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009629(.in0(tmp02_16_75), .in1(tmp02_17_75), .out(tmp03_8_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009630(.in0(tmp02_18_75), .in1(tmp02_19_75), .out(tmp03_9_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009631(.in0(tmp02_20_75), .in1(tmp02_21_75), .out(tmp03_10_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009632(.in0(tmp02_22_75), .in1(tmp02_23_75), .out(tmp03_11_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009633(.in0(tmp02_24_75), .in1(tmp02_25_75), .out(tmp03_12_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009634(.in0(tmp02_26_75), .in1(tmp02_27_75), .out(tmp03_13_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009635(.in0(tmp02_28_75), .in1(tmp02_29_75), .out(tmp03_14_75));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009636(.in0(tmp02_30_75), .in1(tmp02_31_75), .out(tmp03_15_75));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009637(.in0(tmp03_0_75), .in1(tmp03_1_75), .out(tmp04_0_75));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009638(.in0(tmp03_2_75), .in1(tmp03_3_75), .out(tmp04_1_75));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009639(.in0(tmp03_4_75), .in1(tmp03_5_75), .out(tmp04_2_75));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009640(.in0(tmp03_6_75), .in1(tmp03_7_75), .out(tmp04_3_75));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009641(.in0(tmp03_8_75), .in1(tmp03_9_75), .out(tmp04_4_75));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009642(.in0(tmp03_10_75), .in1(tmp03_11_75), .out(tmp04_5_75));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009643(.in0(tmp03_12_75), .in1(tmp03_13_75), .out(tmp04_6_75));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009644(.in0(tmp03_14_75), .in1(tmp03_15_75), .out(tmp04_7_75));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009645(.in0(tmp04_0_75), .in1(tmp04_1_75), .out(tmp05_0_75));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009646(.in0(tmp04_2_75), .in1(tmp04_3_75), .out(tmp05_1_75));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009647(.in0(tmp04_4_75), .in1(tmp04_5_75), .out(tmp05_2_75));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009648(.in0(tmp04_6_75), .in1(tmp04_7_75), .out(tmp05_3_75));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009649(.in0(tmp05_0_75), .in1(tmp05_1_75), .out(tmp06_0_75));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009650(.in0(tmp05_2_75), .in1(tmp05_3_75), .out(tmp06_1_75));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add009651(.in0(tmp06_0_75), .in1(tmp06_1_75), .out(tmp07_0_75));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009652(.in0(tmp00_0_76), .in1(tmp00_1_76), .out(tmp01_0_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009653(.in0(tmp00_2_76), .in1(tmp00_3_76), .out(tmp01_1_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009654(.in0(tmp00_4_76), .in1(tmp00_5_76), .out(tmp01_2_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009655(.in0(tmp00_6_76), .in1(tmp00_7_76), .out(tmp01_3_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009656(.in0(tmp00_8_76), .in1(tmp00_9_76), .out(tmp01_4_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009657(.in0(tmp00_10_76), .in1(tmp00_11_76), .out(tmp01_5_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009658(.in0(tmp00_12_76), .in1(tmp00_13_76), .out(tmp01_6_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009659(.in0(tmp00_14_76), .in1(tmp00_15_76), .out(tmp01_7_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009660(.in0(tmp00_16_76), .in1(tmp00_17_76), .out(tmp01_8_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009661(.in0(tmp00_18_76), .in1(tmp00_19_76), .out(tmp01_9_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009662(.in0(tmp00_20_76), .in1(tmp00_21_76), .out(tmp01_10_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009663(.in0(tmp00_22_76), .in1(tmp00_23_76), .out(tmp01_11_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009664(.in0(tmp00_24_76), .in1(tmp00_25_76), .out(tmp01_12_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009665(.in0(tmp00_26_76), .in1(tmp00_27_76), .out(tmp01_13_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009666(.in0(tmp00_28_76), .in1(tmp00_29_76), .out(tmp01_14_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009667(.in0(tmp00_30_76), .in1(tmp00_31_76), .out(tmp01_15_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009668(.in0(tmp00_32_76), .in1(tmp00_33_76), .out(tmp01_16_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009669(.in0(tmp00_34_76), .in1(tmp00_35_76), .out(tmp01_17_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009670(.in0(tmp00_36_76), .in1(tmp00_37_76), .out(tmp01_18_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009671(.in0(tmp00_38_76), .in1(tmp00_39_76), .out(tmp01_19_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009672(.in0(tmp00_40_76), .in1(tmp00_41_76), .out(tmp01_20_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009673(.in0(tmp00_42_76), .in1(tmp00_43_76), .out(tmp01_21_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009674(.in0(tmp00_44_76), .in1(tmp00_45_76), .out(tmp01_22_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009675(.in0(tmp00_46_76), .in1(tmp00_47_76), .out(tmp01_23_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009676(.in0(tmp00_48_76), .in1(tmp00_49_76), .out(tmp01_24_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009677(.in0(tmp00_50_76), .in1(tmp00_51_76), .out(tmp01_25_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009678(.in0(tmp00_52_76), .in1(tmp00_53_76), .out(tmp01_26_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009679(.in0(tmp00_54_76), .in1(tmp00_55_76), .out(tmp01_27_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009680(.in0(tmp00_56_76), .in1(tmp00_57_76), .out(tmp01_28_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009681(.in0(tmp00_58_76), .in1(tmp00_59_76), .out(tmp01_29_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009682(.in0(tmp00_60_76), .in1(tmp00_61_76), .out(tmp01_30_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009683(.in0(tmp00_62_76), .in1(tmp00_63_76), .out(tmp01_31_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009684(.in0(tmp00_64_76), .in1(tmp00_65_76), .out(tmp01_32_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009685(.in0(tmp00_66_76), .in1(tmp00_67_76), .out(tmp01_33_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009686(.in0(tmp00_68_76), .in1(tmp00_69_76), .out(tmp01_34_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009687(.in0(tmp00_70_76), .in1(tmp00_71_76), .out(tmp01_35_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009688(.in0(tmp00_72_76), .in1(tmp00_73_76), .out(tmp01_36_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009689(.in0(tmp00_74_76), .in1(tmp00_75_76), .out(tmp01_37_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009690(.in0(tmp00_76_76), .in1(tmp00_77_76), .out(tmp01_38_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009691(.in0(tmp00_78_76), .in1(tmp00_79_76), .out(tmp01_39_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009692(.in0(tmp00_80_76), .in1(tmp00_81_76), .out(tmp01_40_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009693(.in0(tmp00_82_76), .in1(tmp00_83_76), .out(tmp01_41_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009694(.in0(tmp00_84_76), .in1(tmp00_85_76), .out(tmp01_42_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009695(.in0(tmp00_86_76), .in1(tmp00_87_76), .out(tmp01_43_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009696(.in0(tmp00_88_76), .in1(tmp00_89_76), .out(tmp01_44_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009697(.in0(tmp00_90_76), .in1(tmp00_91_76), .out(tmp01_45_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009698(.in0(tmp00_92_76), .in1(tmp00_93_76), .out(tmp01_46_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009699(.in0(tmp00_94_76), .in1(tmp00_95_76), .out(tmp01_47_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009700(.in0(tmp00_96_76), .in1(tmp00_97_76), .out(tmp01_48_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009701(.in0(tmp00_98_76), .in1(tmp00_99_76), .out(tmp01_49_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009702(.in0(tmp00_100_76), .in1(tmp00_101_76), .out(tmp01_50_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009703(.in0(tmp00_102_76), .in1(tmp00_103_76), .out(tmp01_51_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009704(.in0(tmp00_104_76), .in1(tmp00_105_76), .out(tmp01_52_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009705(.in0(tmp00_106_76), .in1(tmp00_107_76), .out(tmp01_53_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009706(.in0(tmp00_108_76), .in1(tmp00_109_76), .out(tmp01_54_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009707(.in0(tmp00_110_76), .in1(tmp00_111_76), .out(tmp01_55_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009708(.in0(tmp00_112_76), .in1(tmp00_113_76), .out(tmp01_56_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009709(.in0(tmp00_114_76), .in1(tmp00_115_76), .out(tmp01_57_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009710(.in0(tmp00_116_76), .in1(tmp00_117_76), .out(tmp01_58_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009711(.in0(tmp00_118_76), .in1(tmp00_119_76), .out(tmp01_59_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009712(.in0(tmp00_120_76), .in1(tmp00_121_76), .out(tmp01_60_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009713(.in0(tmp00_122_76), .in1(tmp00_123_76), .out(tmp01_61_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009714(.in0(tmp00_124_76), .in1(tmp00_125_76), .out(tmp01_62_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009715(.in0(tmp00_126_76), .in1(tmp00_127_76), .out(tmp01_63_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009716(.in0(tmp01_0_76), .in1(tmp01_1_76), .out(tmp02_0_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009717(.in0(tmp01_2_76), .in1(tmp01_3_76), .out(tmp02_1_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009718(.in0(tmp01_4_76), .in1(tmp01_5_76), .out(tmp02_2_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009719(.in0(tmp01_6_76), .in1(tmp01_7_76), .out(tmp02_3_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009720(.in0(tmp01_8_76), .in1(tmp01_9_76), .out(tmp02_4_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009721(.in0(tmp01_10_76), .in1(tmp01_11_76), .out(tmp02_5_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009722(.in0(tmp01_12_76), .in1(tmp01_13_76), .out(tmp02_6_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009723(.in0(tmp01_14_76), .in1(tmp01_15_76), .out(tmp02_7_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009724(.in0(tmp01_16_76), .in1(tmp01_17_76), .out(tmp02_8_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009725(.in0(tmp01_18_76), .in1(tmp01_19_76), .out(tmp02_9_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009726(.in0(tmp01_20_76), .in1(tmp01_21_76), .out(tmp02_10_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009727(.in0(tmp01_22_76), .in1(tmp01_23_76), .out(tmp02_11_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009728(.in0(tmp01_24_76), .in1(tmp01_25_76), .out(tmp02_12_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009729(.in0(tmp01_26_76), .in1(tmp01_27_76), .out(tmp02_13_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009730(.in0(tmp01_28_76), .in1(tmp01_29_76), .out(tmp02_14_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009731(.in0(tmp01_30_76), .in1(tmp01_31_76), .out(tmp02_15_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009732(.in0(tmp01_32_76), .in1(tmp01_33_76), .out(tmp02_16_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009733(.in0(tmp01_34_76), .in1(tmp01_35_76), .out(tmp02_17_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009734(.in0(tmp01_36_76), .in1(tmp01_37_76), .out(tmp02_18_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009735(.in0(tmp01_38_76), .in1(tmp01_39_76), .out(tmp02_19_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009736(.in0(tmp01_40_76), .in1(tmp01_41_76), .out(tmp02_20_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009737(.in0(tmp01_42_76), .in1(tmp01_43_76), .out(tmp02_21_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009738(.in0(tmp01_44_76), .in1(tmp01_45_76), .out(tmp02_22_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009739(.in0(tmp01_46_76), .in1(tmp01_47_76), .out(tmp02_23_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009740(.in0(tmp01_48_76), .in1(tmp01_49_76), .out(tmp02_24_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009741(.in0(tmp01_50_76), .in1(tmp01_51_76), .out(tmp02_25_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009742(.in0(tmp01_52_76), .in1(tmp01_53_76), .out(tmp02_26_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009743(.in0(tmp01_54_76), .in1(tmp01_55_76), .out(tmp02_27_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009744(.in0(tmp01_56_76), .in1(tmp01_57_76), .out(tmp02_28_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009745(.in0(tmp01_58_76), .in1(tmp01_59_76), .out(tmp02_29_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009746(.in0(tmp01_60_76), .in1(tmp01_61_76), .out(tmp02_30_76));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009747(.in0(tmp01_62_76), .in1(tmp01_63_76), .out(tmp02_31_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009748(.in0(tmp02_0_76), .in1(tmp02_1_76), .out(tmp03_0_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009749(.in0(tmp02_2_76), .in1(tmp02_3_76), .out(tmp03_1_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009750(.in0(tmp02_4_76), .in1(tmp02_5_76), .out(tmp03_2_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009751(.in0(tmp02_6_76), .in1(tmp02_7_76), .out(tmp03_3_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009752(.in0(tmp02_8_76), .in1(tmp02_9_76), .out(tmp03_4_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009753(.in0(tmp02_10_76), .in1(tmp02_11_76), .out(tmp03_5_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009754(.in0(tmp02_12_76), .in1(tmp02_13_76), .out(tmp03_6_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009755(.in0(tmp02_14_76), .in1(tmp02_15_76), .out(tmp03_7_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009756(.in0(tmp02_16_76), .in1(tmp02_17_76), .out(tmp03_8_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009757(.in0(tmp02_18_76), .in1(tmp02_19_76), .out(tmp03_9_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009758(.in0(tmp02_20_76), .in1(tmp02_21_76), .out(tmp03_10_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009759(.in0(tmp02_22_76), .in1(tmp02_23_76), .out(tmp03_11_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009760(.in0(tmp02_24_76), .in1(tmp02_25_76), .out(tmp03_12_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009761(.in0(tmp02_26_76), .in1(tmp02_27_76), .out(tmp03_13_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009762(.in0(tmp02_28_76), .in1(tmp02_29_76), .out(tmp03_14_76));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009763(.in0(tmp02_30_76), .in1(tmp02_31_76), .out(tmp03_15_76));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009764(.in0(tmp03_0_76), .in1(tmp03_1_76), .out(tmp04_0_76));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009765(.in0(tmp03_2_76), .in1(tmp03_3_76), .out(tmp04_1_76));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009766(.in0(tmp03_4_76), .in1(tmp03_5_76), .out(tmp04_2_76));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009767(.in0(tmp03_6_76), .in1(tmp03_7_76), .out(tmp04_3_76));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009768(.in0(tmp03_8_76), .in1(tmp03_9_76), .out(tmp04_4_76));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009769(.in0(tmp03_10_76), .in1(tmp03_11_76), .out(tmp04_5_76));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009770(.in0(tmp03_12_76), .in1(tmp03_13_76), .out(tmp04_6_76));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009771(.in0(tmp03_14_76), .in1(tmp03_15_76), .out(tmp04_7_76));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009772(.in0(tmp04_0_76), .in1(tmp04_1_76), .out(tmp05_0_76));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009773(.in0(tmp04_2_76), .in1(tmp04_3_76), .out(tmp05_1_76));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009774(.in0(tmp04_4_76), .in1(tmp04_5_76), .out(tmp05_2_76));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009775(.in0(tmp04_6_76), .in1(tmp04_7_76), .out(tmp05_3_76));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009776(.in0(tmp05_0_76), .in1(tmp05_1_76), .out(tmp06_0_76));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009777(.in0(tmp05_2_76), .in1(tmp05_3_76), .out(tmp06_1_76));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add009778(.in0(tmp06_0_76), .in1(tmp06_1_76), .out(tmp07_0_76));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009779(.in0(tmp00_0_77), .in1(tmp00_1_77), .out(tmp01_0_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009780(.in0(tmp00_2_77), .in1(tmp00_3_77), .out(tmp01_1_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009781(.in0(tmp00_4_77), .in1(tmp00_5_77), .out(tmp01_2_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009782(.in0(tmp00_6_77), .in1(tmp00_7_77), .out(tmp01_3_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009783(.in0(tmp00_8_77), .in1(tmp00_9_77), .out(tmp01_4_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009784(.in0(tmp00_10_77), .in1(tmp00_11_77), .out(tmp01_5_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009785(.in0(tmp00_12_77), .in1(tmp00_13_77), .out(tmp01_6_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009786(.in0(tmp00_14_77), .in1(tmp00_15_77), .out(tmp01_7_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009787(.in0(tmp00_16_77), .in1(tmp00_17_77), .out(tmp01_8_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009788(.in0(tmp00_18_77), .in1(tmp00_19_77), .out(tmp01_9_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009789(.in0(tmp00_20_77), .in1(tmp00_21_77), .out(tmp01_10_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009790(.in0(tmp00_22_77), .in1(tmp00_23_77), .out(tmp01_11_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009791(.in0(tmp00_24_77), .in1(tmp00_25_77), .out(tmp01_12_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009792(.in0(tmp00_26_77), .in1(tmp00_27_77), .out(tmp01_13_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009793(.in0(tmp00_28_77), .in1(tmp00_29_77), .out(tmp01_14_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009794(.in0(tmp00_30_77), .in1(tmp00_31_77), .out(tmp01_15_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009795(.in0(tmp00_32_77), .in1(tmp00_33_77), .out(tmp01_16_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009796(.in0(tmp00_34_77), .in1(tmp00_35_77), .out(tmp01_17_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009797(.in0(tmp00_36_77), .in1(tmp00_37_77), .out(tmp01_18_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009798(.in0(tmp00_38_77), .in1(tmp00_39_77), .out(tmp01_19_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009799(.in0(tmp00_40_77), .in1(tmp00_41_77), .out(tmp01_20_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009800(.in0(tmp00_42_77), .in1(tmp00_43_77), .out(tmp01_21_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009801(.in0(tmp00_44_77), .in1(tmp00_45_77), .out(tmp01_22_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009802(.in0(tmp00_46_77), .in1(tmp00_47_77), .out(tmp01_23_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009803(.in0(tmp00_48_77), .in1(tmp00_49_77), .out(tmp01_24_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009804(.in0(tmp00_50_77), .in1(tmp00_51_77), .out(tmp01_25_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009805(.in0(tmp00_52_77), .in1(tmp00_53_77), .out(tmp01_26_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009806(.in0(tmp00_54_77), .in1(tmp00_55_77), .out(tmp01_27_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009807(.in0(tmp00_56_77), .in1(tmp00_57_77), .out(tmp01_28_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009808(.in0(tmp00_58_77), .in1(tmp00_59_77), .out(tmp01_29_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009809(.in0(tmp00_60_77), .in1(tmp00_61_77), .out(tmp01_30_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009810(.in0(tmp00_62_77), .in1(tmp00_63_77), .out(tmp01_31_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009811(.in0(tmp00_64_77), .in1(tmp00_65_77), .out(tmp01_32_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009812(.in0(tmp00_66_77), .in1(tmp00_67_77), .out(tmp01_33_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009813(.in0(tmp00_68_77), .in1(tmp00_69_77), .out(tmp01_34_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009814(.in0(tmp00_70_77), .in1(tmp00_71_77), .out(tmp01_35_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009815(.in0(tmp00_72_77), .in1(tmp00_73_77), .out(tmp01_36_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009816(.in0(tmp00_74_77), .in1(tmp00_75_77), .out(tmp01_37_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009817(.in0(tmp00_76_77), .in1(tmp00_77_77), .out(tmp01_38_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009818(.in0(tmp00_78_77), .in1(tmp00_79_77), .out(tmp01_39_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009819(.in0(tmp00_80_77), .in1(tmp00_81_77), .out(tmp01_40_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009820(.in0(tmp00_82_77), .in1(tmp00_83_77), .out(tmp01_41_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009821(.in0(tmp00_84_77), .in1(tmp00_85_77), .out(tmp01_42_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009822(.in0(tmp00_86_77), .in1(tmp00_87_77), .out(tmp01_43_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009823(.in0(tmp00_88_77), .in1(tmp00_89_77), .out(tmp01_44_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009824(.in0(tmp00_90_77), .in1(tmp00_91_77), .out(tmp01_45_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009825(.in0(tmp00_92_77), .in1(tmp00_93_77), .out(tmp01_46_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009826(.in0(tmp00_94_77), .in1(tmp00_95_77), .out(tmp01_47_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009827(.in0(tmp00_96_77), .in1(tmp00_97_77), .out(tmp01_48_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009828(.in0(tmp00_98_77), .in1(tmp00_99_77), .out(tmp01_49_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009829(.in0(tmp00_100_77), .in1(tmp00_101_77), .out(tmp01_50_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009830(.in0(tmp00_102_77), .in1(tmp00_103_77), .out(tmp01_51_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009831(.in0(tmp00_104_77), .in1(tmp00_105_77), .out(tmp01_52_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009832(.in0(tmp00_106_77), .in1(tmp00_107_77), .out(tmp01_53_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009833(.in0(tmp00_108_77), .in1(tmp00_109_77), .out(tmp01_54_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009834(.in0(tmp00_110_77), .in1(tmp00_111_77), .out(tmp01_55_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009835(.in0(tmp00_112_77), .in1(tmp00_113_77), .out(tmp01_56_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009836(.in0(tmp00_114_77), .in1(tmp00_115_77), .out(tmp01_57_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009837(.in0(tmp00_116_77), .in1(tmp00_117_77), .out(tmp01_58_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009838(.in0(tmp00_118_77), .in1(tmp00_119_77), .out(tmp01_59_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009839(.in0(tmp00_120_77), .in1(tmp00_121_77), .out(tmp01_60_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009840(.in0(tmp00_122_77), .in1(tmp00_123_77), .out(tmp01_61_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009841(.in0(tmp00_124_77), .in1(tmp00_125_77), .out(tmp01_62_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009842(.in0(tmp00_126_77), .in1(tmp00_127_77), .out(tmp01_63_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009843(.in0(tmp01_0_77), .in1(tmp01_1_77), .out(tmp02_0_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009844(.in0(tmp01_2_77), .in1(tmp01_3_77), .out(tmp02_1_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009845(.in0(tmp01_4_77), .in1(tmp01_5_77), .out(tmp02_2_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009846(.in0(tmp01_6_77), .in1(tmp01_7_77), .out(tmp02_3_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009847(.in0(tmp01_8_77), .in1(tmp01_9_77), .out(tmp02_4_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009848(.in0(tmp01_10_77), .in1(tmp01_11_77), .out(tmp02_5_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009849(.in0(tmp01_12_77), .in1(tmp01_13_77), .out(tmp02_6_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009850(.in0(tmp01_14_77), .in1(tmp01_15_77), .out(tmp02_7_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009851(.in0(tmp01_16_77), .in1(tmp01_17_77), .out(tmp02_8_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009852(.in0(tmp01_18_77), .in1(tmp01_19_77), .out(tmp02_9_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009853(.in0(tmp01_20_77), .in1(tmp01_21_77), .out(tmp02_10_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009854(.in0(tmp01_22_77), .in1(tmp01_23_77), .out(tmp02_11_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009855(.in0(tmp01_24_77), .in1(tmp01_25_77), .out(tmp02_12_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009856(.in0(tmp01_26_77), .in1(tmp01_27_77), .out(tmp02_13_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009857(.in0(tmp01_28_77), .in1(tmp01_29_77), .out(tmp02_14_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009858(.in0(tmp01_30_77), .in1(tmp01_31_77), .out(tmp02_15_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009859(.in0(tmp01_32_77), .in1(tmp01_33_77), .out(tmp02_16_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009860(.in0(tmp01_34_77), .in1(tmp01_35_77), .out(tmp02_17_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009861(.in0(tmp01_36_77), .in1(tmp01_37_77), .out(tmp02_18_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009862(.in0(tmp01_38_77), .in1(tmp01_39_77), .out(tmp02_19_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009863(.in0(tmp01_40_77), .in1(tmp01_41_77), .out(tmp02_20_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009864(.in0(tmp01_42_77), .in1(tmp01_43_77), .out(tmp02_21_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009865(.in0(tmp01_44_77), .in1(tmp01_45_77), .out(tmp02_22_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009866(.in0(tmp01_46_77), .in1(tmp01_47_77), .out(tmp02_23_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009867(.in0(tmp01_48_77), .in1(tmp01_49_77), .out(tmp02_24_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009868(.in0(tmp01_50_77), .in1(tmp01_51_77), .out(tmp02_25_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009869(.in0(tmp01_52_77), .in1(tmp01_53_77), .out(tmp02_26_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009870(.in0(tmp01_54_77), .in1(tmp01_55_77), .out(tmp02_27_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009871(.in0(tmp01_56_77), .in1(tmp01_57_77), .out(tmp02_28_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009872(.in0(tmp01_58_77), .in1(tmp01_59_77), .out(tmp02_29_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009873(.in0(tmp01_60_77), .in1(tmp01_61_77), .out(tmp02_30_77));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009874(.in0(tmp01_62_77), .in1(tmp01_63_77), .out(tmp02_31_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009875(.in0(tmp02_0_77), .in1(tmp02_1_77), .out(tmp03_0_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009876(.in0(tmp02_2_77), .in1(tmp02_3_77), .out(tmp03_1_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009877(.in0(tmp02_4_77), .in1(tmp02_5_77), .out(tmp03_2_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009878(.in0(tmp02_6_77), .in1(tmp02_7_77), .out(tmp03_3_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009879(.in0(tmp02_8_77), .in1(tmp02_9_77), .out(tmp03_4_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009880(.in0(tmp02_10_77), .in1(tmp02_11_77), .out(tmp03_5_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009881(.in0(tmp02_12_77), .in1(tmp02_13_77), .out(tmp03_6_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009882(.in0(tmp02_14_77), .in1(tmp02_15_77), .out(tmp03_7_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009883(.in0(tmp02_16_77), .in1(tmp02_17_77), .out(tmp03_8_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009884(.in0(tmp02_18_77), .in1(tmp02_19_77), .out(tmp03_9_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009885(.in0(tmp02_20_77), .in1(tmp02_21_77), .out(tmp03_10_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009886(.in0(tmp02_22_77), .in1(tmp02_23_77), .out(tmp03_11_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009887(.in0(tmp02_24_77), .in1(tmp02_25_77), .out(tmp03_12_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009888(.in0(tmp02_26_77), .in1(tmp02_27_77), .out(tmp03_13_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009889(.in0(tmp02_28_77), .in1(tmp02_29_77), .out(tmp03_14_77));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add009890(.in0(tmp02_30_77), .in1(tmp02_31_77), .out(tmp03_15_77));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009891(.in0(tmp03_0_77), .in1(tmp03_1_77), .out(tmp04_0_77));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009892(.in0(tmp03_2_77), .in1(tmp03_3_77), .out(tmp04_1_77));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009893(.in0(tmp03_4_77), .in1(tmp03_5_77), .out(tmp04_2_77));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009894(.in0(tmp03_6_77), .in1(tmp03_7_77), .out(tmp04_3_77));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009895(.in0(tmp03_8_77), .in1(tmp03_9_77), .out(tmp04_4_77));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009896(.in0(tmp03_10_77), .in1(tmp03_11_77), .out(tmp04_5_77));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009897(.in0(tmp03_12_77), .in1(tmp03_13_77), .out(tmp04_6_77));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add009898(.in0(tmp03_14_77), .in1(tmp03_15_77), .out(tmp04_7_77));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009899(.in0(tmp04_0_77), .in1(tmp04_1_77), .out(tmp05_0_77));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009900(.in0(tmp04_2_77), .in1(tmp04_3_77), .out(tmp05_1_77));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009901(.in0(tmp04_4_77), .in1(tmp04_5_77), .out(tmp05_2_77));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add009902(.in0(tmp04_6_77), .in1(tmp04_7_77), .out(tmp05_3_77));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009903(.in0(tmp05_0_77), .in1(tmp05_1_77), .out(tmp06_0_77));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add009904(.in0(tmp05_2_77), .in1(tmp05_3_77), .out(tmp06_1_77));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add009905(.in0(tmp06_0_77), .in1(tmp06_1_77), .out(tmp07_0_77));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009906(.in0(tmp00_0_78), .in1(tmp00_1_78), .out(tmp01_0_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009907(.in0(tmp00_2_78), .in1(tmp00_3_78), .out(tmp01_1_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009908(.in0(tmp00_4_78), .in1(tmp00_5_78), .out(tmp01_2_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009909(.in0(tmp00_6_78), .in1(tmp00_7_78), .out(tmp01_3_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009910(.in0(tmp00_8_78), .in1(tmp00_9_78), .out(tmp01_4_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009911(.in0(tmp00_10_78), .in1(tmp00_11_78), .out(tmp01_5_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009912(.in0(tmp00_12_78), .in1(tmp00_13_78), .out(tmp01_6_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009913(.in0(tmp00_14_78), .in1(tmp00_15_78), .out(tmp01_7_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009914(.in0(tmp00_16_78), .in1(tmp00_17_78), .out(tmp01_8_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009915(.in0(tmp00_18_78), .in1(tmp00_19_78), .out(tmp01_9_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009916(.in0(tmp00_20_78), .in1(tmp00_21_78), .out(tmp01_10_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009917(.in0(tmp00_22_78), .in1(tmp00_23_78), .out(tmp01_11_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009918(.in0(tmp00_24_78), .in1(tmp00_25_78), .out(tmp01_12_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009919(.in0(tmp00_26_78), .in1(tmp00_27_78), .out(tmp01_13_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009920(.in0(tmp00_28_78), .in1(tmp00_29_78), .out(tmp01_14_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009921(.in0(tmp00_30_78), .in1(tmp00_31_78), .out(tmp01_15_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009922(.in0(tmp00_32_78), .in1(tmp00_33_78), .out(tmp01_16_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009923(.in0(tmp00_34_78), .in1(tmp00_35_78), .out(tmp01_17_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009924(.in0(tmp00_36_78), .in1(tmp00_37_78), .out(tmp01_18_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009925(.in0(tmp00_38_78), .in1(tmp00_39_78), .out(tmp01_19_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009926(.in0(tmp00_40_78), .in1(tmp00_41_78), .out(tmp01_20_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009927(.in0(tmp00_42_78), .in1(tmp00_43_78), .out(tmp01_21_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009928(.in0(tmp00_44_78), .in1(tmp00_45_78), .out(tmp01_22_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009929(.in0(tmp00_46_78), .in1(tmp00_47_78), .out(tmp01_23_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009930(.in0(tmp00_48_78), .in1(tmp00_49_78), .out(tmp01_24_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009931(.in0(tmp00_50_78), .in1(tmp00_51_78), .out(tmp01_25_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009932(.in0(tmp00_52_78), .in1(tmp00_53_78), .out(tmp01_26_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009933(.in0(tmp00_54_78), .in1(tmp00_55_78), .out(tmp01_27_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009934(.in0(tmp00_56_78), .in1(tmp00_57_78), .out(tmp01_28_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009935(.in0(tmp00_58_78), .in1(tmp00_59_78), .out(tmp01_29_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009936(.in0(tmp00_60_78), .in1(tmp00_61_78), .out(tmp01_30_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009937(.in0(tmp00_62_78), .in1(tmp00_63_78), .out(tmp01_31_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009938(.in0(tmp00_64_78), .in1(tmp00_65_78), .out(tmp01_32_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009939(.in0(tmp00_66_78), .in1(tmp00_67_78), .out(tmp01_33_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009940(.in0(tmp00_68_78), .in1(tmp00_69_78), .out(tmp01_34_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009941(.in0(tmp00_70_78), .in1(tmp00_71_78), .out(tmp01_35_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009942(.in0(tmp00_72_78), .in1(tmp00_73_78), .out(tmp01_36_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009943(.in0(tmp00_74_78), .in1(tmp00_75_78), .out(tmp01_37_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009944(.in0(tmp00_76_78), .in1(tmp00_77_78), .out(tmp01_38_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009945(.in0(tmp00_78_78), .in1(tmp00_79_78), .out(tmp01_39_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009946(.in0(tmp00_80_78), .in1(tmp00_81_78), .out(tmp01_40_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009947(.in0(tmp00_82_78), .in1(tmp00_83_78), .out(tmp01_41_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009948(.in0(tmp00_84_78), .in1(tmp00_85_78), .out(tmp01_42_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009949(.in0(tmp00_86_78), .in1(tmp00_87_78), .out(tmp01_43_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009950(.in0(tmp00_88_78), .in1(tmp00_89_78), .out(tmp01_44_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009951(.in0(tmp00_90_78), .in1(tmp00_91_78), .out(tmp01_45_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009952(.in0(tmp00_92_78), .in1(tmp00_93_78), .out(tmp01_46_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009953(.in0(tmp00_94_78), .in1(tmp00_95_78), .out(tmp01_47_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009954(.in0(tmp00_96_78), .in1(tmp00_97_78), .out(tmp01_48_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009955(.in0(tmp00_98_78), .in1(tmp00_99_78), .out(tmp01_49_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009956(.in0(tmp00_100_78), .in1(tmp00_101_78), .out(tmp01_50_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009957(.in0(tmp00_102_78), .in1(tmp00_103_78), .out(tmp01_51_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009958(.in0(tmp00_104_78), .in1(tmp00_105_78), .out(tmp01_52_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009959(.in0(tmp00_106_78), .in1(tmp00_107_78), .out(tmp01_53_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009960(.in0(tmp00_108_78), .in1(tmp00_109_78), .out(tmp01_54_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009961(.in0(tmp00_110_78), .in1(tmp00_111_78), .out(tmp01_55_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009962(.in0(tmp00_112_78), .in1(tmp00_113_78), .out(tmp01_56_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009963(.in0(tmp00_114_78), .in1(tmp00_115_78), .out(tmp01_57_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009964(.in0(tmp00_116_78), .in1(tmp00_117_78), .out(tmp01_58_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009965(.in0(tmp00_118_78), .in1(tmp00_119_78), .out(tmp01_59_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009966(.in0(tmp00_120_78), .in1(tmp00_121_78), .out(tmp01_60_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009967(.in0(tmp00_122_78), .in1(tmp00_123_78), .out(tmp01_61_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009968(.in0(tmp00_124_78), .in1(tmp00_125_78), .out(tmp01_62_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add009969(.in0(tmp00_126_78), .in1(tmp00_127_78), .out(tmp01_63_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009970(.in0(tmp01_0_78), .in1(tmp01_1_78), .out(tmp02_0_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009971(.in0(tmp01_2_78), .in1(tmp01_3_78), .out(tmp02_1_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009972(.in0(tmp01_4_78), .in1(tmp01_5_78), .out(tmp02_2_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009973(.in0(tmp01_6_78), .in1(tmp01_7_78), .out(tmp02_3_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009974(.in0(tmp01_8_78), .in1(tmp01_9_78), .out(tmp02_4_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009975(.in0(tmp01_10_78), .in1(tmp01_11_78), .out(tmp02_5_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009976(.in0(tmp01_12_78), .in1(tmp01_13_78), .out(tmp02_6_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009977(.in0(tmp01_14_78), .in1(tmp01_15_78), .out(tmp02_7_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009978(.in0(tmp01_16_78), .in1(tmp01_17_78), .out(tmp02_8_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009979(.in0(tmp01_18_78), .in1(tmp01_19_78), .out(tmp02_9_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009980(.in0(tmp01_20_78), .in1(tmp01_21_78), .out(tmp02_10_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009981(.in0(tmp01_22_78), .in1(tmp01_23_78), .out(tmp02_11_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009982(.in0(tmp01_24_78), .in1(tmp01_25_78), .out(tmp02_12_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009983(.in0(tmp01_26_78), .in1(tmp01_27_78), .out(tmp02_13_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009984(.in0(tmp01_28_78), .in1(tmp01_29_78), .out(tmp02_14_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009985(.in0(tmp01_30_78), .in1(tmp01_31_78), .out(tmp02_15_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009986(.in0(tmp01_32_78), .in1(tmp01_33_78), .out(tmp02_16_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009987(.in0(tmp01_34_78), .in1(tmp01_35_78), .out(tmp02_17_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009988(.in0(tmp01_36_78), .in1(tmp01_37_78), .out(tmp02_18_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009989(.in0(tmp01_38_78), .in1(tmp01_39_78), .out(tmp02_19_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009990(.in0(tmp01_40_78), .in1(tmp01_41_78), .out(tmp02_20_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009991(.in0(tmp01_42_78), .in1(tmp01_43_78), .out(tmp02_21_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009992(.in0(tmp01_44_78), .in1(tmp01_45_78), .out(tmp02_22_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009993(.in0(tmp01_46_78), .in1(tmp01_47_78), .out(tmp02_23_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009994(.in0(tmp01_48_78), .in1(tmp01_49_78), .out(tmp02_24_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009995(.in0(tmp01_50_78), .in1(tmp01_51_78), .out(tmp02_25_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009996(.in0(tmp01_52_78), .in1(tmp01_53_78), .out(tmp02_26_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009997(.in0(tmp01_54_78), .in1(tmp01_55_78), .out(tmp02_27_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009998(.in0(tmp01_56_78), .in1(tmp01_57_78), .out(tmp02_28_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add009999(.in0(tmp01_58_78), .in1(tmp01_59_78), .out(tmp02_29_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010000(.in0(tmp01_60_78), .in1(tmp01_61_78), .out(tmp02_30_78));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010001(.in0(tmp01_62_78), .in1(tmp01_63_78), .out(tmp02_31_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010002(.in0(tmp02_0_78), .in1(tmp02_1_78), .out(tmp03_0_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010003(.in0(tmp02_2_78), .in1(tmp02_3_78), .out(tmp03_1_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010004(.in0(tmp02_4_78), .in1(tmp02_5_78), .out(tmp03_2_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010005(.in0(tmp02_6_78), .in1(tmp02_7_78), .out(tmp03_3_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010006(.in0(tmp02_8_78), .in1(tmp02_9_78), .out(tmp03_4_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010007(.in0(tmp02_10_78), .in1(tmp02_11_78), .out(tmp03_5_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010008(.in0(tmp02_12_78), .in1(tmp02_13_78), .out(tmp03_6_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010009(.in0(tmp02_14_78), .in1(tmp02_15_78), .out(tmp03_7_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010010(.in0(tmp02_16_78), .in1(tmp02_17_78), .out(tmp03_8_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010011(.in0(tmp02_18_78), .in1(tmp02_19_78), .out(tmp03_9_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010012(.in0(tmp02_20_78), .in1(tmp02_21_78), .out(tmp03_10_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010013(.in0(tmp02_22_78), .in1(tmp02_23_78), .out(tmp03_11_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010014(.in0(tmp02_24_78), .in1(tmp02_25_78), .out(tmp03_12_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010015(.in0(tmp02_26_78), .in1(tmp02_27_78), .out(tmp03_13_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010016(.in0(tmp02_28_78), .in1(tmp02_29_78), .out(tmp03_14_78));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010017(.in0(tmp02_30_78), .in1(tmp02_31_78), .out(tmp03_15_78));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010018(.in0(tmp03_0_78), .in1(tmp03_1_78), .out(tmp04_0_78));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010019(.in0(tmp03_2_78), .in1(tmp03_3_78), .out(tmp04_1_78));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010020(.in0(tmp03_4_78), .in1(tmp03_5_78), .out(tmp04_2_78));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010021(.in0(tmp03_6_78), .in1(tmp03_7_78), .out(tmp04_3_78));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010022(.in0(tmp03_8_78), .in1(tmp03_9_78), .out(tmp04_4_78));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010023(.in0(tmp03_10_78), .in1(tmp03_11_78), .out(tmp04_5_78));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010024(.in0(tmp03_12_78), .in1(tmp03_13_78), .out(tmp04_6_78));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010025(.in0(tmp03_14_78), .in1(tmp03_15_78), .out(tmp04_7_78));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010026(.in0(tmp04_0_78), .in1(tmp04_1_78), .out(tmp05_0_78));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010027(.in0(tmp04_2_78), .in1(tmp04_3_78), .out(tmp05_1_78));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010028(.in0(tmp04_4_78), .in1(tmp04_5_78), .out(tmp05_2_78));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010029(.in0(tmp04_6_78), .in1(tmp04_7_78), .out(tmp05_3_78));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010030(.in0(tmp05_0_78), .in1(tmp05_1_78), .out(tmp06_0_78));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010031(.in0(tmp05_2_78), .in1(tmp05_3_78), .out(tmp06_1_78));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add010032(.in0(tmp06_0_78), .in1(tmp06_1_78), .out(tmp07_0_78));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010033(.in0(tmp00_0_79), .in1(tmp00_1_79), .out(tmp01_0_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010034(.in0(tmp00_2_79), .in1(tmp00_3_79), .out(tmp01_1_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010035(.in0(tmp00_4_79), .in1(tmp00_5_79), .out(tmp01_2_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010036(.in0(tmp00_6_79), .in1(tmp00_7_79), .out(tmp01_3_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010037(.in0(tmp00_8_79), .in1(tmp00_9_79), .out(tmp01_4_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010038(.in0(tmp00_10_79), .in1(tmp00_11_79), .out(tmp01_5_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010039(.in0(tmp00_12_79), .in1(tmp00_13_79), .out(tmp01_6_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010040(.in0(tmp00_14_79), .in1(tmp00_15_79), .out(tmp01_7_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010041(.in0(tmp00_16_79), .in1(tmp00_17_79), .out(tmp01_8_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010042(.in0(tmp00_18_79), .in1(tmp00_19_79), .out(tmp01_9_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010043(.in0(tmp00_20_79), .in1(tmp00_21_79), .out(tmp01_10_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010044(.in0(tmp00_22_79), .in1(tmp00_23_79), .out(tmp01_11_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010045(.in0(tmp00_24_79), .in1(tmp00_25_79), .out(tmp01_12_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010046(.in0(tmp00_26_79), .in1(tmp00_27_79), .out(tmp01_13_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010047(.in0(tmp00_28_79), .in1(tmp00_29_79), .out(tmp01_14_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010048(.in0(tmp00_30_79), .in1(tmp00_31_79), .out(tmp01_15_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010049(.in0(tmp00_32_79), .in1(tmp00_33_79), .out(tmp01_16_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010050(.in0(tmp00_34_79), .in1(tmp00_35_79), .out(tmp01_17_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010051(.in0(tmp00_36_79), .in1(tmp00_37_79), .out(tmp01_18_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010052(.in0(tmp00_38_79), .in1(tmp00_39_79), .out(tmp01_19_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010053(.in0(tmp00_40_79), .in1(tmp00_41_79), .out(tmp01_20_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010054(.in0(tmp00_42_79), .in1(tmp00_43_79), .out(tmp01_21_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010055(.in0(tmp00_44_79), .in1(tmp00_45_79), .out(tmp01_22_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010056(.in0(tmp00_46_79), .in1(tmp00_47_79), .out(tmp01_23_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010057(.in0(tmp00_48_79), .in1(tmp00_49_79), .out(tmp01_24_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010058(.in0(tmp00_50_79), .in1(tmp00_51_79), .out(tmp01_25_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010059(.in0(tmp00_52_79), .in1(tmp00_53_79), .out(tmp01_26_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010060(.in0(tmp00_54_79), .in1(tmp00_55_79), .out(tmp01_27_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010061(.in0(tmp00_56_79), .in1(tmp00_57_79), .out(tmp01_28_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010062(.in0(tmp00_58_79), .in1(tmp00_59_79), .out(tmp01_29_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010063(.in0(tmp00_60_79), .in1(tmp00_61_79), .out(tmp01_30_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010064(.in0(tmp00_62_79), .in1(tmp00_63_79), .out(tmp01_31_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010065(.in0(tmp00_64_79), .in1(tmp00_65_79), .out(tmp01_32_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010066(.in0(tmp00_66_79), .in1(tmp00_67_79), .out(tmp01_33_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010067(.in0(tmp00_68_79), .in1(tmp00_69_79), .out(tmp01_34_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010068(.in0(tmp00_70_79), .in1(tmp00_71_79), .out(tmp01_35_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010069(.in0(tmp00_72_79), .in1(tmp00_73_79), .out(tmp01_36_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010070(.in0(tmp00_74_79), .in1(tmp00_75_79), .out(tmp01_37_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010071(.in0(tmp00_76_79), .in1(tmp00_77_79), .out(tmp01_38_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010072(.in0(tmp00_78_79), .in1(tmp00_79_79), .out(tmp01_39_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010073(.in0(tmp00_80_79), .in1(tmp00_81_79), .out(tmp01_40_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010074(.in0(tmp00_82_79), .in1(tmp00_83_79), .out(tmp01_41_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010075(.in0(tmp00_84_79), .in1(tmp00_85_79), .out(tmp01_42_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010076(.in0(tmp00_86_79), .in1(tmp00_87_79), .out(tmp01_43_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010077(.in0(tmp00_88_79), .in1(tmp00_89_79), .out(tmp01_44_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010078(.in0(tmp00_90_79), .in1(tmp00_91_79), .out(tmp01_45_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010079(.in0(tmp00_92_79), .in1(tmp00_93_79), .out(tmp01_46_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010080(.in0(tmp00_94_79), .in1(tmp00_95_79), .out(tmp01_47_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010081(.in0(tmp00_96_79), .in1(tmp00_97_79), .out(tmp01_48_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010082(.in0(tmp00_98_79), .in1(tmp00_99_79), .out(tmp01_49_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010083(.in0(tmp00_100_79), .in1(tmp00_101_79), .out(tmp01_50_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010084(.in0(tmp00_102_79), .in1(tmp00_103_79), .out(tmp01_51_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010085(.in0(tmp00_104_79), .in1(tmp00_105_79), .out(tmp01_52_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010086(.in0(tmp00_106_79), .in1(tmp00_107_79), .out(tmp01_53_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010087(.in0(tmp00_108_79), .in1(tmp00_109_79), .out(tmp01_54_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010088(.in0(tmp00_110_79), .in1(tmp00_111_79), .out(tmp01_55_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010089(.in0(tmp00_112_79), .in1(tmp00_113_79), .out(tmp01_56_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010090(.in0(tmp00_114_79), .in1(tmp00_115_79), .out(tmp01_57_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010091(.in0(tmp00_116_79), .in1(tmp00_117_79), .out(tmp01_58_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010092(.in0(tmp00_118_79), .in1(tmp00_119_79), .out(tmp01_59_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010093(.in0(tmp00_120_79), .in1(tmp00_121_79), .out(tmp01_60_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010094(.in0(tmp00_122_79), .in1(tmp00_123_79), .out(tmp01_61_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010095(.in0(tmp00_124_79), .in1(tmp00_125_79), .out(tmp01_62_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010096(.in0(tmp00_126_79), .in1(tmp00_127_79), .out(tmp01_63_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010097(.in0(tmp01_0_79), .in1(tmp01_1_79), .out(tmp02_0_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010098(.in0(tmp01_2_79), .in1(tmp01_3_79), .out(tmp02_1_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010099(.in0(tmp01_4_79), .in1(tmp01_5_79), .out(tmp02_2_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010100(.in0(tmp01_6_79), .in1(tmp01_7_79), .out(tmp02_3_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010101(.in0(tmp01_8_79), .in1(tmp01_9_79), .out(tmp02_4_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010102(.in0(tmp01_10_79), .in1(tmp01_11_79), .out(tmp02_5_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010103(.in0(tmp01_12_79), .in1(tmp01_13_79), .out(tmp02_6_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010104(.in0(tmp01_14_79), .in1(tmp01_15_79), .out(tmp02_7_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010105(.in0(tmp01_16_79), .in1(tmp01_17_79), .out(tmp02_8_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010106(.in0(tmp01_18_79), .in1(tmp01_19_79), .out(tmp02_9_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010107(.in0(tmp01_20_79), .in1(tmp01_21_79), .out(tmp02_10_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010108(.in0(tmp01_22_79), .in1(tmp01_23_79), .out(tmp02_11_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010109(.in0(tmp01_24_79), .in1(tmp01_25_79), .out(tmp02_12_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010110(.in0(tmp01_26_79), .in1(tmp01_27_79), .out(tmp02_13_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010111(.in0(tmp01_28_79), .in1(tmp01_29_79), .out(tmp02_14_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010112(.in0(tmp01_30_79), .in1(tmp01_31_79), .out(tmp02_15_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010113(.in0(tmp01_32_79), .in1(tmp01_33_79), .out(tmp02_16_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010114(.in0(tmp01_34_79), .in1(tmp01_35_79), .out(tmp02_17_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010115(.in0(tmp01_36_79), .in1(tmp01_37_79), .out(tmp02_18_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010116(.in0(tmp01_38_79), .in1(tmp01_39_79), .out(tmp02_19_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010117(.in0(tmp01_40_79), .in1(tmp01_41_79), .out(tmp02_20_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010118(.in0(tmp01_42_79), .in1(tmp01_43_79), .out(tmp02_21_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010119(.in0(tmp01_44_79), .in1(tmp01_45_79), .out(tmp02_22_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010120(.in0(tmp01_46_79), .in1(tmp01_47_79), .out(tmp02_23_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010121(.in0(tmp01_48_79), .in1(tmp01_49_79), .out(tmp02_24_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010122(.in0(tmp01_50_79), .in1(tmp01_51_79), .out(tmp02_25_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010123(.in0(tmp01_52_79), .in1(tmp01_53_79), .out(tmp02_26_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010124(.in0(tmp01_54_79), .in1(tmp01_55_79), .out(tmp02_27_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010125(.in0(tmp01_56_79), .in1(tmp01_57_79), .out(tmp02_28_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010126(.in0(tmp01_58_79), .in1(tmp01_59_79), .out(tmp02_29_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010127(.in0(tmp01_60_79), .in1(tmp01_61_79), .out(tmp02_30_79));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010128(.in0(tmp01_62_79), .in1(tmp01_63_79), .out(tmp02_31_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010129(.in0(tmp02_0_79), .in1(tmp02_1_79), .out(tmp03_0_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010130(.in0(tmp02_2_79), .in1(tmp02_3_79), .out(tmp03_1_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010131(.in0(tmp02_4_79), .in1(tmp02_5_79), .out(tmp03_2_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010132(.in0(tmp02_6_79), .in1(tmp02_7_79), .out(tmp03_3_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010133(.in0(tmp02_8_79), .in1(tmp02_9_79), .out(tmp03_4_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010134(.in0(tmp02_10_79), .in1(tmp02_11_79), .out(tmp03_5_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010135(.in0(tmp02_12_79), .in1(tmp02_13_79), .out(tmp03_6_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010136(.in0(tmp02_14_79), .in1(tmp02_15_79), .out(tmp03_7_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010137(.in0(tmp02_16_79), .in1(tmp02_17_79), .out(tmp03_8_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010138(.in0(tmp02_18_79), .in1(tmp02_19_79), .out(tmp03_9_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010139(.in0(tmp02_20_79), .in1(tmp02_21_79), .out(tmp03_10_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010140(.in0(tmp02_22_79), .in1(tmp02_23_79), .out(tmp03_11_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010141(.in0(tmp02_24_79), .in1(tmp02_25_79), .out(tmp03_12_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010142(.in0(tmp02_26_79), .in1(tmp02_27_79), .out(tmp03_13_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010143(.in0(tmp02_28_79), .in1(tmp02_29_79), .out(tmp03_14_79));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010144(.in0(tmp02_30_79), .in1(tmp02_31_79), .out(tmp03_15_79));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010145(.in0(tmp03_0_79), .in1(tmp03_1_79), .out(tmp04_0_79));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010146(.in0(tmp03_2_79), .in1(tmp03_3_79), .out(tmp04_1_79));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010147(.in0(tmp03_4_79), .in1(tmp03_5_79), .out(tmp04_2_79));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010148(.in0(tmp03_6_79), .in1(tmp03_7_79), .out(tmp04_3_79));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010149(.in0(tmp03_8_79), .in1(tmp03_9_79), .out(tmp04_4_79));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010150(.in0(tmp03_10_79), .in1(tmp03_11_79), .out(tmp04_5_79));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010151(.in0(tmp03_12_79), .in1(tmp03_13_79), .out(tmp04_6_79));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010152(.in0(tmp03_14_79), .in1(tmp03_15_79), .out(tmp04_7_79));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010153(.in0(tmp04_0_79), .in1(tmp04_1_79), .out(tmp05_0_79));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010154(.in0(tmp04_2_79), .in1(tmp04_3_79), .out(tmp05_1_79));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010155(.in0(tmp04_4_79), .in1(tmp04_5_79), .out(tmp05_2_79));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010156(.in0(tmp04_6_79), .in1(tmp04_7_79), .out(tmp05_3_79));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010157(.in0(tmp05_0_79), .in1(tmp05_1_79), .out(tmp06_0_79));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010158(.in0(tmp05_2_79), .in1(tmp05_3_79), .out(tmp06_1_79));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add010159(.in0(tmp06_0_79), .in1(tmp06_1_79), .out(tmp07_0_79));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010160(.in0(tmp00_0_80), .in1(tmp00_1_80), .out(tmp01_0_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010161(.in0(tmp00_2_80), .in1(tmp00_3_80), .out(tmp01_1_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010162(.in0(tmp00_4_80), .in1(tmp00_5_80), .out(tmp01_2_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010163(.in0(tmp00_6_80), .in1(tmp00_7_80), .out(tmp01_3_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010164(.in0(tmp00_8_80), .in1(tmp00_9_80), .out(tmp01_4_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010165(.in0(tmp00_10_80), .in1(tmp00_11_80), .out(tmp01_5_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010166(.in0(tmp00_12_80), .in1(tmp00_13_80), .out(tmp01_6_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010167(.in0(tmp00_14_80), .in1(tmp00_15_80), .out(tmp01_7_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010168(.in0(tmp00_16_80), .in1(tmp00_17_80), .out(tmp01_8_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010169(.in0(tmp00_18_80), .in1(tmp00_19_80), .out(tmp01_9_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010170(.in0(tmp00_20_80), .in1(tmp00_21_80), .out(tmp01_10_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010171(.in0(tmp00_22_80), .in1(tmp00_23_80), .out(tmp01_11_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010172(.in0(tmp00_24_80), .in1(tmp00_25_80), .out(tmp01_12_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010173(.in0(tmp00_26_80), .in1(tmp00_27_80), .out(tmp01_13_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010174(.in0(tmp00_28_80), .in1(tmp00_29_80), .out(tmp01_14_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010175(.in0(tmp00_30_80), .in1(tmp00_31_80), .out(tmp01_15_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010176(.in0(tmp00_32_80), .in1(tmp00_33_80), .out(tmp01_16_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010177(.in0(tmp00_34_80), .in1(tmp00_35_80), .out(tmp01_17_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010178(.in0(tmp00_36_80), .in1(tmp00_37_80), .out(tmp01_18_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010179(.in0(tmp00_38_80), .in1(tmp00_39_80), .out(tmp01_19_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010180(.in0(tmp00_40_80), .in1(tmp00_41_80), .out(tmp01_20_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010181(.in0(tmp00_42_80), .in1(tmp00_43_80), .out(tmp01_21_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010182(.in0(tmp00_44_80), .in1(tmp00_45_80), .out(tmp01_22_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010183(.in0(tmp00_46_80), .in1(tmp00_47_80), .out(tmp01_23_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010184(.in0(tmp00_48_80), .in1(tmp00_49_80), .out(tmp01_24_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010185(.in0(tmp00_50_80), .in1(tmp00_51_80), .out(tmp01_25_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010186(.in0(tmp00_52_80), .in1(tmp00_53_80), .out(tmp01_26_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010187(.in0(tmp00_54_80), .in1(tmp00_55_80), .out(tmp01_27_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010188(.in0(tmp00_56_80), .in1(tmp00_57_80), .out(tmp01_28_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010189(.in0(tmp00_58_80), .in1(tmp00_59_80), .out(tmp01_29_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010190(.in0(tmp00_60_80), .in1(tmp00_61_80), .out(tmp01_30_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010191(.in0(tmp00_62_80), .in1(tmp00_63_80), .out(tmp01_31_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010192(.in0(tmp00_64_80), .in1(tmp00_65_80), .out(tmp01_32_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010193(.in0(tmp00_66_80), .in1(tmp00_67_80), .out(tmp01_33_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010194(.in0(tmp00_68_80), .in1(tmp00_69_80), .out(tmp01_34_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010195(.in0(tmp00_70_80), .in1(tmp00_71_80), .out(tmp01_35_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010196(.in0(tmp00_72_80), .in1(tmp00_73_80), .out(tmp01_36_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010197(.in0(tmp00_74_80), .in1(tmp00_75_80), .out(tmp01_37_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010198(.in0(tmp00_76_80), .in1(tmp00_77_80), .out(tmp01_38_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010199(.in0(tmp00_78_80), .in1(tmp00_79_80), .out(tmp01_39_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010200(.in0(tmp00_80_80), .in1(tmp00_81_80), .out(tmp01_40_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010201(.in0(tmp00_82_80), .in1(tmp00_83_80), .out(tmp01_41_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010202(.in0(tmp00_84_80), .in1(tmp00_85_80), .out(tmp01_42_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010203(.in0(tmp00_86_80), .in1(tmp00_87_80), .out(tmp01_43_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010204(.in0(tmp00_88_80), .in1(tmp00_89_80), .out(tmp01_44_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010205(.in0(tmp00_90_80), .in1(tmp00_91_80), .out(tmp01_45_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010206(.in0(tmp00_92_80), .in1(tmp00_93_80), .out(tmp01_46_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010207(.in0(tmp00_94_80), .in1(tmp00_95_80), .out(tmp01_47_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010208(.in0(tmp00_96_80), .in1(tmp00_97_80), .out(tmp01_48_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010209(.in0(tmp00_98_80), .in1(tmp00_99_80), .out(tmp01_49_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010210(.in0(tmp00_100_80), .in1(tmp00_101_80), .out(tmp01_50_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010211(.in0(tmp00_102_80), .in1(tmp00_103_80), .out(tmp01_51_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010212(.in0(tmp00_104_80), .in1(tmp00_105_80), .out(tmp01_52_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010213(.in0(tmp00_106_80), .in1(tmp00_107_80), .out(tmp01_53_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010214(.in0(tmp00_108_80), .in1(tmp00_109_80), .out(tmp01_54_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010215(.in0(tmp00_110_80), .in1(tmp00_111_80), .out(tmp01_55_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010216(.in0(tmp00_112_80), .in1(tmp00_113_80), .out(tmp01_56_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010217(.in0(tmp00_114_80), .in1(tmp00_115_80), .out(tmp01_57_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010218(.in0(tmp00_116_80), .in1(tmp00_117_80), .out(tmp01_58_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010219(.in0(tmp00_118_80), .in1(tmp00_119_80), .out(tmp01_59_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010220(.in0(tmp00_120_80), .in1(tmp00_121_80), .out(tmp01_60_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010221(.in0(tmp00_122_80), .in1(tmp00_123_80), .out(tmp01_61_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010222(.in0(tmp00_124_80), .in1(tmp00_125_80), .out(tmp01_62_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010223(.in0(tmp00_126_80), .in1(tmp00_127_80), .out(tmp01_63_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010224(.in0(tmp01_0_80), .in1(tmp01_1_80), .out(tmp02_0_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010225(.in0(tmp01_2_80), .in1(tmp01_3_80), .out(tmp02_1_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010226(.in0(tmp01_4_80), .in1(tmp01_5_80), .out(tmp02_2_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010227(.in0(tmp01_6_80), .in1(tmp01_7_80), .out(tmp02_3_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010228(.in0(tmp01_8_80), .in1(tmp01_9_80), .out(tmp02_4_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010229(.in0(tmp01_10_80), .in1(tmp01_11_80), .out(tmp02_5_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010230(.in0(tmp01_12_80), .in1(tmp01_13_80), .out(tmp02_6_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010231(.in0(tmp01_14_80), .in1(tmp01_15_80), .out(tmp02_7_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010232(.in0(tmp01_16_80), .in1(tmp01_17_80), .out(tmp02_8_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010233(.in0(tmp01_18_80), .in1(tmp01_19_80), .out(tmp02_9_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010234(.in0(tmp01_20_80), .in1(tmp01_21_80), .out(tmp02_10_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010235(.in0(tmp01_22_80), .in1(tmp01_23_80), .out(tmp02_11_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010236(.in0(tmp01_24_80), .in1(tmp01_25_80), .out(tmp02_12_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010237(.in0(tmp01_26_80), .in1(tmp01_27_80), .out(tmp02_13_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010238(.in0(tmp01_28_80), .in1(tmp01_29_80), .out(tmp02_14_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010239(.in0(tmp01_30_80), .in1(tmp01_31_80), .out(tmp02_15_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010240(.in0(tmp01_32_80), .in1(tmp01_33_80), .out(tmp02_16_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010241(.in0(tmp01_34_80), .in1(tmp01_35_80), .out(tmp02_17_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010242(.in0(tmp01_36_80), .in1(tmp01_37_80), .out(tmp02_18_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010243(.in0(tmp01_38_80), .in1(tmp01_39_80), .out(tmp02_19_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010244(.in0(tmp01_40_80), .in1(tmp01_41_80), .out(tmp02_20_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010245(.in0(tmp01_42_80), .in1(tmp01_43_80), .out(tmp02_21_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010246(.in0(tmp01_44_80), .in1(tmp01_45_80), .out(tmp02_22_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010247(.in0(tmp01_46_80), .in1(tmp01_47_80), .out(tmp02_23_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010248(.in0(tmp01_48_80), .in1(tmp01_49_80), .out(tmp02_24_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010249(.in0(tmp01_50_80), .in1(tmp01_51_80), .out(tmp02_25_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010250(.in0(tmp01_52_80), .in1(tmp01_53_80), .out(tmp02_26_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010251(.in0(tmp01_54_80), .in1(tmp01_55_80), .out(tmp02_27_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010252(.in0(tmp01_56_80), .in1(tmp01_57_80), .out(tmp02_28_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010253(.in0(tmp01_58_80), .in1(tmp01_59_80), .out(tmp02_29_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010254(.in0(tmp01_60_80), .in1(tmp01_61_80), .out(tmp02_30_80));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010255(.in0(tmp01_62_80), .in1(tmp01_63_80), .out(tmp02_31_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010256(.in0(tmp02_0_80), .in1(tmp02_1_80), .out(tmp03_0_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010257(.in0(tmp02_2_80), .in1(tmp02_3_80), .out(tmp03_1_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010258(.in0(tmp02_4_80), .in1(tmp02_5_80), .out(tmp03_2_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010259(.in0(tmp02_6_80), .in1(tmp02_7_80), .out(tmp03_3_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010260(.in0(tmp02_8_80), .in1(tmp02_9_80), .out(tmp03_4_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010261(.in0(tmp02_10_80), .in1(tmp02_11_80), .out(tmp03_5_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010262(.in0(tmp02_12_80), .in1(tmp02_13_80), .out(tmp03_6_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010263(.in0(tmp02_14_80), .in1(tmp02_15_80), .out(tmp03_7_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010264(.in0(tmp02_16_80), .in1(tmp02_17_80), .out(tmp03_8_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010265(.in0(tmp02_18_80), .in1(tmp02_19_80), .out(tmp03_9_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010266(.in0(tmp02_20_80), .in1(tmp02_21_80), .out(tmp03_10_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010267(.in0(tmp02_22_80), .in1(tmp02_23_80), .out(tmp03_11_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010268(.in0(tmp02_24_80), .in1(tmp02_25_80), .out(tmp03_12_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010269(.in0(tmp02_26_80), .in1(tmp02_27_80), .out(tmp03_13_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010270(.in0(tmp02_28_80), .in1(tmp02_29_80), .out(tmp03_14_80));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010271(.in0(tmp02_30_80), .in1(tmp02_31_80), .out(tmp03_15_80));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010272(.in0(tmp03_0_80), .in1(tmp03_1_80), .out(tmp04_0_80));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010273(.in0(tmp03_2_80), .in1(tmp03_3_80), .out(tmp04_1_80));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010274(.in0(tmp03_4_80), .in1(tmp03_5_80), .out(tmp04_2_80));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010275(.in0(tmp03_6_80), .in1(tmp03_7_80), .out(tmp04_3_80));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010276(.in0(tmp03_8_80), .in1(tmp03_9_80), .out(tmp04_4_80));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010277(.in0(tmp03_10_80), .in1(tmp03_11_80), .out(tmp04_5_80));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010278(.in0(tmp03_12_80), .in1(tmp03_13_80), .out(tmp04_6_80));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010279(.in0(tmp03_14_80), .in1(tmp03_15_80), .out(tmp04_7_80));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010280(.in0(tmp04_0_80), .in1(tmp04_1_80), .out(tmp05_0_80));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010281(.in0(tmp04_2_80), .in1(tmp04_3_80), .out(tmp05_1_80));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010282(.in0(tmp04_4_80), .in1(tmp04_5_80), .out(tmp05_2_80));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010283(.in0(tmp04_6_80), .in1(tmp04_7_80), .out(tmp05_3_80));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010284(.in0(tmp05_0_80), .in1(tmp05_1_80), .out(tmp06_0_80));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010285(.in0(tmp05_2_80), .in1(tmp05_3_80), .out(tmp06_1_80));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add010286(.in0(tmp06_0_80), .in1(tmp06_1_80), .out(tmp07_0_80));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010287(.in0(tmp00_0_81), .in1(tmp00_1_81), .out(tmp01_0_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010288(.in0(tmp00_2_81), .in1(tmp00_3_81), .out(tmp01_1_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010289(.in0(tmp00_4_81), .in1(tmp00_5_81), .out(tmp01_2_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010290(.in0(tmp00_6_81), .in1(tmp00_7_81), .out(tmp01_3_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010291(.in0(tmp00_8_81), .in1(tmp00_9_81), .out(tmp01_4_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010292(.in0(tmp00_10_81), .in1(tmp00_11_81), .out(tmp01_5_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010293(.in0(tmp00_12_81), .in1(tmp00_13_81), .out(tmp01_6_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010294(.in0(tmp00_14_81), .in1(tmp00_15_81), .out(tmp01_7_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010295(.in0(tmp00_16_81), .in1(tmp00_17_81), .out(tmp01_8_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010296(.in0(tmp00_18_81), .in1(tmp00_19_81), .out(tmp01_9_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010297(.in0(tmp00_20_81), .in1(tmp00_21_81), .out(tmp01_10_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010298(.in0(tmp00_22_81), .in1(tmp00_23_81), .out(tmp01_11_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010299(.in0(tmp00_24_81), .in1(tmp00_25_81), .out(tmp01_12_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010300(.in0(tmp00_26_81), .in1(tmp00_27_81), .out(tmp01_13_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010301(.in0(tmp00_28_81), .in1(tmp00_29_81), .out(tmp01_14_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010302(.in0(tmp00_30_81), .in1(tmp00_31_81), .out(tmp01_15_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010303(.in0(tmp00_32_81), .in1(tmp00_33_81), .out(tmp01_16_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010304(.in0(tmp00_34_81), .in1(tmp00_35_81), .out(tmp01_17_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010305(.in0(tmp00_36_81), .in1(tmp00_37_81), .out(tmp01_18_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010306(.in0(tmp00_38_81), .in1(tmp00_39_81), .out(tmp01_19_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010307(.in0(tmp00_40_81), .in1(tmp00_41_81), .out(tmp01_20_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010308(.in0(tmp00_42_81), .in1(tmp00_43_81), .out(tmp01_21_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010309(.in0(tmp00_44_81), .in1(tmp00_45_81), .out(tmp01_22_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010310(.in0(tmp00_46_81), .in1(tmp00_47_81), .out(tmp01_23_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010311(.in0(tmp00_48_81), .in1(tmp00_49_81), .out(tmp01_24_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010312(.in0(tmp00_50_81), .in1(tmp00_51_81), .out(tmp01_25_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010313(.in0(tmp00_52_81), .in1(tmp00_53_81), .out(tmp01_26_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010314(.in0(tmp00_54_81), .in1(tmp00_55_81), .out(tmp01_27_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010315(.in0(tmp00_56_81), .in1(tmp00_57_81), .out(tmp01_28_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010316(.in0(tmp00_58_81), .in1(tmp00_59_81), .out(tmp01_29_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010317(.in0(tmp00_60_81), .in1(tmp00_61_81), .out(tmp01_30_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010318(.in0(tmp00_62_81), .in1(tmp00_63_81), .out(tmp01_31_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010319(.in0(tmp00_64_81), .in1(tmp00_65_81), .out(tmp01_32_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010320(.in0(tmp00_66_81), .in1(tmp00_67_81), .out(tmp01_33_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010321(.in0(tmp00_68_81), .in1(tmp00_69_81), .out(tmp01_34_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010322(.in0(tmp00_70_81), .in1(tmp00_71_81), .out(tmp01_35_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010323(.in0(tmp00_72_81), .in1(tmp00_73_81), .out(tmp01_36_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010324(.in0(tmp00_74_81), .in1(tmp00_75_81), .out(tmp01_37_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010325(.in0(tmp00_76_81), .in1(tmp00_77_81), .out(tmp01_38_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010326(.in0(tmp00_78_81), .in1(tmp00_79_81), .out(tmp01_39_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010327(.in0(tmp00_80_81), .in1(tmp00_81_81), .out(tmp01_40_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010328(.in0(tmp00_82_81), .in1(tmp00_83_81), .out(tmp01_41_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010329(.in0(tmp00_84_81), .in1(tmp00_85_81), .out(tmp01_42_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010330(.in0(tmp00_86_81), .in1(tmp00_87_81), .out(tmp01_43_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010331(.in0(tmp00_88_81), .in1(tmp00_89_81), .out(tmp01_44_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010332(.in0(tmp00_90_81), .in1(tmp00_91_81), .out(tmp01_45_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010333(.in0(tmp00_92_81), .in1(tmp00_93_81), .out(tmp01_46_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010334(.in0(tmp00_94_81), .in1(tmp00_95_81), .out(tmp01_47_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010335(.in0(tmp00_96_81), .in1(tmp00_97_81), .out(tmp01_48_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010336(.in0(tmp00_98_81), .in1(tmp00_99_81), .out(tmp01_49_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010337(.in0(tmp00_100_81), .in1(tmp00_101_81), .out(tmp01_50_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010338(.in0(tmp00_102_81), .in1(tmp00_103_81), .out(tmp01_51_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010339(.in0(tmp00_104_81), .in1(tmp00_105_81), .out(tmp01_52_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010340(.in0(tmp00_106_81), .in1(tmp00_107_81), .out(tmp01_53_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010341(.in0(tmp00_108_81), .in1(tmp00_109_81), .out(tmp01_54_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010342(.in0(tmp00_110_81), .in1(tmp00_111_81), .out(tmp01_55_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010343(.in0(tmp00_112_81), .in1(tmp00_113_81), .out(tmp01_56_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010344(.in0(tmp00_114_81), .in1(tmp00_115_81), .out(tmp01_57_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010345(.in0(tmp00_116_81), .in1(tmp00_117_81), .out(tmp01_58_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010346(.in0(tmp00_118_81), .in1(tmp00_119_81), .out(tmp01_59_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010347(.in0(tmp00_120_81), .in1(tmp00_121_81), .out(tmp01_60_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010348(.in0(tmp00_122_81), .in1(tmp00_123_81), .out(tmp01_61_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010349(.in0(tmp00_124_81), .in1(tmp00_125_81), .out(tmp01_62_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010350(.in0(tmp00_126_81), .in1(tmp00_127_81), .out(tmp01_63_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010351(.in0(tmp01_0_81), .in1(tmp01_1_81), .out(tmp02_0_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010352(.in0(tmp01_2_81), .in1(tmp01_3_81), .out(tmp02_1_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010353(.in0(tmp01_4_81), .in1(tmp01_5_81), .out(tmp02_2_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010354(.in0(tmp01_6_81), .in1(tmp01_7_81), .out(tmp02_3_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010355(.in0(tmp01_8_81), .in1(tmp01_9_81), .out(tmp02_4_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010356(.in0(tmp01_10_81), .in1(tmp01_11_81), .out(tmp02_5_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010357(.in0(tmp01_12_81), .in1(tmp01_13_81), .out(tmp02_6_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010358(.in0(tmp01_14_81), .in1(tmp01_15_81), .out(tmp02_7_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010359(.in0(tmp01_16_81), .in1(tmp01_17_81), .out(tmp02_8_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010360(.in0(tmp01_18_81), .in1(tmp01_19_81), .out(tmp02_9_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010361(.in0(tmp01_20_81), .in1(tmp01_21_81), .out(tmp02_10_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010362(.in0(tmp01_22_81), .in1(tmp01_23_81), .out(tmp02_11_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010363(.in0(tmp01_24_81), .in1(tmp01_25_81), .out(tmp02_12_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010364(.in0(tmp01_26_81), .in1(tmp01_27_81), .out(tmp02_13_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010365(.in0(tmp01_28_81), .in1(tmp01_29_81), .out(tmp02_14_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010366(.in0(tmp01_30_81), .in1(tmp01_31_81), .out(tmp02_15_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010367(.in0(tmp01_32_81), .in1(tmp01_33_81), .out(tmp02_16_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010368(.in0(tmp01_34_81), .in1(tmp01_35_81), .out(tmp02_17_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010369(.in0(tmp01_36_81), .in1(tmp01_37_81), .out(tmp02_18_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010370(.in0(tmp01_38_81), .in1(tmp01_39_81), .out(tmp02_19_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010371(.in0(tmp01_40_81), .in1(tmp01_41_81), .out(tmp02_20_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010372(.in0(tmp01_42_81), .in1(tmp01_43_81), .out(tmp02_21_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010373(.in0(tmp01_44_81), .in1(tmp01_45_81), .out(tmp02_22_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010374(.in0(tmp01_46_81), .in1(tmp01_47_81), .out(tmp02_23_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010375(.in0(tmp01_48_81), .in1(tmp01_49_81), .out(tmp02_24_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010376(.in0(tmp01_50_81), .in1(tmp01_51_81), .out(tmp02_25_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010377(.in0(tmp01_52_81), .in1(tmp01_53_81), .out(tmp02_26_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010378(.in0(tmp01_54_81), .in1(tmp01_55_81), .out(tmp02_27_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010379(.in0(tmp01_56_81), .in1(tmp01_57_81), .out(tmp02_28_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010380(.in0(tmp01_58_81), .in1(tmp01_59_81), .out(tmp02_29_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010381(.in0(tmp01_60_81), .in1(tmp01_61_81), .out(tmp02_30_81));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010382(.in0(tmp01_62_81), .in1(tmp01_63_81), .out(tmp02_31_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010383(.in0(tmp02_0_81), .in1(tmp02_1_81), .out(tmp03_0_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010384(.in0(tmp02_2_81), .in1(tmp02_3_81), .out(tmp03_1_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010385(.in0(tmp02_4_81), .in1(tmp02_5_81), .out(tmp03_2_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010386(.in0(tmp02_6_81), .in1(tmp02_7_81), .out(tmp03_3_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010387(.in0(tmp02_8_81), .in1(tmp02_9_81), .out(tmp03_4_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010388(.in0(tmp02_10_81), .in1(tmp02_11_81), .out(tmp03_5_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010389(.in0(tmp02_12_81), .in1(tmp02_13_81), .out(tmp03_6_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010390(.in0(tmp02_14_81), .in1(tmp02_15_81), .out(tmp03_7_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010391(.in0(tmp02_16_81), .in1(tmp02_17_81), .out(tmp03_8_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010392(.in0(tmp02_18_81), .in1(tmp02_19_81), .out(tmp03_9_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010393(.in0(tmp02_20_81), .in1(tmp02_21_81), .out(tmp03_10_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010394(.in0(tmp02_22_81), .in1(tmp02_23_81), .out(tmp03_11_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010395(.in0(tmp02_24_81), .in1(tmp02_25_81), .out(tmp03_12_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010396(.in0(tmp02_26_81), .in1(tmp02_27_81), .out(tmp03_13_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010397(.in0(tmp02_28_81), .in1(tmp02_29_81), .out(tmp03_14_81));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010398(.in0(tmp02_30_81), .in1(tmp02_31_81), .out(tmp03_15_81));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010399(.in0(tmp03_0_81), .in1(tmp03_1_81), .out(tmp04_0_81));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010400(.in0(tmp03_2_81), .in1(tmp03_3_81), .out(tmp04_1_81));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010401(.in0(tmp03_4_81), .in1(tmp03_5_81), .out(tmp04_2_81));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010402(.in0(tmp03_6_81), .in1(tmp03_7_81), .out(tmp04_3_81));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010403(.in0(tmp03_8_81), .in1(tmp03_9_81), .out(tmp04_4_81));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010404(.in0(tmp03_10_81), .in1(tmp03_11_81), .out(tmp04_5_81));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010405(.in0(tmp03_12_81), .in1(tmp03_13_81), .out(tmp04_6_81));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010406(.in0(tmp03_14_81), .in1(tmp03_15_81), .out(tmp04_7_81));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010407(.in0(tmp04_0_81), .in1(tmp04_1_81), .out(tmp05_0_81));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010408(.in0(tmp04_2_81), .in1(tmp04_3_81), .out(tmp05_1_81));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010409(.in0(tmp04_4_81), .in1(tmp04_5_81), .out(tmp05_2_81));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010410(.in0(tmp04_6_81), .in1(tmp04_7_81), .out(tmp05_3_81));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010411(.in0(tmp05_0_81), .in1(tmp05_1_81), .out(tmp06_0_81));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010412(.in0(tmp05_2_81), .in1(tmp05_3_81), .out(tmp06_1_81));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add010413(.in0(tmp06_0_81), .in1(tmp06_1_81), .out(tmp07_0_81));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010414(.in0(tmp00_0_82), .in1(tmp00_1_82), .out(tmp01_0_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010415(.in0(tmp00_2_82), .in1(tmp00_3_82), .out(tmp01_1_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010416(.in0(tmp00_4_82), .in1(tmp00_5_82), .out(tmp01_2_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010417(.in0(tmp00_6_82), .in1(tmp00_7_82), .out(tmp01_3_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010418(.in0(tmp00_8_82), .in1(tmp00_9_82), .out(tmp01_4_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010419(.in0(tmp00_10_82), .in1(tmp00_11_82), .out(tmp01_5_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010420(.in0(tmp00_12_82), .in1(tmp00_13_82), .out(tmp01_6_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010421(.in0(tmp00_14_82), .in1(tmp00_15_82), .out(tmp01_7_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010422(.in0(tmp00_16_82), .in1(tmp00_17_82), .out(tmp01_8_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010423(.in0(tmp00_18_82), .in1(tmp00_19_82), .out(tmp01_9_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010424(.in0(tmp00_20_82), .in1(tmp00_21_82), .out(tmp01_10_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010425(.in0(tmp00_22_82), .in1(tmp00_23_82), .out(tmp01_11_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010426(.in0(tmp00_24_82), .in1(tmp00_25_82), .out(tmp01_12_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010427(.in0(tmp00_26_82), .in1(tmp00_27_82), .out(tmp01_13_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010428(.in0(tmp00_28_82), .in1(tmp00_29_82), .out(tmp01_14_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010429(.in0(tmp00_30_82), .in1(tmp00_31_82), .out(tmp01_15_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010430(.in0(tmp00_32_82), .in1(tmp00_33_82), .out(tmp01_16_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010431(.in0(tmp00_34_82), .in1(tmp00_35_82), .out(tmp01_17_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010432(.in0(tmp00_36_82), .in1(tmp00_37_82), .out(tmp01_18_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010433(.in0(tmp00_38_82), .in1(tmp00_39_82), .out(tmp01_19_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010434(.in0(tmp00_40_82), .in1(tmp00_41_82), .out(tmp01_20_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010435(.in0(tmp00_42_82), .in1(tmp00_43_82), .out(tmp01_21_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010436(.in0(tmp00_44_82), .in1(tmp00_45_82), .out(tmp01_22_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010437(.in0(tmp00_46_82), .in1(tmp00_47_82), .out(tmp01_23_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010438(.in0(tmp00_48_82), .in1(tmp00_49_82), .out(tmp01_24_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010439(.in0(tmp00_50_82), .in1(tmp00_51_82), .out(tmp01_25_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010440(.in0(tmp00_52_82), .in1(tmp00_53_82), .out(tmp01_26_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010441(.in0(tmp00_54_82), .in1(tmp00_55_82), .out(tmp01_27_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010442(.in0(tmp00_56_82), .in1(tmp00_57_82), .out(tmp01_28_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010443(.in0(tmp00_58_82), .in1(tmp00_59_82), .out(tmp01_29_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010444(.in0(tmp00_60_82), .in1(tmp00_61_82), .out(tmp01_30_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010445(.in0(tmp00_62_82), .in1(tmp00_63_82), .out(tmp01_31_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010446(.in0(tmp00_64_82), .in1(tmp00_65_82), .out(tmp01_32_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010447(.in0(tmp00_66_82), .in1(tmp00_67_82), .out(tmp01_33_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010448(.in0(tmp00_68_82), .in1(tmp00_69_82), .out(tmp01_34_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010449(.in0(tmp00_70_82), .in1(tmp00_71_82), .out(tmp01_35_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010450(.in0(tmp00_72_82), .in1(tmp00_73_82), .out(tmp01_36_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010451(.in0(tmp00_74_82), .in1(tmp00_75_82), .out(tmp01_37_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010452(.in0(tmp00_76_82), .in1(tmp00_77_82), .out(tmp01_38_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010453(.in0(tmp00_78_82), .in1(tmp00_79_82), .out(tmp01_39_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010454(.in0(tmp00_80_82), .in1(tmp00_81_82), .out(tmp01_40_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010455(.in0(tmp00_82_82), .in1(tmp00_83_82), .out(tmp01_41_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010456(.in0(tmp00_84_82), .in1(tmp00_85_82), .out(tmp01_42_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010457(.in0(tmp00_86_82), .in1(tmp00_87_82), .out(tmp01_43_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010458(.in0(tmp00_88_82), .in1(tmp00_89_82), .out(tmp01_44_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010459(.in0(tmp00_90_82), .in1(tmp00_91_82), .out(tmp01_45_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010460(.in0(tmp00_92_82), .in1(tmp00_93_82), .out(tmp01_46_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010461(.in0(tmp00_94_82), .in1(tmp00_95_82), .out(tmp01_47_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010462(.in0(tmp00_96_82), .in1(tmp00_97_82), .out(tmp01_48_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010463(.in0(tmp00_98_82), .in1(tmp00_99_82), .out(tmp01_49_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010464(.in0(tmp00_100_82), .in1(tmp00_101_82), .out(tmp01_50_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010465(.in0(tmp00_102_82), .in1(tmp00_103_82), .out(tmp01_51_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010466(.in0(tmp00_104_82), .in1(tmp00_105_82), .out(tmp01_52_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010467(.in0(tmp00_106_82), .in1(tmp00_107_82), .out(tmp01_53_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010468(.in0(tmp00_108_82), .in1(tmp00_109_82), .out(tmp01_54_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010469(.in0(tmp00_110_82), .in1(tmp00_111_82), .out(tmp01_55_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010470(.in0(tmp00_112_82), .in1(tmp00_113_82), .out(tmp01_56_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010471(.in0(tmp00_114_82), .in1(tmp00_115_82), .out(tmp01_57_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010472(.in0(tmp00_116_82), .in1(tmp00_117_82), .out(tmp01_58_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010473(.in0(tmp00_118_82), .in1(tmp00_119_82), .out(tmp01_59_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010474(.in0(tmp00_120_82), .in1(tmp00_121_82), .out(tmp01_60_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010475(.in0(tmp00_122_82), .in1(tmp00_123_82), .out(tmp01_61_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010476(.in0(tmp00_124_82), .in1(tmp00_125_82), .out(tmp01_62_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010477(.in0(tmp00_126_82), .in1(tmp00_127_82), .out(tmp01_63_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010478(.in0(tmp01_0_82), .in1(tmp01_1_82), .out(tmp02_0_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010479(.in0(tmp01_2_82), .in1(tmp01_3_82), .out(tmp02_1_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010480(.in0(tmp01_4_82), .in1(tmp01_5_82), .out(tmp02_2_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010481(.in0(tmp01_6_82), .in1(tmp01_7_82), .out(tmp02_3_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010482(.in0(tmp01_8_82), .in1(tmp01_9_82), .out(tmp02_4_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010483(.in0(tmp01_10_82), .in1(tmp01_11_82), .out(tmp02_5_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010484(.in0(tmp01_12_82), .in1(tmp01_13_82), .out(tmp02_6_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010485(.in0(tmp01_14_82), .in1(tmp01_15_82), .out(tmp02_7_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010486(.in0(tmp01_16_82), .in1(tmp01_17_82), .out(tmp02_8_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010487(.in0(tmp01_18_82), .in1(tmp01_19_82), .out(tmp02_9_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010488(.in0(tmp01_20_82), .in1(tmp01_21_82), .out(tmp02_10_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010489(.in0(tmp01_22_82), .in1(tmp01_23_82), .out(tmp02_11_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010490(.in0(tmp01_24_82), .in1(tmp01_25_82), .out(tmp02_12_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010491(.in0(tmp01_26_82), .in1(tmp01_27_82), .out(tmp02_13_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010492(.in0(tmp01_28_82), .in1(tmp01_29_82), .out(tmp02_14_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010493(.in0(tmp01_30_82), .in1(tmp01_31_82), .out(tmp02_15_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010494(.in0(tmp01_32_82), .in1(tmp01_33_82), .out(tmp02_16_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010495(.in0(tmp01_34_82), .in1(tmp01_35_82), .out(tmp02_17_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010496(.in0(tmp01_36_82), .in1(tmp01_37_82), .out(tmp02_18_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010497(.in0(tmp01_38_82), .in1(tmp01_39_82), .out(tmp02_19_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010498(.in0(tmp01_40_82), .in1(tmp01_41_82), .out(tmp02_20_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010499(.in0(tmp01_42_82), .in1(tmp01_43_82), .out(tmp02_21_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010500(.in0(tmp01_44_82), .in1(tmp01_45_82), .out(tmp02_22_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010501(.in0(tmp01_46_82), .in1(tmp01_47_82), .out(tmp02_23_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010502(.in0(tmp01_48_82), .in1(tmp01_49_82), .out(tmp02_24_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010503(.in0(tmp01_50_82), .in1(tmp01_51_82), .out(tmp02_25_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010504(.in0(tmp01_52_82), .in1(tmp01_53_82), .out(tmp02_26_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010505(.in0(tmp01_54_82), .in1(tmp01_55_82), .out(tmp02_27_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010506(.in0(tmp01_56_82), .in1(tmp01_57_82), .out(tmp02_28_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010507(.in0(tmp01_58_82), .in1(tmp01_59_82), .out(tmp02_29_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010508(.in0(tmp01_60_82), .in1(tmp01_61_82), .out(tmp02_30_82));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010509(.in0(tmp01_62_82), .in1(tmp01_63_82), .out(tmp02_31_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010510(.in0(tmp02_0_82), .in1(tmp02_1_82), .out(tmp03_0_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010511(.in0(tmp02_2_82), .in1(tmp02_3_82), .out(tmp03_1_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010512(.in0(tmp02_4_82), .in1(tmp02_5_82), .out(tmp03_2_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010513(.in0(tmp02_6_82), .in1(tmp02_7_82), .out(tmp03_3_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010514(.in0(tmp02_8_82), .in1(tmp02_9_82), .out(tmp03_4_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010515(.in0(tmp02_10_82), .in1(tmp02_11_82), .out(tmp03_5_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010516(.in0(tmp02_12_82), .in1(tmp02_13_82), .out(tmp03_6_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010517(.in0(tmp02_14_82), .in1(tmp02_15_82), .out(tmp03_7_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010518(.in0(tmp02_16_82), .in1(tmp02_17_82), .out(tmp03_8_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010519(.in0(tmp02_18_82), .in1(tmp02_19_82), .out(tmp03_9_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010520(.in0(tmp02_20_82), .in1(tmp02_21_82), .out(tmp03_10_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010521(.in0(tmp02_22_82), .in1(tmp02_23_82), .out(tmp03_11_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010522(.in0(tmp02_24_82), .in1(tmp02_25_82), .out(tmp03_12_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010523(.in0(tmp02_26_82), .in1(tmp02_27_82), .out(tmp03_13_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010524(.in0(tmp02_28_82), .in1(tmp02_29_82), .out(tmp03_14_82));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010525(.in0(tmp02_30_82), .in1(tmp02_31_82), .out(tmp03_15_82));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010526(.in0(tmp03_0_82), .in1(tmp03_1_82), .out(tmp04_0_82));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010527(.in0(tmp03_2_82), .in1(tmp03_3_82), .out(tmp04_1_82));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010528(.in0(tmp03_4_82), .in1(tmp03_5_82), .out(tmp04_2_82));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010529(.in0(tmp03_6_82), .in1(tmp03_7_82), .out(tmp04_3_82));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010530(.in0(tmp03_8_82), .in1(tmp03_9_82), .out(tmp04_4_82));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010531(.in0(tmp03_10_82), .in1(tmp03_11_82), .out(tmp04_5_82));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010532(.in0(tmp03_12_82), .in1(tmp03_13_82), .out(tmp04_6_82));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010533(.in0(tmp03_14_82), .in1(tmp03_15_82), .out(tmp04_7_82));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010534(.in0(tmp04_0_82), .in1(tmp04_1_82), .out(tmp05_0_82));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010535(.in0(tmp04_2_82), .in1(tmp04_3_82), .out(tmp05_1_82));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010536(.in0(tmp04_4_82), .in1(tmp04_5_82), .out(tmp05_2_82));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010537(.in0(tmp04_6_82), .in1(tmp04_7_82), .out(tmp05_3_82));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010538(.in0(tmp05_0_82), .in1(tmp05_1_82), .out(tmp06_0_82));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010539(.in0(tmp05_2_82), .in1(tmp05_3_82), .out(tmp06_1_82));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add010540(.in0(tmp06_0_82), .in1(tmp06_1_82), .out(tmp07_0_82));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010541(.in0(tmp00_0_83), .in1(tmp00_1_83), .out(tmp01_0_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010542(.in0(tmp00_2_83), .in1(tmp00_3_83), .out(tmp01_1_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010543(.in0(tmp00_4_83), .in1(tmp00_5_83), .out(tmp01_2_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010544(.in0(tmp00_6_83), .in1(tmp00_7_83), .out(tmp01_3_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010545(.in0(tmp00_8_83), .in1(tmp00_9_83), .out(tmp01_4_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010546(.in0(tmp00_10_83), .in1(tmp00_11_83), .out(tmp01_5_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010547(.in0(tmp00_12_83), .in1(tmp00_13_83), .out(tmp01_6_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010548(.in0(tmp00_14_83), .in1(tmp00_15_83), .out(tmp01_7_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010549(.in0(tmp00_16_83), .in1(tmp00_17_83), .out(tmp01_8_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010550(.in0(tmp00_18_83), .in1(tmp00_19_83), .out(tmp01_9_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010551(.in0(tmp00_20_83), .in1(tmp00_21_83), .out(tmp01_10_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010552(.in0(tmp00_22_83), .in1(tmp00_23_83), .out(tmp01_11_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010553(.in0(tmp00_24_83), .in1(tmp00_25_83), .out(tmp01_12_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010554(.in0(tmp00_26_83), .in1(tmp00_27_83), .out(tmp01_13_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010555(.in0(tmp00_28_83), .in1(tmp00_29_83), .out(tmp01_14_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010556(.in0(tmp00_30_83), .in1(tmp00_31_83), .out(tmp01_15_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010557(.in0(tmp00_32_83), .in1(tmp00_33_83), .out(tmp01_16_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010558(.in0(tmp00_34_83), .in1(tmp00_35_83), .out(tmp01_17_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010559(.in0(tmp00_36_83), .in1(tmp00_37_83), .out(tmp01_18_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010560(.in0(tmp00_38_83), .in1(tmp00_39_83), .out(tmp01_19_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010561(.in0(tmp00_40_83), .in1(tmp00_41_83), .out(tmp01_20_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010562(.in0(tmp00_42_83), .in1(tmp00_43_83), .out(tmp01_21_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010563(.in0(tmp00_44_83), .in1(tmp00_45_83), .out(tmp01_22_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010564(.in0(tmp00_46_83), .in1(tmp00_47_83), .out(tmp01_23_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010565(.in0(tmp00_48_83), .in1(tmp00_49_83), .out(tmp01_24_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010566(.in0(tmp00_50_83), .in1(tmp00_51_83), .out(tmp01_25_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010567(.in0(tmp00_52_83), .in1(tmp00_53_83), .out(tmp01_26_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010568(.in0(tmp00_54_83), .in1(tmp00_55_83), .out(tmp01_27_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010569(.in0(tmp00_56_83), .in1(tmp00_57_83), .out(tmp01_28_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010570(.in0(tmp00_58_83), .in1(tmp00_59_83), .out(tmp01_29_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010571(.in0(tmp00_60_83), .in1(tmp00_61_83), .out(tmp01_30_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010572(.in0(tmp00_62_83), .in1(tmp00_63_83), .out(tmp01_31_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010573(.in0(tmp00_64_83), .in1(tmp00_65_83), .out(tmp01_32_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010574(.in0(tmp00_66_83), .in1(tmp00_67_83), .out(tmp01_33_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010575(.in0(tmp00_68_83), .in1(tmp00_69_83), .out(tmp01_34_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010576(.in0(tmp00_70_83), .in1(tmp00_71_83), .out(tmp01_35_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010577(.in0(tmp00_72_83), .in1(tmp00_73_83), .out(tmp01_36_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010578(.in0(tmp00_74_83), .in1(tmp00_75_83), .out(tmp01_37_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010579(.in0(tmp00_76_83), .in1(tmp00_77_83), .out(tmp01_38_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010580(.in0(tmp00_78_83), .in1(tmp00_79_83), .out(tmp01_39_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010581(.in0(tmp00_80_83), .in1(tmp00_81_83), .out(tmp01_40_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010582(.in0(tmp00_82_83), .in1(tmp00_83_83), .out(tmp01_41_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010583(.in0(tmp00_84_83), .in1(tmp00_85_83), .out(tmp01_42_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010584(.in0(tmp00_86_83), .in1(tmp00_87_83), .out(tmp01_43_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010585(.in0(tmp00_88_83), .in1(tmp00_89_83), .out(tmp01_44_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010586(.in0(tmp00_90_83), .in1(tmp00_91_83), .out(tmp01_45_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010587(.in0(tmp00_92_83), .in1(tmp00_93_83), .out(tmp01_46_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010588(.in0(tmp00_94_83), .in1(tmp00_95_83), .out(tmp01_47_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010589(.in0(tmp00_96_83), .in1(tmp00_97_83), .out(tmp01_48_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010590(.in0(tmp00_98_83), .in1(tmp00_99_83), .out(tmp01_49_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010591(.in0(tmp00_100_83), .in1(tmp00_101_83), .out(tmp01_50_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010592(.in0(tmp00_102_83), .in1(tmp00_103_83), .out(tmp01_51_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010593(.in0(tmp00_104_83), .in1(tmp00_105_83), .out(tmp01_52_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010594(.in0(tmp00_106_83), .in1(tmp00_107_83), .out(tmp01_53_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010595(.in0(tmp00_108_83), .in1(tmp00_109_83), .out(tmp01_54_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010596(.in0(tmp00_110_83), .in1(tmp00_111_83), .out(tmp01_55_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010597(.in0(tmp00_112_83), .in1(tmp00_113_83), .out(tmp01_56_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010598(.in0(tmp00_114_83), .in1(tmp00_115_83), .out(tmp01_57_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010599(.in0(tmp00_116_83), .in1(tmp00_117_83), .out(tmp01_58_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010600(.in0(tmp00_118_83), .in1(tmp00_119_83), .out(tmp01_59_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010601(.in0(tmp00_120_83), .in1(tmp00_121_83), .out(tmp01_60_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010602(.in0(tmp00_122_83), .in1(tmp00_123_83), .out(tmp01_61_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010603(.in0(tmp00_124_83), .in1(tmp00_125_83), .out(tmp01_62_83));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add010604(.in0(tmp00_126_83), .in1(tmp00_127_83), .out(tmp01_63_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010605(.in0(tmp01_0_83), .in1(tmp01_1_83), .out(tmp02_0_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010606(.in0(tmp01_2_83), .in1(tmp01_3_83), .out(tmp02_1_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010607(.in0(tmp01_4_83), .in1(tmp01_5_83), .out(tmp02_2_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010608(.in0(tmp01_6_83), .in1(tmp01_7_83), .out(tmp02_3_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010609(.in0(tmp01_8_83), .in1(tmp01_9_83), .out(tmp02_4_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010610(.in0(tmp01_10_83), .in1(tmp01_11_83), .out(tmp02_5_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010611(.in0(tmp01_12_83), .in1(tmp01_13_83), .out(tmp02_6_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010612(.in0(tmp01_14_83), .in1(tmp01_15_83), .out(tmp02_7_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010613(.in0(tmp01_16_83), .in1(tmp01_17_83), .out(tmp02_8_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010614(.in0(tmp01_18_83), .in1(tmp01_19_83), .out(tmp02_9_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010615(.in0(tmp01_20_83), .in1(tmp01_21_83), .out(tmp02_10_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010616(.in0(tmp01_22_83), .in1(tmp01_23_83), .out(tmp02_11_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010617(.in0(tmp01_24_83), .in1(tmp01_25_83), .out(tmp02_12_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010618(.in0(tmp01_26_83), .in1(tmp01_27_83), .out(tmp02_13_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010619(.in0(tmp01_28_83), .in1(tmp01_29_83), .out(tmp02_14_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010620(.in0(tmp01_30_83), .in1(tmp01_31_83), .out(tmp02_15_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010621(.in0(tmp01_32_83), .in1(tmp01_33_83), .out(tmp02_16_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010622(.in0(tmp01_34_83), .in1(tmp01_35_83), .out(tmp02_17_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010623(.in0(tmp01_36_83), .in1(tmp01_37_83), .out(tmp02_18_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010624(.in0(tmp01_38_83), .in1(tmp01_39_83), .out(tmp02_19_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010625(.in0(tmp01_40_83), .in1(tmp01_41_83), .out(tmp02_20_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010626(.in0(tmp01_42_83), .in1(tmp01_43_83), .out(tmp02_21_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010627(.in0(tmp01_44_83), .in1(tmp01_45_83), .out(tmp02_22_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010628(.in0(tmp01_46_83), .in1(tmp01_47_83), .out(tmp02_23_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010629(.in0(tmp01_48_83), .in1(tmp01_49_83), .out(tmp02_24_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010630(.in0(tmp01_50_83), .in1(tmp01_51_83), .out(tmp02_25_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010631(.in0(tmp01_52_83), .in1(tmp01_53_83), .out(tmp02_26_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010632(.in0(tmp01_54_83), .in1(tmp01_55_83), .out(tmp02_27_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010633(.in0(tmp01_56_83), .in1(tmp01_57_83), .out(tmp02_28_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010634(.in0(tmp01_58_83), .in1(tmp01_59_83), .out(tmp02_29_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010635(.in0(tmp01_60_83), .in1(tmp01_61_83), .out(tmp02_30_83));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add010636(.in0(tmp01_62_83), .in1(tmp01_63_83), .out(tmp02_31_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010637(.in0(tmp02_0_83), .in1(tmp02_1_83), .out(tmp03_0_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010638(.in0(tmp02_2_83), .in1(tmp02_3_83), .out(tmp03_1_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010639(.in0(tmp02_4_83), .in1(tmp02_5_83), .out(tmp03_2_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010640(.in0(tmp02_6_83), .in1(tmp02_7_83), .out(tmp03_3_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010641(.in0(tmp02_8_83), .in1(tmp02_9_83), .out(tmp03_4_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010642(.in0(tmp02_10_83), .in1(tmp02_11_83), .out(tmp03_5_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010643(.in0(tmp02_12_83), .in1(tmp02_13_83), .out(tmp03_6_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010644(.in0(tmp02_14_83), .in1(tmp02_15_83), .out(tmp03_7_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010645(.in0(tmp02_16_83), .in1(tmp02_17_83), .out(tmp03_8_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010646(.in0(tmp02_18_83), .in1(tmp02_19_83), .out(tmp03_9_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010647(.in0(tmp02_20_83), .in1(tmp02_21_83), .out(tmp03_10_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010648(.in0(tmp02_22_83), .in1(tmp02_23_83), .out(tmp03_11_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010649(.in0(tmp02_24_83), .in1(tmp02_25_83), .out(tmp03_12_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010650(.in0(tmp02_26_83), .in1(tmp02_27_83), .out(tmp03_13_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010651(.in0(tmp02_28_83), .in1(tmp02_29_83), .out(tmp03_14_83));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add010652(.in0(tmp02_30_83), .in1(tmp02_31_83), .out(tmp03_15_83));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010653(.in0(tmp03_0_83), .in1(tmp03_1_83), .out(tmp04_0_83));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010654(.in0(tmp03_2_83), .in1(tmp03_3_83), .out(tmp04_1_83));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010655(.in0(tmp03_4_83), .in1(tmp03_5_83), .out(tmp04_2_83));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010656(.in0(tmp03_6_83), .in1(tmp03_7_83), .out(tmp04_3_83));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010657(.in0(tmp03_8_83), .in1(tmp03_9_83), .out(tmp04_4_83));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010658(.in0(tmp03_10_83), .in1(tmp03_11_83), .out(tmp04_5_83));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010659(.in0(tmp03_12_83), .in1(tmp03_13_83), .out(tmp04_6_83));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add010660(.in0(tmp03_14_83), .in1(tmp03_15_83), .out(tmp04_7_83));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010661(.in0(tmp04_0_83), .in1(tmp04_1_83), .out(tmp05_0_83));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010662(.in0(tmp04_2_83), .in1(tmp04_3_83), .out(tmp05_1_83));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010663(.in0(tmp04_4_83), .in1(tmp04_5_83), .out(tmp05_2_83));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add010664(.in0(tmp04_6_83), .in1(tmp04_7_83), .out(tmp05_3_83));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010665(.in0(tmp05_0_83), .in1(tmp05_1_83), .out(tmp06_0_83));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add010666(.in0(tmp05_2_83), .in1(tmp05_3_83), .out(tmp06_1_83));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add010667(.in0(tmp06_0_83), .in1(tmp06_1_83), .out(tmp07_0_83));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU000(.a(tmp07_0_0), .b(23'h0), .sel(tmp07_0_0[WIDTH*2+$clog2(IN)-1]), .out(z_0));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU001(.a(tmp07_0_1), .b(23'h0), .sel(tmp07_0_1[WIDTH*2+$clog2(IN)-1]), .out(z_1));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU002(.a(tmp07_0_2), .b(23'h0), .sel(tmp07_0_2[WIDTH*2+$clog2(IN)-1]), .out(z_2));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU003(.a(tmp07_0_3), .b(23'h0), .sel(tmp07_0_3[WIDTH*2+$clog2(IN)-1]), .out(z_3));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU004(.a(tmp07_0_4), .b(23'h0), .sel(tmp07_0_4[WIDTH*2+$clog2(IN)-1]), .out(z_4));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU005(.a(tmp07_0_5), .b(23'h0), .sel(tmp07_0_5[WIDTH*2+$clog2(IN)-1]), .out(z_5));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU006(.a(tmp07_0_6), .b(23'h0), .sel(tmp07_0_6[WIDTH*2+$clog2(IN)-1]), .out(z_6));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU007(.a(tmp07_0_7), .b(23'h0), .sel(tmp07_0_7[WIDTH*2+$clog2(IN)-1]), .out(z_7));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU008(.a(tmp07_0_8), .b(23'h0), .sel(tmp07_0_8[WIDTH*2+$clog2(IN)-1]), .out(z_8));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU009(.a(tmp07_0_9), .b(23'h0), .sel(tmp07_0_9[WIDTH*2+$clog2(IN)-1]), .out(z_9));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU010(.a(tmp07_0_10), .b(23'h0), .sel(tmp07_0_10[WIDTH*2+$clog2(IN)-1]), .out(z_10));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU011(.a(tmp07_0_11), .b(23'h0), .sel(tmp07_0_11[WIDTH*2+$clog2(IN)-1]), .out(z_11));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU012(.a(tmp07_0_12), .b(23'h0), .sel(tmp07_0_12[WIDTH*2+$clog2(IN)-1]), .out(z_12));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU013(.a(tmp07_0_13), .b(23'h0), .sel(tmp07_0_13[WIDTH*2+$clog2(IN)-1]), .out(z_13));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU014(.a(tmp07_0_14), .b(23'h0), .sel(tmp07_0_14[WIDTH*2+$clog2(IN)-1]), .out(z_14));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU015(.a(tmp07_0_15), .b(23'h0), .sel(tmp07_0_15[WIDTH*2+$clog2(IN)-1]), .out(z_15));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU016(.a(tmp07_0_16), .b(23'h0), .sel(tmp07_0_16[WIDTH*2+$clog2(IN)-1]), .out(z_16));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU017(.a(tmp07_0_17), .b(23'h0), .sel(tmp07_0_17[WIDTH*2+$clog2(IN)-1]), .out(z_17));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU018(.a(tmp07_0_18), .b(23'h0), .sel(tmp07_0_18[WIDTH*2+$clog2(IN)-1]), .out(z_18));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU019(.a(tmp07_0_19), .b(23'h0), .sel(tmp07_0_19[WIDTH*2+$clog2(IN)-1]), .out(z_19));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU020(.a(tmp07_0_20), .b(23'h0), .sel(tmp07_0_20[WIDTH*2+$clog2(IN)-1]), .out(z_20));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU021(.a(tmp07_0_21), .b(23'h0), .sel(tmp07_0_21[WIDTH*2+$clog2(IN)-1]), .out(z_21));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU022(.a(tmp07_0_22), .b(23'h0), .sel(tmp07_0_22[WIDTH*2+$clog2(IN)-1]), .out(z_22));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU023(.a(tmp07_0_23), .b(23'h0), .sel(tmp07_0_23[WIDTH*2+$clog2(IN)-1]), .out(z_23));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU024(.a(tmp07_0_24), .b(23'h0), .sel(tmp07_0_24[WIDTH*2+$clog2(IN)-1]), .out(z_24));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU025(.a(tmp07_0_25), .b(23'h0), .sel(tmp07_0_25[WIDTH*2+$clog2(IN)-1]), .out(z_25));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU026(.a(tmp07_0_26), .b(23'h0), .sel(tmp07_0_26[WIDTH*2+$clog2(IN)-1]), .out(z_26));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU027(.a(tmp07_0_27), .b(23'h0), .sel(tmp07_0_27[WIDTH*2+$clog2(IN)-1]), .out(z_27));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU028(.a(tmp07_0_28), .b(23'h0), .sel(tmp07_0_28[WIDTH*2+$clog2(IN)-1]), .out(z_28));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU029(.a(tmp07_0_29), .b(23'h0), .sel(tmp07_0_29[WIDTH*2+$clog2(IN)-1]), .out(z_29));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU030(.a(tmp07_0_30), .b(23'h0), .sel(tmp07_0_30[WIDTH*2+$clog2(IN)-1]), .out(z_30));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU031(.a(tmp07_0_31), .b(23'h0), .sel(tmp07_0_31[WIDTH*2+$clog2(IN)-1]), .out(z_31));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU032(.a(tmp07_0_32), .b(23'h0), .sel(tmp07_0_32[WIDTH*2+$clog2(IN)-1]), .out(z_32));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU033(.a(tmp07_0_33), .b(23'h0), .sel(tmp07_0_33[WIDTH*2+$clog2(IN)-1]), .out(z_33));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU034(.a(tmp07_0_34), .b(23'h0), .sel(tmp07_0_34[WIDTH*2+$clog2(IN)-1]), .out(z_34));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU035(.a(tmp07_0_35), .b(23'h0), .sel(tmp07_0_35[WIDTH*2+$clog2(IN)-1]), .out(z_35));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU036(.a(tmp07_0_36), .b(23'h0), .sel(tmp07_0_36[WIDTH*2+$clog2(IN)-1]), .out(z_36));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU037(.a(tmp07_0_37), .b(23'h0), .sel(tmp07_0_37[WIDTH*2+$clog2(IN)-1]), .out(z_37));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU038(.a(tmp07_0_38), .b(23'h0), .sel(tmp07_0_38[WIDTH*2+$clog2(IN)-1]), .out(z_38));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU039(.a(tmp07_0_39), .b(23'h0), .sel(tmp07_0_39[WIDTH*2+$clog2(IN)-1]), .out(z_39));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU040(.a(tmp07_0_40), .b(23'h0), .sel(tmp07_0_40[WIDTH*2+$clog2(IN)-1]), .out(z_40));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU041(.a(tmp07_0_41), .b(23'h0), .sel(tmp07_0_41[WIDTH*2+$clog2(IN)-1]), .out(z_41));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU042(.a(tmp07_0_42), .b(23'h0), .sel(tmp07_0_42[WIDTH*2+$clog2(IN)-1]), .out(z_42));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU043(.a(tmp07_0_43), .b(23'h0), .sel(tmp07_0_43[WIDTH*2+$clog2(IN)-1]), .out(z_43));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU044(.a(tmp07_0_44), .b(23'h0), .sel(tmp07_0_44[WIDTH*2+$clog2(IN)-1]), .out(z_44));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU045(.a(tmp07_0_45), .b(23'h0), .sel(tmp07_0_45[WIDTH*2+$clog2(IN)-1]), .out(z_45));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU046(.a(tmp07_0_46), .b(23'h0), .sel(tmp07_0_46[WIDTH*2+$clog2(IN)-1]), .out(z_46));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU047(.a(tmp07_0_47), .b(23'h0), .sel(tmp07_0_47[WIDTH*2+$clog2(IN)-1]), .out(z_47));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU048(.a(tmp07_0_48), .b(23'h0), .sel(tmp07_0_48[WIDTH*2+$clog2(IN)-1]), .out(z_48));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU049(.a(tmp07_0_49), .b(23'h0), .sel(tmp07_0_49[WIDTH*2+$clog2(IN)-1]), .out(z_49));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU050(.a(tmp07_0_50), .b(23'h0), .sel(tmp07_0_50[WIDTH*2+$clog2(IN)-1]), .out(z_50));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU051(.a(tmp07_0_51), .b(23'h0), .sel(tmp07_0_51[WIDTH*2+$clog2(IN)-1]), .out(z_51));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU052(.a(tmp07_0_52), .b(23'h0), .sel(tmp07_0_52[WIDTH*2+$clog2(IN)-1]), .out(z_52));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU053(.a(tmp07_0_53), .b(23'h0), .sel(tmp07_0_53[WIDTH*2+$clog2(IN)-1]), .out(z_53));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU054(.a(tmp07_0_54), .b(23'h0), .sel(tmp07_0_54[WIDTH*2+$clog2(IN)-1]), .out(z_54));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU055(.a(tmp07_0_55), .b(23'h0), .sel(tmp07_0_55[WIDTH*2+$clog2(IN)-1]), .out(z_55));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU056(.a(tmp07_0_56), .b(23'h0), .sel(tmp07_0_56[WIDTH*2+$clog2(IN)-1]), .out(z_56));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU057(.a(tmp07_0_57), .b(23'h0), .sel(tmp07_0_57[WIDTH*2+$clog2(IN)-1]), .out(z_57));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU058(.a(tmp07_0_58), .b(23'h0), .sel(tmp07_0_58[WIDTH*2+$clog2(IN)-1]), .out(z_58));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU059(.a(tmp07_0_59), .b(23'h0), .sel(tmp07_0_59[WIDTH*2+$clog2(IN)-1]), .out(z_59));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU060(.a(tmp07_0_60), .b(23'h0), .sel(tmp07_0_60[WIDTH*2+$clog2(IN)-1]), .out(z_60));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU061(.a(tmp07_0_61), .b(23'h0), .sel(tmp07_0_61[WIDTH*2+$clog2(IN)-1]), .out(z_61));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU062(.a(tmp07_0_62), .b(23'h0), .sel(tmp07_0_62[WIDTH*2+$clog2(IN)-1]), .out(z_62));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU063(.a(tmp07_0_63), .b(23'h0), .sel(tmp07_0_63[WIDTH*2+$clog2(IN)-1]), .out(z_63));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU064(.a(tmp07_0_64), .b(23'h0), .sel(tmp07_0_64[WIDTH*2+$clog2(IN)-1]), .out(z_64));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU065(.a(tmp07_0_65), .b(23'h0), .sel(tmp07_0_65[WIDTH*2+$clog2(IN)-1]), .out(z_65));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU066(.a(tmp07_0_66), .b(23'h0), .sel(tmp07_0_66[WIDTH*2+$clog2(IN)-1]), .out(z_66));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU067(.a(tmp07_0_67), .b(23'h0), .sel(tmp07_0_67[WIDTH*2+$clog2(IN)-1]), .out(z_67));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU068(.a(tmp07_0_68), .b(23'h0), .sel(tmp07_0_68[WIDTH*2+$clog2(IN)-1]), .out(z_68));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU069(.a(tmp07_0_69), .b(23'h0), .sel(tmp07_0_69[WIDTH*2+$clog2(IN)-1]), .out(z_69));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU070(.a(tmp07_0_70), .b(23'h0), .sel(tmp07_0_70[WIDTH*2+$clog2(IN)-1]), .out(z_70));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU071(.a(tmp07_0_71), .b(23'h0), .sel(tmp07_0_71[WIDTH*2+$clog2(IN)-1]), .out(z_71));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU072(.a(tmp07_0_72), .b(23'h0), .sel(tmp07_0_72[WIDTH*2+$clog2(IN)-1]), .out(z_72));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU073(.a(tmp07_0_73), .b(23'h0), .sel(tmp07_0_73[WIDTH*2+$clog2(IN)-1]), .out(z_73));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU074(.a(tmp07_0_74), .b(23'h0), .sel(tmp07_0_74[WIDTH*2+$clog2(IN)-1]), .out(z_74));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU075(.a(tmp07_0_75), .b(23'h0), .sel(tmp07_0_75[WIDTH*2+$clog2(IN)-1]), .out(z_75));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU076(.a(tmp07_0_76), .b(23'h0), .sel(tmp07_0_76[WIDTH*2+$clog2(IN)-1]), .out(z_76));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU077(.a(tmp07_0_77), .b(23'h0), .sel(tmp07_0_77[WIDTH*2+$clog2(IN)-1]), .out(z_77));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU078(.a(tmp07_0_78), .b(23'h0), .sel(tmp07_0_78[WIDTH*2+$clog2(IN)-1]), .out(z_78));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU079(.a(tmp07_0_79), .b(23'h0), .sel(tmp07_0_79[WIDTH*2+$clog2(IN)-1]), .out(z_79));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU080(.a(tmp07_0_80), .b(23'h0), .sel(tmp07_0_80[WIDTH*2+$clog2(IN)-1]), .out(z_80));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU081(.a(tmp07_0_81), .b(23'h0), .sel(tmp07_0_81[WIDTH*2+$clog2(IN)-1]), .out(z_81));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU082(.a(tmp07_0_82), .b(23'h0), .sel(tmp07_0_82[WIDTH*2+$clog2(IN)-1]), .out(z_82));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU083(.a(tmp07_0_83), .b(23'h0), .sel(tmp07_0_83[WIDTH*2+$clog2(IN)-1]), .out(z_83));
endmodule

