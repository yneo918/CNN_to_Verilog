module tb;
	localparam WIDTH = 8;
	localparam IN = 256;
	localparam OUT = 128;
	logic [WIDTH-1:0] x[0:IN-1];
	logic [WIDTH*2+$clog2(IN)-1:0] z[0:OUT-1];
	logic [WIDTH*2+$clog2(IN)-1:0] exp[0:OUT-1];
	fc256_128 #(.WIDTH(WIDTH)) fc(.x(x), .z(z));
	initial begin
		$readmemh("exp",exp);
		x <= '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};

		#10
		x <= '{ 8'ha5, 8'h59, 8'h39, 8'h78, 8'hb2, 8'h71, 8'ha1, 8'hfc, 8'h15, 8'hd0, 8'hfc, 8'hb6, 8'he1, 8'h45, 8'hd2, 8'h7, 8'h5f, 8'haa, 8'h6b, 8'hd4, 8'ha7, 8'h31, 8'hd7, 8'h4c, 8'h4b, 8'h63, 8'h3d, 8'h28, 8'h32, 8'h13, 8'h4, 8'hd6, 8'hd, 8'h6f, 8'h27, 8'hf5, 8'h64, 8'hd8, 8'h57, 8'h23, 8'h6f, 8'h6, 8'h6f, 8'hfb, 8'h1f, 8'h52, 8'h38, 8'hc5, 8'hee, 8'h2b, 8'he9, 8'h96, 8'h1f, 8'h85, 8'h60, 8'h25, 8'h79, 8'h8, 8'h3e, 8'h7c, 8'h82, 8'h6e, 8'he2, 8'h6a, 8'h86, 8'hf1, 8'ha2, 8'h76, 8'h48, 8'h8a, 8'h4b, 8'h18, 8'hd, 8'h18, 8'h8c, 8'hfa, 8'h4f, 8'h7c, 8'h45, 8'h6f, 8'hdb, 8'h18, 8'h47, 8'he4, 8'h1f, 8'h91, 8'h6a, 8'hdf, 8'hd9, 8'h9c, 8'h56, 8'hd1, 8'hfa, 8'h99, 8'h98, 8'h2d, 8'h4, 8'h8, 8'h5d, 8'h53, 8'h25, 8'he1, 8'h5d, 8'h86, 8'h9f, 8'h52, 8'ha8, 8'hb8, 8'h49, 8'h99, 8'h54, 8'h9a, 8'h93, 8'h68, 8'h40, 8'h4f, 8'h34, 8'haa, 8'h6a, 8'h43, 8'h9d, 8'h87, 8'hd7, 8'h6f, 8'h1f, 8'h38, 8'h5f, 8'ha7, 8'ha5, 8'hab, 8'h7d, 8'h21, 8'h84, 8'h7f, 8'h58, 8'haf, 8'h3c, 8'ha3, 8'h92, 8'hb9, 8'h6d, 8'ha6, 8'h1a, 8'hf3, 8'h1a, 8'h51, 8'h89, 8'h4a, 8'h6c, 8'h72, 8'h41, 8'h60, 8'h66, 8'h55, 8'h92, 8'h39, 8'h8f, 8'h70, 8'h56, 8'h16, 8'h1d, 8'h1a, 8'hdf, 8'hfa, 8'h1d, 8'he4, 8'h55, 8'h2a, 8'he1, 8'h4e, 8'hfb, 8'h37, 8'h59, 8'hce, 8'hd8, 8'h8f, 8'h3b, 8'h8b, 8'h9b, 8'hf7, 8'h31, 8'h15, 8'h52, 8'h2f, 8'h2, 8'he2, 8'hcb, 8'h82, 8'h96, 8'h8, 8'h5a, 8'hfb, 8'hdf, 8'h80, 8'h16, 8'hc, 8'h45, 8'h5, 8'h7, 8'h94, 8'h5, 8'hb1, 8'h36, 8'h39, 8'h84, 8'h7c, 8'h11, 8'h34, 8'h4d, 8'hf, 8'h95, 8'h8b, 8'hd, 8'h54, 8'hb9, 8'h12, 8'h8e, 8'hbf, 8'h4d, 8'h1e, 8'h2a, 8'hc8, 8'hf5, 8'h1a, 8'h6c, 8'hdc, 8'hf6, 8'hb2, 8'hb0, 8'h67, 8'hb3, 8'ha0, 8'h1a, 8'h43, 8'hd5, 8'h21, 8'he3, 8'hf0, 8'h92, 8'h3c, 8'ha, 8'hb4, 8'h79, 8'h8d, 8'h82, 8'h4c, 8'hd6, 8'h21, 8'h4d, 8'h4d, 8'h8c, 8'h98, 8'he8, 8'h81, 8'h2a, 8'h9d };
		#10
		if (exp !== z)begin
			$display("Mismatch Error");
			$display("out: z0=0x%0h z1=0x%0h z2=0x%0h z3=0x%0h z4=0x%0h z5=0x%0h z6=0x%0h z7=0x%0h z8=0x%0h z9=0x%0h ",z[0], z[1], z[2], z[3], z[4], z[5], z[6], z[7], z[8], z[9]);
			$display("exp: z0=0x%0h z1=0x%0h z2=0x%0h z3=0x%0h z4=0x%0h z5=0x%0h z6=0x%0h z7=0x%0h z8=0x%0h z9=0x%0h ",exp[0], exp[1], exp[2], exp[3], exp[4], exp[5], exp[6], exp[7], exp[8], exp[9]);
		end
		if (exp == z)begin
			$display("\nPASS\n");
		end
		#10 $finish;

	end
endmodule
