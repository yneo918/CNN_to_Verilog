module fc84_10
	#(parameter WIDTH = 8)
	(x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7, x_8, x_9, x_10, x_11, x_12, x_13, x_14, x_15, x_16, x_17, x_18, x_19, x_20, x_21, x_22, x_23, x_24, x_25, x_26, x_27, x_28, x_29, x_30, x_31, x_32, x_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, z_0, z_1, z_2, z_3, z_4, z_5, z_6, z_7, z_8, z_9 );
	localparam IN = 84, OUT = 10;
	input [WIDTH-1:0] x_0;
	input [WIDTH-1:0] x_1;
	input [WIDTH-1:0] x_2;
	input [WIDTH-1:0] x_3;
	input [WIDTH-1:0] x_4;
	input [WIDTH-1:0] x_5;
	input [WIDTH-1:0] x_6;
	input [WIDTH-1:0] x_7;
	input [WIDTH-1:0] x_8;
	input [WIDTH-1:0] x_9;
	input [WIDTH-1:0] x_10;
	input [WIDTH-1:0] x_11;
	input [WIDTH-1:0] x_12;
	input [WIDTH-1:0] x_13;
	input [WIDTH-1:0] x_14;
	input [WIDTH-1:0] x_15;
	input [WIDTH-1:0] x_16;
	input [WIDTH-1:0] x_17;
	input [WIDTH-1:0] x_18;
	input [WIDTH-1:0] x_19;
	input [WIDTH-1:0] x_20;
	input [WIDTH-1:0] x_21;
	input [WIDTH-1:0] x_22;
	input [WIDTH-1:0] x_23;
	input [WIDTH-1:0] x_24;
	input [WIDTH-1:0] x_25;
	input [WIDTH-1:0] x_26;
	input [WIDTH-1:0] x_27;
	input [WIDTH-1:0] x_28;
	input [WIDTH-1:0] x_29;
	input [WIDTH-1:0] x_30;
	input [WIDTH-1:0] x_31;
	input [WIDTH-1:0] x_32;
	input [WIDTH-1:0] x_33;
	input [WIDTH-1:0] x_34;
	input [WIDTH-1:0] x_35;
	input [WIDTH-1:0] x_36;
	input [WIDTH-1:0] x_37;
	input [WIDTH-1:0] x_38;
	input [WIDTH-1:0] x_39;
	input [WIDTH-1:0] x_40;
	input [WIDTH-1:0] x_41;
	input [WIDTH-1:0] x_42;
	input [WIDTH-1:0] x_43;
	input [WIDTH-1:0] x_44;
	input [WIDTH-1:0] x_45;
	input [WIDTH-1:0] x_46;
	input [WIDTH-1:0] x_47;
	input [WIDTH-1:0] x_48;
	input [WIDTH-1:0] x_49;
	input [WIDTH-1:0] x_50;
	input [WIDTH-1:0] x_51;
	input [WIDTH-1:0] x_52;
	input [WIDTH-1:0] x_53;
	input [WIDTH-1:0] x_54;
	input [WIDTH-1:0] x_55;
	input [WIDTH-1:0] x_56;
	input [WIDTH-1:0] x_57;
	input [WIDTH-1:0] x_58;
	input [WIDTH-1:0] x_59;
	input [WIDTH-1:0] x_60;
	input [WIDTH-1:0] x_61;
	input [WIDTH-1:0] x_62;
	input [WIDTH-1:0] x_63;
	input [WIDTH-1:0] x_64;
	input [WIDTH-1:0] x_65;
	input [WIDTH-1:0] x_66;
	input [WIDTH-1:0] x_67;
	input [WIDTH-1:0] x_68;
	input [WIDTH-1:0] x_69;
	input [WIDTH-1:0] x_70;
	input [WIDTH-1:0] x_71;
	input [WIDTH-1:0] x_72;
	input [WIDTH-1:0] x_73;
	input [WIDTH-1:0] x_74;
	input [WIDTH-1:0] x_75;
	input [WIDTH-1:0] x_76;
	input [WIDTH-1:0] x_77;
	input [WIDTH-1:0] x_78;
	input [WIDTH-1:0] x_79;
	input [WIDTH-1:0] x_80;
	input [WIDTH-1:0] x_81;
	input [WIDTH-1:0] x_82;
	input [WIDTH-1:0] x_83;
	output [WIDTH-1:0] z_0;
	output [WIDTH-1:0] z_1;
	output [WIDTH-1:0] z_2;
	output [WIDTH-1:0] z_3;
	output [WIDTH-1:0] z_4;
	output [WIDTH-1:0] z_5;
	output [WIDTH-1:0] z_6;
	output [WIDTH-1:0] z_7;
	output [WIDTH-1:0] z_8;
	output [WIDTH-1:0] z_9;
	wire [WIDTH*2-1+0:0] tmp00_0_0;
	wire [WIDTH*2-1+0:0] tmp00_0_1;
	wire [WIDTH*2-1+0:0] tmp00_0_2;
	wire [WIDTH*2-1+0:0] tmp00_0_3;
	wire [WIDTH*2-1+0:0] tmp00_0_4;
	wire [WIDTH*2-1+0:0] tmp00_0_5;
	wire [WIDTH*2-1+0:0] tmp00_0_6;
	wire [WIDTH*2-1+0:0] tmp00_0_7;
	wire [WIDTH*2-1+0:0] tmp00_0_8;
	wire [WIDTH*2-1+0:0] tmp00_0_9;
	wire [WIDTH*2-1+0:0] tmp00_1_0;
	wire [WIDTH*2-1+0:0] tmp00_1_1;
	wire [WIDTH*2-1+0:0] tmp00_1_2;
	wire [WIDTH*2-1+0:0] tmp00_1_3;
	wire [WIDTH*2-1+0:0] tmp00_1_4;
	wire [WIDTH*2-1+0:0] tmp00_1_5;
	wire [WIDTH*2-1+0:0] tmp00_1_6;
	wire [WIDTH*2-1+0:0] tmp00_1_7;
	wire [WIDTH*2-1+0:0] tmp00_1_8;
	wire [WIDTH*2-1+0:0] tmp00_1_9;
	wire [WIDTH*2-1+0:0] tmp00_2_0;
	wire [WIDTH*2-1+0:0] tmp00_2_1;
	wire [WIDTH*2-1+0:0] tmp00_2_2;
	wire [WIDTH*2-1+0:0] tmp00_2_3;
	wire [WIDTH*2-1+0:0] tmp00_2_4;
	wire [WIDTH*2-1+0:0] tmp00_2_5;
	wire [WIDTH*2-1+0:0] tmp00_2_6;
	wire [WIDTH*2-1+0:0] tmp00_2_7;
	wire [WIDTH*2-1+0:0] tmp00_2_8;
	wire [WIDTH*2-1+0:0] tmp00_2_9;
	wire [WIDTH*2-1+0:0] tmp00_3_0;
	wire [WIDTH*2-1+0:0] tmp00_3_1;
	wire [WIDTH*2-1+0:0] tmp00_3_2;
	wire [WIDTH*2-1+0:0] tmp00_3_3;
	wire [WIDTH*2-1+0:0] tmp00_3_4;
	wire [WIDTH*2-1+0:0] tmp00_3_5;
	wire [WIDTH*2-1+0:0] tmp00_3_6;
	wire [WIDTH*2-1+0:0] tmp00_3_7;
	wire [WIDTH*2-1+0:0] tmp00_3_8;
	wire [WIDTH*2-1+0:0] tmp00_3_9;
	wire [WIDTH*2-1+0:0] tmp00_4_0;
	wire [WIDTH*2-1+0:0] tmp00_4_1;
	wire [WIDTH*2-1+0:0] tmp00_4_2;
	wire [WIDTH*2-1+0:0] tmp00_4_3;
	wire [WIDTH*2-1+0:0] tmp00_4_4;
	wire [WIDTH*2-1+0:0] tmp00_4_5;
	wire [WIDTH*2-1+0:0] tmp00_4_6;
	wire [WIDTH*2-1+0:0] tmp00_4_7;
	wire [WIDTH*2-1+0:0] tmp00_4_8;
	wire [WIDTH*2-1+0:0] tmp00_4_9;
	wire [WIDTH*2-1+0:0] tmp00_5_0;
	wire [WIDTH*2-1+0:0] tmp00_5_1;
	wire [WIDTH*2-1+0:0] tmp00_5_2;
	wire [WIDTH*2-1+0:0] tmp00_5_3;
	wire [WIDTH*2-1+0:0] tmp00_5_4;
	wire [WIDTH*2-1+0:0] tmp00_5_5;
	wire [WIDTH*2-1+0:0] tmp00_5_6;
	wire [WIDTH*2-1+0:0] tmp00_5_7;
	wire [WIDTH*2-1+0:0] tmp00_5_8;
	wire [WIDTH*2-1+0:0] tmp00_5_9;
	wire [WIDTH*2-1+0:0] tmp00_6_0;
	wire [WIDTH*2-1+0:0] tmp00_6_1;
	wire [WIDTH*2-1+0:0] tmp00_6_2;
	wire [WIDTH*2-1+0:0] tmp00_6_3;
	wire [WIDTH*2-1+0:0] tmp00_6_4;
	wire [WIDTH*2-1+0:0] tmp00_6_5;
	wire [WIDTH*2-1+0:0] tmp00_6_6;
	wire [WIDTH*2-1+0:0] tmp00_6_7;
	wire [WIDTH*2-1+0:0] tmp00_6_8;
	wire [WIDTH*2-1+0:0] tmp00_6_9;
	wire [WIDTH*2-1+0:0] tmp00_7_0;
	wire [WIDTH*2-1+0:0] tmp00_7_1;
	wire [WIDTH*2-1+0:0] tmp00_7_2;
	wire [WIDTH*2-1+0:0] tmp00_7_3;
	wire [WIDTH*2-1+0:0] tmp00_7_4;
	wire [WIDTH*2-1+0:0] tmp00_7_5;
	wire [WIDTH*2-1+0:0] tmp00_7_6;
	wire [WIDTH*2-1+0:0] tmp00_7_7;
	wire [WIDTH*2-1+0:0] tmp00_7_8;
	wire [WIDTH*2-1+0:0] tmp00_7_9;
	wire [WIDTH*2-1+0:0] tmp00_8_0;
	wire [WIDTH*2-1+0:0] tmp00_8_1;
	wire [WIDTH*2-1+0:0] tmp00_8_2;
	wire [WIDTH*2-1+0:0] tmp00_8_3;
	wire [WIDTH*2-1+0:0] tmp00_8_4;
	wire [WIDTH*2-1+0:0] tmp00_8_5;
	wire [WIDTH*2-1+0:0] tmp00_8_6;
	wire [WIDTH*2-1+0:0] tmp00_8_7;
	wire [WIDTH*2-1+0:0] tmp00_8_8;
	wire [WIDTH*2-1+0:0] tmp00_8_9;
	wire [WIDTH*2-1+0:0] tmp00_9_0;
	wire [WIDTH*2-1+0:0] tmp00_9_1;
	wire [WIDTH*2-1+0:0] tmp00_9_2;
	wire [WIDTH*2-1+0:0] tmp00_9_3;
	wire [WIDTH*2-1+0:0] tmp00_9_4;
	wire [WIDTH*2-1+0:0] tmp00_9_5;
	wire [WIDTH*2-1+0:0] tmp00_9_6;
	wire [WIDTH*2-1+0:0] tmp00_9_7;
	wire [WIDTH*2-1+0:0] tmp00_9_8;
	wire [WIDTH*2-1+0:0] tmp00_9_9;
	wire [WIDTH*2-1+0:0] tmp00_10_0;
	wire [WIDTH*2-1+0:0] tmp00_10_1;
	wire [WIDTH*2-1+0:0] tmp00_10_2;
	wire [WIDTH*2-1+0:0] tmp00_10_3;
	wire [WIDTH*2-1+0:0] tmp00_10_4;
	wire [WIDTH*2-1+0:0] tmp00_10_5;
	wire [WIDTH*2-1+0:0] tmp00_10_6;
	wire [WIDTH*2-1+0:0] tmp00_10_7;
	wire [WIDTH*2-1+0:0] tmp00_10_8;
	wire [WIDTH*2-1+0:0] tmp00_10_9;
	wire [WIDTH*2-1+0:0] tmp00_11_0;
	wire [WIDTH*2-1+0:0] tmp00_11_1;
	wire [WIDTH*2-1+0:0] tmp00_11_2;
	wire [WIDTH*2-1+0:0] tmp00_11_3;
	wire [WIDTH*2-1+0:0] tmp00_11_4;
	wire [WIDTH*2-1+0:0] tmp00_11_5;
	wire [WIDTH*2-1+0:0] tmp00_11_6;
	wire [WIDTH*2-1+0:0] tmp00_11_7;
	wire [WIDTH*2-1+0:0] tmp00_11_8;
	wire [WIDTH*2-1+0:0] tmp00_11_9;
	wire [WIDTH*2-1+0:0] tmp00_12_0;
	wire [WIDTH*2-1+0:0] tmp00_12_1;
	wire [WIDTH*2-1+0:0] tmp00_12_2;
	wire [WIDTH*2-1+0:0] tmp00_12_3;
	wire [WIDTH*2-1+0:0] tmp00_12_4;
	wire [WIDTH*2-1+0:0] tmp00_12_5;
	wire [WIDTH*2-1+0:0] tmp00_12_6;
	wire [WIDTH*2-1+0:0] tmp00_12_7;
	wire [WIDTH*2-1+0:0] tmp00_12_8;
	wire [WIDTH*2-1+0:0] tmp00_12_9;
	wire [WIDTH*2-1+0:0] tmp00_13_0;
	wire [WIDTH*2-1+0:0] tmp00_13_1;
	wire [WIDTH*2-1+0:0] tmp00_13_2;
	wire [WIDTH*2-1+0:0] tmp00_13_3;
	wire [WIDTH*2-1+0:0] tmp00_13_4;
	wire [WIDTH*2-1+0:0] tmp00_13_5;
	wire [WIDTH*2-1+0:0] tmp00_13_6;
	wire [WIDTH*2-1+0:0] tmp00_13_7;
	wire [WIDTH*2-1+0:0] tmp00_13_8;
	wire [WIDTH*2-1+0:0] tmp00_13_9;
	wire [WIDTH*2-1+0:0] tmp00_14_0;
	wire [WIDTH*2-1+0:0] tmp00_14_1;
	wire [WIDTH*2-1+0:0] tmp00_14_2;
	wire [WIDTH*2-1+0:0] tmp00_14_3;
	wire [WIDTH*2-1+0:0] tmp00_14_4;
	wire [WIDTH*2-1+0:0] tmp00_14_5;
	wire [WIDTH*2-1+0:0] tmp00_14_6;
	wire [WIDTH*2-1+0:0] tmp00_14_7;
	wire [WIDTH*2-1+0:0] tmp00_14_8;
	wire [WIDTH*2-1+0:0] tmp00_14_9;
	wire [WIDTH*2-1+0:0] tmp00_15_0;
	wire [WIDTH*2-1+0:0] tmp00_15_1;
	wire [WIDTH*2-1+0:0] tmp00_15_2;
	wire [WIDTH*2-1+0:0] tmp00_15_3;
	wire [WIDTH*2-1+0:0] tmp00_15_4;
	wire [WIDTH*2-1+0:0] tmp00_15_5;
	wire [WIDTH*2-1+0:0] tmp00_15_6;
	wire [WIDTH*2-1+0:0] tmp00_15_7;
	wire [WIDTH*2-1+0:0] tmp00_15_8;
	wire [WIDTH*2-1+0:0] tmp00_15_9;
	wire [WIDTH*2-1+0:0] tmp00_16_0;
	wire [WIDTH*2-1+0:0] tmp00_16_1;
	wire [WIDTH*2-1+0:0] tmp00_16_2;
	wire [WIDTH*2-1+0:0] tmp00_16_3;
	wire [WIDTH*2-1+0:0] tmp00_16_4;
	wire [WIDTH*2-1+0:0] tmp00_16_5;
	wire [WIDTH*2-1+0:0] tmp00_16_6;
	wire [WIDTH*2-1+0:0] tmp00_16_7;
	wire [WIDTH*2-1+0:0] tmp00_16_8;
	wire [WIDTH*2-1+0:0] tmp00_16_9;
	wire [WIDTH*2-1+0:0] tmp00_17_0;
	wire [WIDTH*2-1+0:0] tmp00_17_1;
	wire [WIDTH*2-1+0:0] tmp00_17_2;
	wire [WIDTH*2-1+0:0] tmp00_17_3;
	wire [WIDTH*2-1+0:0] tmp00_17_4;
	wire [WIDTH*2-1+0:0] tmp00_17_5;
	wire [WIDTH*2-1+0:0] tmp00_17_6;
	wire [WIDTH*2-1+0:0] tmp00_17_7;
	wire [WIDTH*2-1+0:0] tmp00_17_8;
	wire [WIDTH*2-1+0:0] tmp00_17_9;
	wire [WIDTH*2-1+0:0] tmp00_18_0;
	wire [WIDTH*2-1+0:0] tmp00_18_1;
	wire [WIDTH*2-1+0:0] tmp00_18_2;
	wire [WIDTH*2-1+0:0] tmp00_18_3;
	wire [WIDTH*2-1+0:0] tmp00_18_4;
	wire [WIDTH*2-1+0:0] tmp00_18_5;
	wire [WIDTH*2-1+0:0] tmp00_18_6;
	wire [WIDTH*2-1+0:0] tmp00_18_7;
	wire [WIDTH*2-1+0:0] tmp00_18_8;
	wire [WIDTH*2-1+0:0] tmp00_18_9;
	wire [WIDTH*2-1+0:0] tmp00_19_0;
	wire [WIDTH*2-1+0:0] tmp00_19_1;
	wire [WIDTH*2-1+0:0] tmp00_19_2;
	wire [WIDTH*2-1+0:0] tmp00_19_3;
	wire [WIDTH*2-1+0:0] tmp00_19_4;
	wire [WIDTH*2-1+0:0] tmp00_19_5;
	wire [WIDTH*2-1+0:0] tmp00_19_6;
	wire [WIDTH*2-1+0:0] tmp00_19_7;
	wire [WIDTH*2-1+0:0] tmp00_19_8;
	wire [WIDTH*2-1+0:0] tmp00_19_9;
	wire [WIDTH*2-1+0:0] tmp00_20_0;
	wire [WIDTH*2-1+0:0] tmp00_20_1;
	wire [WIDTH*2-1+0:0] tmp00_20_2;
	wire [WIDTH*2-1+0:0] tmp00_20_3;
	wire [WIDTH*2-1+0:0] tmp00_20_4;
	wire [WIDTH*2-1+0:0] tmp00_20_5;
	wire [WIDTH*2-1+0:0] tmp00_20_6;
	wire [WIDTH*2-1+0:0] tmp00_20_7;
	wire [WIDTH*2-1+0:0] tmp00_20_8;
	wire [WIDTH*2-1+0:0] tmp00_20_9;
	wire [WIDTH*2-1+0:0] tmp00_21_0;
	wire [WIDTH*2-1+0:0] tmp00_21_1;
	wire [WIDTH*2-1+0:0] tmp00_21_2;
	wire [WIDTH*2-1+0:0] tmp00_21_3;
	wire [WIDTH*2-1+0:0] tmp00_21_4;
	wire [WIDTH*2-1+0:0] tmp00_21_5;
	wire [WIDTH*2-1+0:0] tmp00_21_6;
	wire [WIDTH*2-1+0:0] tmp00_21_7;
	wire [WIDTH*2-1+0:0] tmp00_21_8;
	wire [WIDTH*2-1+0:0] tmp00_21_9;
	wire [WIDTH*2-1+0:0] tmp00_22_0;
	wire [WIDTH*2-1+0:0] tmp00_22_1;
	wire [WIDTH*2-1+0:0] tmp00_22_2;
	wire [WIDTH*2-1+0:0] tmp00_22_3;
	wire [WIDTH*2-1+0:0] tmp00_22_4;
	wire [WIDTH*2-1+0:0] tmp00_22_5;
	wire [WIDTH*2-1+0:0] tmp00_22_6;
	wire [WIDTH*2-1+0:0] tmp00_22_7;
	wire [WIDTH*2-1+0:0] tmp00_22_8;
	wire [WIDTH*2-1+0:0] tmp00_22_9;
	wire [WIDTH*2-1+0:0] tmp00_23_0;
	wire [WIDTH*2-1+0:0] tmp00_23_1;
	wire [WIDTH*2-1+0:0] tmp00_23_2;
	wire [WIDTH*2-1+0:0] tmp00_23_3;
	wire [WIDTH*2-1+0:0] tmp00_23_4;
	wire [WIDTH*2-1+0:0] tmp00_23_5;
	wire [WIDTH*2-1+0:0] tmp00_23_6;
	wire [WIDTH*2-1+0:0] tmp00_23_7;
	wire [WIDTH*2-1+0:0] tmp00_23_8;
	wire [WIDTH*2-1+0:0] tmp00_23_9;
	wire [WIDTH*2-1+0:0] tmp00_24_0;
	wire [WIDTH*2-1+0:0] tmp00_24_1;
	wire [WIDTH*2-1+0:0] tmp00_24_2;
	wire [WIDTH*2-1+0:0] tmp00_24_3;
	wire [WIDTH*2-1+0:0] tmp00_24_4;
	wire [WIDTH*2-1+0:0] tmp00_24_5;
	wire [WIDTH*2-1+0:0] tmp00_24_6;
	wire [WIDTH*2-1+0:0] tmp00_24_7;
	wire [WIDTH*2-1+0:0] tmp00_24_8;
	wire [WIDTH*2-1+0:0] tmp00_24_9;
	wire [WIDTH*2-1+0:0] tmp00_25_0;
	wire [WIDTH*2-1+0:0] tmp00_25_1;
	wire [WIDTH*2-1+0:0] tmp00_25_2;
	wire [WIDTH*2-1+0:0] tmp00_25_3;
	wire [WIDTH*2-1+0:0] tmp00_25_4;
	wire [WIDTH*2-1+0:0] tmp00_25_5;
	wire [WIDTH*2-1+0:0] tmp00_25_6;
	wire [WIDTH*2-1+0:0] tmp00_25_7;
	wire [WIDTH*2-1+0:0] tmp00_25_8;
	wire [WIDTH*2-1+0:0] tmp00_25_9;
	wire [WIDTH*2-1+0:0] tmp00_26_0;
	wire [WIDTH*2-1+0:0] tmp00_26_1;
	wire [WIDTH*2-1+0:0] tmp00_26_2;
	wire [WIDTH*2-1+0:0] tmp00_26_3;
	wire [WIDTH*2-1+0:0] tmp00_26_4;
	wire [WIDTH*2-1+0:0] tmp00_26_5;
	wire [WIDTH*2-1+0:0] tmp00_26_6;
	wire [WIDTH*2-1+0:0] tmp00_26_7;
	wire [WIDTH*2-1+0:0] tmp00_26_8;
	wire [WIDTH*2-1+0:0] tmp00_26_9;
	wire [WIDTH*2-1+0:0] tmp00_27_0;
	wire [WIDTH*2-1+0:0] tmp00_27_1;
	wire [WIDTH*2-1+0:0] tmp00_27_2;
	wire [WIDTH*2-1+0:0] tmp00_27_3;
	wire [WIDTH*2-1+0:0] tmp00_27_4;
	wire [WIDTH*2-1+0:0] tmp00_27_5;
	wire [WIDTH*2-1+0:0] tmp00_27_6;
	wire [WIDTH*2-1+0:0] tmp00_27_7;
	wire [WIDTH*2-1+0:0] tmp00_27_8;
	wire [WIDTH*2-1+0:0] tmp00_27_9;
	wire [WIDTH*2-1+0:0] tmp00_28_0;
	wire [WIDTH*2-1+0:0] tmp00_28_1;
	wire [WIDTH*2-1+0:0] tmp00_28_2;
	wire [WIDTH*2-1+0:0] tmp00_28_3;
	wire [WIDTH*2-1+0:0] tmp00_28_4;
	wire [WIDTH*2-1+0:0] tmp00_28_5;
	wire [WIDTH*2-1+0:0] tmp00_28_6;
	wire [WIDTH*2-1+0:0] tmp00_28_7;
	wire [WIDTH*2-1+0:0] tmp00_28_8;
	wire [WIDTH*2-1+0:0] tmp00_28_9;
	wire [WIDTH*2-1+0:0] tmp00_29_0;
	wire [WIDTH*2-1+0:0] tmp00_29_1;
	wire [WIDTH*2-1+0:0] tmp00_29_2;
	wire [WIDTH*2-1+0:0] tmp00_29_3;
	wire [WIDTH*2-1+0:0] tmp00_29_4;
	wire [WIDTH*2-1+0:0] tmp00_29_5;
	wire [WIDTH*2-1+0:0] tmp00_29_6;
	wire [WIDTH*2-1+0:0] tmp00_29_7;
	wire [WIDTH*2-1+0:0] tmp00_29_8;
	wire [WIDTH*2-1+0:0] tmp00_29_9;
	wire [WIDTH*2-1+0:0] tmp00_30_0;
	wire [WIDTH*2-1+0:0] tmp00_30_1;
	wire [WIDTH*2-1+0:0] tmp00_30_2;
	wire [WIDTH*2-1+0:0] tmp00_30_3;
	wire [WIDTH*2-1+0:0] tmp00_30_4;
	wire [WIDTH*2-1+0:0] tmp00_30_5;
	wire [WIDTH*2-1+0:0] tmp00_30_6;
	wire [WIDTH*2-1+0:0] tmp00_30_7;
	wire [WIDTH*2-1+0:0] tmp00_30_8;
	wire [WIDTH*2-1+0:0] tmp00_30_9;
	wire [WIDTH*2-1+0:0] tmp00_31_0;
	wire [WIDTH*2-1+0:0] tmp00_31_1;
	wire [WIDTH*2-1+0:0] tmp00_31_2;
	wire [WIDTH*2-1+0:0] tmp00_31_3;
	wire [WIDTH*2-1+0:0] tmp00_31_4;
	wire [WIDTH*2-1+0:0] tmp00_31_5;
	wire [WIDTH*2-1+0:0] tmp00_31_6;
	wire [WIDTH*2-1+0:0] tmp00_31_7;
	wire [WIDTH*2-1+0:0] tmp00_31_8;
	wire [WIDTH*2-1+0:0] tmp00_31_9;
	wire [WIDTH*2-1+0:0] tmp00_32_0;
	wire [WIDTH*2-1+0:0] tmp00_32_1;
	wire [WIDTH*2-1+0:0] tmp00_32_2;
	wire [WIDTH*2-1+0:0] tmp00_32_3;
	wire [WIDTH*2-1+0:0] tmp00_32_4;
	wire [WIDTH*2-1+0:0] tmp00_32_5;
	wire [WIDTH*2-1+0:0] tmp00_32_6;
	wire [WIDTH*2-1+0:0] tmp00_32_7;
	wire [WIDTH*2-1+0:0] tmp00_32_8;
	wire [WIDTH*2-1+0:0] tmp00_32_9;
	wire [WIDTH*2-1+0:0] tmp00_33_0;
	wire [WIDTH*2-1+0:0] tmp00_33_1;
	wire [WIDTH*2-1+0:0] tmp00_33_2;
	wire [WIDTH*2-1+0:0] tmp00_33_3;
	wire [WIDTH*2-1+0:0] tmp00_33_4;
	wire [WIDTH*2-1+0:0] tmp00_33_5;
	wire [WIDTH*2-1+0:0] tmp00_33_6;
	wire [WIDTH*2-1+0:0] tmp00_33_7;
	wire [WIDTH*2-1+0:0] tmp00_33_8;
	wire [WIDTH*2-1+0:0] tmp00_33_9;
	wire [WIDTH*2-1+0:0] tmp00_34_0;
	wire [WIDTH*2-1+0:0] tmp00_34_1;
	wire [WIDTH*2-1+0:0] tmp00_34_2;
	wire [WIDTH*2-1+0:0] tmp00_34_3;
	wire [WIDTH*2-1+0:0] tmp00_34_4;
	wire [WIDTH*2-1+0:0] tmp00_34_5;
	wire [WIDTH*2-1+0:0] tmp00_34_6;
	wire [WIDTH*2-1+0:0] tmp00_34_7;
	wire [WIDTH*2-1+0:0] tmp00_34_8;
	wire [WIDTH*2-1+0:0] tmp00_34_9;
	wire [WIDTH*2-1+0:0] tmp00_35_0;
	wire [WIDTH*2-1+0:0] tmp00_35_1;
	wire [WIDTH*2-1+0:0] tmp00_35_2;
	wire [WIDTH*2-1+0:0] tmp00_35_3;
	wire [WIDTH*2-1+0:0] tmp00_35_4;
	wire [WIDTH*2-1+0:0] tmp00_35_5;
	wire [WIDTH*2-1+0:0] tmp00_35_6;
	wire [WIDTH*2-1+0:0] tmp00_35_7;
	wire [WIDTH*2-1+0:0] tmp00_35_8;
	wire [WIDTH*2-1+0:0] tmp00_35_9;
	wire [WIDTH*2-1+0:0] tmp00_36_0;
	wire [WIDTH*2-1+0:0] tmp00_36_1;
	wire [WIDTH*2-1+0:0] tmp00_36_2;
	wire [WIDTH*2-1+0:0] tmp00_36_3;
	wire [WIDTH*2-1+0:0] tmp00_36_4;
	wire [WIDTH*2-1+0:0] tmp00_36_5;
	wire [WIDTH*2-1+0:0] tmp00_36_6;
	wire [WIDTH*2-1+0:0] tmp00_36_7;
	wire [WIDTH*2-1+0:0] tmp00_36_8;
	wire [WIDTH*2-1+0:0] tmp00_36_9;
	wire [WIDTH*2-1+0:0] tmp00_37_0;
	wire [WIDTH*2-1+0:0] tmp00_37_1;
	wire [WIDTH*2-1+0:0] tmp00_37_2;
	wire [WIDTH*2-1+0:0] tmp00_37_3;
	wire [WIDTH*2-1+0:0] tmp00_37_4;
	wire [WIDTH*2-1+0:0] tmp00_37_5;
	wire [WIDTH*2-1+0:0] tmp00_37_6;
	wire [WIDTH*2-1+0:0] tmp00_37_7;
	wire [WIDTH*2-1+0:0] tmp00_37_8;
	wire [WIDTH*2-1+0:0] tmp00_37_9;
	wire [WIDTH*2-1+0:0] tmp00_38_0;
	wire [WIDTH*2-1+0:0] tmp00_38_1;
	wire [WIDTH*2-1+0:0] tmp00_38_2;
	wire [WIDTH*2-1+0:0] tmp00_38_3;
	wire [WIDTH*2-1+0:0] tmp00_38_4;
	wire [WIDTH*2-1+0:0] tmp00_38_5;
	wire [WIDTH*2-1+0:0] tmp00_38_6;
	wire [WIDTH*2-1+0:0] tmp00_38_7;
	wire [WIDTH*2-1+0:0] tmp00_38_8;
	wire [WIDTH*2-1+0:0] tmp00_38_9;
	wire [WIDTH*2-1+0:0] tmp00_39_0;
	wire [WIDTH*2-1+0:0] tmp00_39_1;
	wire [WIDTH*2-1+0:0] tmp00_39_2;
	wire [WIDTH*2-1+0:0] tmp00_39_3;
	wire [WIDTH*2-1+0:0] tmp00_39_4;
	wire [WIDTH*2-1+0:0] tmp00_39_5;
	wire [WIDTH*2-1+0:0] tmp00_39_6;
	wire [WIDTH*2-1+0:0] tmp00_39_7;
	wire [WIDTH*2-1+0:0] tmp00_39_8;
	wire [WIDTH*2-1+0:0] tmp00_39_9;
	wire [WIDTH*2-1+0:0] tmp00_40_0;
	wire [WIDTH*2-1+0:0] tmp00_40_1;
	wire [WIDTH*2-1+0:0] tmp00_40_2;
	wire [WIDTH*2-1+0:0] tmp00_40_3;
	wire [WIDTH*2-1+0:0] tmp00_40_4;
	wire [WIDTH*2-1+0:0] tmp00_40_5;
	wire [WIDTH*2-1+0:0] tmp00_40_6;
	wire [WIDTH*2-1+0:0] tmp00_40_7;
	wire [WIDTH*2-1+0:0] tmp00_40_8;
	wire [WIDTH*2-1+0:0] tmp00_40_9;
	wire [WIDTH*2-1+0:0] tmp00_41_0;
	wire [WIDTH*2-1+0:0] tmp00_41_1;
	wire [WIDTH*2-1+0:0] tmp00_41_2;
	wire [WIDTH*2-1+0:0] tmp00_41_3;
	wire [WIDTH*2-1+0:0] tmp00_41_4;
	wire [WIDTH*2-1+0:0] tmp00_41_5;
	wire [WIDTH*2-1+0:0] tmp00_41_6;
	wire [WIDTH*2-1+0:0] tmp00_41_7;
	wire [WIDTH*2-1+0:0] tmp00_41_8;
	wire [WIDTH*2-1+0:0] tmp00_41_9;
	wire [WIDTH*2-1+0:0] tmp00_42_0;
	wire [WIDTH*2-1+0:0] tmp00_42_1;
	wire [WIDTH*2-1+0:0] tmp00_42_2;
	wire [WIDTH*2-1+0:0] tmp00_42_3;
	wire [WIDTH*2-1+0:0] tmp00_42_4;
	wire [WIDTH*2-1+0:0] tmp00_42_5;
	wire [WIDTH*2-1+0:0] tmp00_42_6;
	wire [WIDTH*2-1+0:0] tmp00_42_7;
	wire [WIDTH*2-1+0:0] tmp00_42_8;
	wire [WIDTH*2-1+0:0] tmp00_42_9;
	wire [WIDTH*2-1+0:0] tmp00_43_0;
	wire [WIDTH*2-1+0:0] tmp00_43_1;
	wire [WIDTH*2-1+0:0] tmp00_43_2;
	wire [WIDTH*2-1+0:0] tmp00_43_3;
	wire [WIDTH*2-1+0:0] tmp00_43_4;
	wire [WIDTH*2-1+0:0] tmp00_43_5;
	wire [WIDTH*2-1+0:0] tmp00_43_6;
	wire [WIDTH*2-1+0:0] tmp00_43_7;
	wire [WIDTH*2-1+0:0] tmp00_43_8;
	wire [WIDTH*2-1+0:0] tmp00_43_9;
	wire [WIDTH*2-1+0:0] tmp00_44_0;
	wire [WIDTH*2-1+0:0] tmp00_44_1;
	wire [WIDTH*2-1+0:0] tmp00_44_2;
	wire [WIDTH*2-1+0:0] tmp00_44_3;
	wire [WIDTH*2-1+0:0] tmp00_44_4;
	wire [WIDTH*2-1+0:0] tmp00_44_5;
	wire [WIDTH*2-1+0:0] tmp00_44_6;
	wire [WIDTH*2-1+0:0] tmp00_44_7;
	wire [WIDTH*2-1+0:0] tmp00_44_8;
	wire [WIDTH*2-1+0:0] tmp00_44_9;
	wire [WIDTH*2-1+0:0] tmp00_45_0;
	wire [WIDTH*2-1+0:0] tmp00_45_1;
	wire [WIDTH*2-1+0:0] tmp00_45_2;
	wire [WIDTH*2-1+0:0] tmp00_45_3;
	wire [WIDTH*2-1+0:0] tmp00_45_4;
	wire [WIDTH*2-1+0:0] tmp00_45_5;
	wire [WIDTH*2-1+0:0] tmp00_45_6;
	wire [WIDTH*2-1+0:0] tmp00_45_7;
	wire [WIDTH*2-1+0:0] tmp00_45_8;
	wire [WIDTH*2-1+0:0] tmp00_45_9;
	wire [WIDTH*2-1+0:0] tmp00_46_0;
	wire [WIDTH*2-1+0:0] tmp00_46_1;
	wire [WIDTH*2-1+0:0] tmp00_46_2;
	wire [WIDTH*2-1+0:0] tmp00_46_3;
	wire [WIDTH*2-1+0:0] tmp00_46_4;
	wire [WIDTH*2-1+0:0] tmp00_46_5;
	wire [WIDTH*2-1+0:0] tmp00_46_6;
	wire [WIDTH*2-1+0:0] tmp00_46_7;
	wire [WIDTH*2-1+0:0] tmp00_46_8;
	wire [WIDTH*2-1+0:0] tmp00_46_9;
	wire [WIDTH*2-1+0:0] tmp00_47_0;
	wire [WIDTH*2-1+0:0] tmp00_47_1;
	wire [WIDTH*2-1+0:0] tmp00_47_2;
	wire [WIDTH*2-1+0:0] tmp00_47_3;
	wire [WIDTH*2-1+0:0] tmp00_47_4;
	wire [WIDTH*2-1+0:0] tmp00_47_5;
	wire [WIDTH*2-1+0:0] tmp00_47_6;
	wire [WIDTH*2-1+0:0] tmp00_47_7;
	wire [WIDTH*2-1+0:0] tmp00_47_8;
	wire [WIDTH*2-1+0:0] tmp00_47_9;
	wire [WIDTH*2-1+0:0] tmp00_48_0;
	wire [WIDTH*2-1+0:0] tmp00_48_1;
	wire [WIDTH*2-1+0:0] tmp00_48_2;
	wire [WIDTH*2-1+0:0] tmp00_48_3;
	wire [WIDTH*2-1+0:0] tmp00_48_4;
	wire [WIDTH*2-1+0:0] tmp00_48_5;
	wire [WIDTH*2-1+0:0] tmp00_48_6;
	wire [WIDTH*2-1+0:0] tmp00_48_7;
	wire [WIDTH*2-1+0:0] tmp00_48_8;
	wire [WIDTH*2-1+0:0] tmp00_48_9;
	wire [WIDTH*2-1+0:0] tmp00_49_0;
	wire [WIDTH*2-1+0:0] tmp00_49_1;
	wire [WIDTH*2-1+0:0] tmp00_49_2;
	wire [WIDTH*2-1+0:0] tmp00_49_3;
	wire [WIDTH*2-1+0:0] tmp00_49_4;
	wire [WIDTH*2-1+0:0] tmp00_49_5;
	wire [WIDTH*2-1+0:0] tmp00_49_6;
	wire [WIDTH*2-1+0:0] tmp00_49_7;
	wire [WIDTH*2-1+0:0] tmp00_49_8;
	wire [WIDTH*2-1+0:0] tmp00_49_9;
	wire [WIDTH*2-1+0:0] tmp00_50_0;
	wire [WIDTH*2-1+0:0] tmp00_50_1;
	wire [WIDTH*2-1+0:0] tmp00_50_2;
	wire [WIDTH*2-1+0:0] tmp00_50_3;
	wire [WIDTH*2-1+0:0] tmp00_50_4;
	wire [WIDTH*2-1+0:0] tmp00_50_5;
	wire [WIDTH*2-1+0:0] tmp00_50_6;
	wire [WIDTH*2-1+0:0] tmp00_50_7;
	wire [WIDTH*2-1+0:0] tmp00_50_8;
	wire [WIDTH*2-1+0:0] tmp00_50_9;
	wire [WIDTH*2-1+0:0] tmp00_51_0;
	wire [WIDTH*2-1+0:0] tmp00_51_1;
	wire [WIDTH*2-1+0:0] tmp00_51_2;
	wire [WIDTH*2-1+0:0] tmp00_51_3;
	wire [WIDTH*2-1+0:0] tmp00_51_4;
	wire [WIDTH*2-1+0:0] tmp00_51_5;
	wire [WIDTH*2-1+0:0] tmp00_51_6;
	wire [WIDTH*2-1+0:0] tmp00_51_7;
	wire [WIDTH*2-1+0:0] tmp00_51_8;
	wire [WIDTH*2-1+0:0] tmp00_51_9;
	wire [WIDTH*2-1+0:0] tmp00_52_0;
	wire [WIDTH*2-1+0:0] tmp00_52_1;
	wire [WIDTH*2-1+0:0] tmp00_52_2;
	wire [WIDTH*2-1+0:0] tmp00_52_3;
	wire [WIDTH*2-1+0:0] tmp00_52_4;
	wire [WIDTH*2-1+0:0] tmp00_52_5;
	wire [WIDTH*2-1+0:0] tmp00_52_6;
	wire [WIDTH*2-1+0:0] tmp00_52_7;
	wire [WIDTH*2-1+0:0] tmp00_52_8;
	wire [WIDTH*2-1+0:0] tmp00_52_9;
	wire [WIDTH*2-1+0:0] tmp00_53_0;
	wire [WIDTH*2-1+0:0] tmp00_53_1;
	wire [WIDTH*2-1+0:0] tmp00_53_2;
	wire [WIDTH*2-1+0:0] tmp00_53_3;
	wire [WIDTH*2-1+0:0] tmp00_53_4;
	wire [WIDTH*2-1+0:0] tmp00_53_5;
	wire [WIDTH*2-1+0:0] tmp00_53_6;
	wire [WIDTH*2-1+0:0] tmp00_53_7;
	wire [WIDTH*2-1+0:0] tmp00_53_8;
	wire [WIDTH*2-1+0:0] tmp00_53_9;
	wire [WIDTH*2-1+0:0] tmp00_54_0;
	wire [WIDTH*2-1+0:0] tmp00_54_1;
	wire [WIDTH*2-1+0:0] tmp00_54_2;
	wire [WIDTH*2-1+0:0] tmp00_54_3;
	wire [WIDTH*2-1+0:0] tmp00_54_4;
	wire [WIDTH*2-1+0:0] tmp00_54_5;
	wire [WIDTH*2-1+0:0] tmp00_54_6;
	wire [WIDTH*2-1+0:0] tmp00_54_7;
	wire [WIDTH*2-1+0:0] tmp00_54_8;
	wire [WIDTH*2-1+0:0] tmp00_54_9;
	wire [WIDTH*2-1+0:0] tmp00_55_0;
	wire [WIDTH*2-1+0:0] tmp00_55_1;
	wire [WIDTH*2-1+0:0] tmp00_55_2;
	wire [WIDTH*2-1+0:0] tmp00_55_3;
	wire [WIDTH*2-1+0:0] tmp00_55_4;
	wire [WIDTH*2-1+0:0] tmp00_55_5;
	wire [WIDTH*2-1+0:0] tmp00_55_6;
	wire [WIDTH*2-1+0:0] tmp00_55_7;
	wire [WIDTH*2-1+0:0] tmp00_55_8;
	wire [WIDTH*2-1+0:0] tmp00_55_9;
	wire [WIDTH*2-1+0:0] tmp00_56_0;
	wire [WIDTH*2-1+0:0] tmp00_56_1;
	wire [WIDTH*2-1+0:0] tmp00_56_2;
	wire [WIDTH*2-1+0:0] tmp00_56_3;
	wire [WIDTH*2-1+0:0] tmp00_56_4;
	wire [WIDTH*2-1+0:0] tmp00_56_5;
	wire [WIDTH*2-1+0:0] tmp00_56_6;
	wire [WIDTH*2-1+0:0] tmp00_56_7;
	wire [WIDTH*2-1+0:0] tmp00_56_8;
	wire [WIDTH*2-1+0:0] tmp00_56_9;
	wire [WIDTH*2-1+0:0] tmp00_57_0;
	wire [WIDTH*2-1+0:0] tmp00_57_1;
	wire [WIDTH*2-1+0:0] tmp00_57_2;
	wire [WIDTH*2-1+0:0] tmp00_57_3;
	wire [WIDTH*2-1+0:0] tmp00_57_4;
	wire [WIDTH*2-1+0:0] tmp00_57_5;
	wire [WIDTH*2-1+0:0] tmp00_57_6;
	wire [WIDTH*2-1+0:0] tmp00_57_7;
	wire [WIDTH*2-1+0:0] tmp00_57_8;
	wire [WIDTH*2-1+0:0] tmp00_57_9;
	wire [WIDTH*2-1+0:0] tmp00_58_0;
	wire [WIDTH*2-1+0:0] tmp00_58_1;
	wire [WIDTH*2-1+0:0] tmp00_58_2;
	wire [WIDTH*2-1+0:0] tmp00_58_3;
	wire [WIDTH*2-1+0:0] tmp00_58_4;
	wire [WIDTH*2-1+0:0] tmp00_58_5;
	wire [WIDTH*2-1+0:0] tmp00_58_6;
	wire [WIDTH*2-1+0:0] tmp00_58_7;
	wire [WIDTH*2-1+0:0] tmp00_58_8;
	wire [WIDTH*2-1+0:0] tmp00_58_9;
	wire [WIDTH*2-1+0:0] tmp00_59_0;
	wire [WIDTH*2-1+0:0] tmp00_59_1;
	wire [WIDTH*2-1+0:0] tmp00_59_2;
	wire [WIDTH*2-1+0:0] tmp00_59_3;
	wire [WIDTH*2-1+0:0] tmp00_59_4;
	wire [WIDTH*2-1+0:0] tmp00_59_5;
	wire [WIDTH*2-1+0:0] tmp00_59_6;
	wire [WIDTH*2-1+0:0] tmp00_59_7;
	wire [WIDTH*2-1+0:0] tmp00_59_8;
	wire [WIDTH*2-1+0:0] tmp00_59_9;
	wire [WIDTH*2-1+0:0] tmp00_60_0;
	wire [WIDTH*2-1+0:0] tmp00_60_1;
	wire [WIDTH*2-1+0:0] tmp00_60_2;
	wire [WIDTH*2-1+0:0] tmp00_60_3;
	wire [WIDTH*2-1+0:0] tmp00_60_4;
	wire [WIDTH*2-1+0:0] tmp00_60_5;
	wire [WIDTH*2-1+0:0] tmp00_60_6;
	wire [WIDTH*2-1+0:0] tmp00_60_7;
	wire [WIDTH*2-1+0:0] tmp00_60_8;
	wire [WIDTH*2-1+0:0] tmp00_60_9;
	wire [WIDTH*2-1+0:0] tmp00_61_0;
	wire [WIDTH*2-1+0:0] tmp00_61_1;
	wire [WIDTH*2-1+0:0] tmp00_61_2;
	wire [WIDTH*2-1+0:0] tmp00_61_3;
	wire [WIDTH*2-1+0:0] tmp00_61_4;
	wire [WIDTH*2-1+0:0] tmp00_61_5;
	wire [WIDTH*2-1+0:0] tmp00_61_6;
	wire [WIDTH*2-1+0:0] tmp00_61_7;
	wire [WIDTH*2-1+0:0] tmp00_61_8;
	wire [WIDTH*2-1+0:0] tmp00_61_9;
	wire [WIDTH*2-1+0:0] tmp00_62_0;
	wire [WIDTH*2-1+0:0] tmp00_62_1;
	wire [WIDTH*2-1+0:0] tmp00_62_2;
	wire [WIDTH*2-1+0:0] tmp00_62_3;
	wire [WIDTH*2-1+0:0] tmp00_62_4;
	wire [WIDTH*2-1+0:0] tmp00_62_5;
	wire [WIDTH*2-1+0:0] tmp00_62_6;
	wire [WIDTH*2-1+0:0] tmp00_62_7;
	wire [WIDTH*2-1+0:0] tmp00_62_8;
	wire [WIDTH*2-1+0:0] tmp00_62_9;
	wire [WIDTH*2-1+0:0] tmp00_63_0;
	wire [WIDTH*2-1+0:0] tmp00_63_1;
	wire [WIDTH*2-1+0:0] tmp00_63_2;
	wire [WIDTH*2-1+0:0] tmp00_63_3;
	wire [WIDTH*2-1+0:0] tmp00_63_4;
	wire [WIDTH*2-1+0:0] tmp00_63_5;
	wire [WIDTH*2-1+0:0] tmp00_63_6;
	wire [WIDTH*2-1+0:0] tmp00_63_7;
	wire [WIDTH*2-1+0:0] tmp00_63_8;
	wire [WIDTH*2-1+0:0] tmp00_63_9;
	wire [WIDTH*2-1+0:0] tmp00_64_0;
	wire [WIDTH*2-1+0:0] tmp00_64_1;
	wire [WIDTH*2-1+0:0] tmp00_64_2;
	wire [WIDTH*2-1+0:0] tmp00_64_3;
	wire [WIDTH*2-1+0:0] tmp00_64_4;
	wire [WIDTH*2-1+0:0] tmp00_64_5;
	wire [WIDTH*2-1+0:0] tmp00_64_6;
	wire [WIDTH*2-1+0:0] tmp00_64_7;
	wire [WIDTH*2-1+0:0] tmp00_64_8;
	wire [WIDTH*2-1+0:0] tmp00_64_9;
	wire [WIDTH*2-1+0:0] tmp00_65_0;
	wire [WIDTH*2-1+0:0] tmp00_65_1;
	wire [WIDTH*2-1+0:0] tmp00_65_2;
	wire [WIDTH*2-1+0:0] tmp00_65_3;
	wire [WIDTH*2-1+0:0] tmp00_65_4;
	wire [WIDTH*2-1+0:0] tmp00_65_5;
	wire [WIDTH*2-1+0:0] tmp00_65_6;
	wire [WIDTH*2-1+0:0] tmp00_65_7;
	wire [WIDTH*2-1+0:0] tmp00_65_8;
	wire [WIDTH*2-1+0:0] tmp00_65_9;
	wire [WIDTH*2-1+0:0] tmp00_66_0;
	wire [WIDTH*2-1+0:0] tmp00_66_1;
	wire [WIDTH*2-1+0:0] tmp00_66_2;
	wire [WIDTH*2-1+0:0] tmp00_66_3;
	wire [WIDTH*2-1+0:0] tmp00_66_4;
	wire [WIDTH*2-1+0:0] tmp00_66_5;
	wire [WIDTH*2-1+0:0] tmp00_66_6;
	wire [WIDTH*2-1+0:0] tmp00_66_7;
	wire [WIDTH*2-1+0:0] tmp00_66_8;
	wire [WIDTH*2-1+0:0] tmp00_66_9;
	wire [WIDTH*2-1+0:0] tmp00_67_0;
	wire [WIDTH*2-1+0:0] tmp00_67_1;
	wire [WIDTH*2-1+0:0] tmp00_67_2;
	wire [WIDTH*2-1+0:0] tmp00_67_3;
	wire [WIDTH*2-1+0:0] tmp00_67_4;
	wire [WIDTH*2-1+0:0] tmp00_67_5;
	wire [WIDTH*2-1+0:0] tmp00_67_6;
	wire [WIDTH*2-1+0:0] tmp00_67_7;
	wire [WIDTH*2-1+0:0] tmp00_67_8;
	wire [WIDTH*2-1+0:0] tmp00_67_9;
	wire [WIDTH*2-1+0:0] tmp00_68_0;
	wire [WIDTH*2-1+0:0] tmp00_68_1;
	wire [WIDTH*2-1+0:0] tmp00_68_2;
	wire [WIDTH*2-1+0:0] tmp00_68_3;
	wire [WIDTH*2-1+0:0] tmp00_68_4;
	wire [WIDTH*2-1+0:0] tmp00_68_5;
	wire [WIDTH*2-1+0:0] tmp00_68_6;
	wire [WIDTH*2-1+0:0] tmp00_68_7;
	wire [WIDTH*2-1+0:0] tmp00_68_8;
	wire [WIDTH*2-1+0:0] tmp00_68_9;
	wire [WIDTH*2-1+0:0] tmp00_69_0;
	wire [WIDTH*2-1+0:0] tmp00_69_1;
	wire [WIDTH*2-1+0:0] tmp00_69_2;
	wire [WIDTH*2-1+0:0] tmp00_69_3;
	wire [WIDTH*2-1+0:0] tmp00_69_4;
	wire [WIDTH*2-1+0:0] tmp00_69_5;
	wire [WIDTH*2-1+0:0] tmp00_69_6;
	wire [WIDTH*2-1+0:0] tmp00_69_7;
	wire [WIDTH*2-1+0:0] tmp00_69_8;
	wire [WIDTH*2-1+0:0] tmp00_69_9;
	wire [WIDTH*2-1+0:0] tmp00_70_0;
	wire [WIDTH*2-1+0:0] tmp00_70_1;
	wire [WIDTH*2-1+0:0] tmp00_70_2;
	wire [WIDTH*2-1+0:0] tmp00_70_3;
	wire [WIDTH*2-1+0:0] tmp00_70_4;
	wire [WIDTH*2-1+0:0] tmp00_70_5;
	wire [WIDTH*2-1+0:0] tmp00_70_6;
	wire [WIDTH*2-1+0:0] tmp00_70_7;
	wire [WIDTH*2-1+0:0] tmp00_70_8;
	wire [WIDTH*2-1+0:0] tmp00_70_9;
	wire [WIDTH*2-1+0:0] tmp00_71_0;
	wire [WIDTH*2-1+0:0] tmp00_71_1;
	wire [WIDTH*2-1+0:0] tmp00_71_2;
	wire [WIDTH*2-1+0:0] tmp00_71_3;
	wire [WIDTH*2-1+0:0] tmp00_71_4;
	wire [WIDTH*2-1+0:0] tmp00_71_5;
	wire [WIDTH*2-1+0:0] tmp00_71_6;
	wire [WIDTH*2-1+0:0] tmp00_71_7;
	wire [WIDTH*2-1+0:0] tmp00_71_8;
	wire [WIDTH*2-1+0:0] tmp00_71_9;
	wire [WIDTH*2-1+0:0] tmp00_72_0;
	wire [WIDTH*2-1+0:0] tmp00_72_1;
	wire [WIDTH*2-1+0:0] tmp00_72_2;
	wire [WIDTH*2-1+0:0] tmp00_72_3;
	wire [WIDTH*2-1+0:0] tmp00_72_4;
	wire [WIDTH*2-1+0:0] tmp00_72_5;
	wire [WIDTH*2-1+0:0] tmp00_72_6;
	wire [WIDTH*2-1+0:0] tmp00_72_7;
	wire [WIDTH*2-1+0:0] tmp00_72_8;
	wire [WIDTH*2-1+0:0] tmp00_72_9;
	wire [WIDTH*2-1+0:0] tmp00_73_0;
	wire [WIDTH*2-1+0:0] tmp00_73_1;
	wire [WIDTH*2-1+0:0] tmp00_73_2;
	wire [WIDTH*2-1+0:0] tmp00_73_3;
	wire [WIDTH*2-1+0:0] tmp00_73_4;
	wire [WIDTH*2-1+0:0] tmp00_73_5;
	wire [WIDTH*2-1+0:0] tmp00_73_6;
	wire [WIDTH*2-1+0:0] tmp00_73_7;
	wire [WIDTH*2-1+0:0] tmp00_73_8;
	wire [WIDTH*2-1+0:0] tmp00_73_9;
	wire [WIDTH*2-1+0:0] tmp00_74_0;
	wire [WIDTH*2-1+0:0] tmp00_74_1;
	wire [WIDTH*2-1+0:0] tmp00_74_2;
	wire [WIDTH*2-1+0:0] tmp00_74_3;
	wire [WIDTH*2-1+0:0] tmp00_74_4;
	wire [WIDTH*2-1+0:0] tmp00_74_5;
	wire [WIDTH*2-1+0:0] tmp00_74_6;
	wire [WIDTH*2-1+0:0] tmp00_74_7;
	wire [WIDTH*2-1+0:0] tmp00_74_8;
	wire [WIDTH*2-1+0:0] tmp00_74_9;
	wire [WIDTH*2-1+0:0] tmp00_75_0;
	wire [WIDTH*2-1+0:0] tmp00_75_1;
	wire [WIDTH*2-1+0:0] tmp00_75_2;
	wire [WIDTH*2-1+0:0] tmp00_75_3;
	wire [WIDTH*2-1+0:0] tmp00_75_4;
	wire [WIDTH*2-1+0:0] tmp00_75_5;
	wire [WIDTH*2-1+0:0] tmp00_75_6;
	wire [WIDTH*2-1+0:0] tmp00_75_7;
	wire [WIDTH*2-1+0:0] tmp00_75_8;
	wire [WIDTH*2-1+0:0] tmp00_75_9;
	wire [WIDTH*2-1+0:0] tmp00_76_0;
	wire [WIDTH*2-1+0:0] tmp00_76_1;
	wire [WIDTH*2-1+0:0] tmp00_76_2;
	wire [WIDTH*2-1+0:0] tmp00_76_3;
	wire [WIDTH*2-1+0:0] tmp00_76_4;
	wire [WIDTH*2-1+0:0] tmp00_76_5;
	wire [WIDTH*2-1+0:0] tmp00_76_6;
	wire [WIDTH*2-1+0:0] tmp00_76_7;
	wire [WIDTH*2-1+0:0] tmp00_76_8;
	wire [WIDTH*2-1+0:0] tmp00_76_9;
	wire [WIDTH*2-1+0:0] tmp00_77_0;
	wire [WIDTH*2-1+0:0] tmp00_77_1;
	wire [WIDTH*2-1+0:0] tmp00_77_2;
	wire [WIDTH*2-1+0:0] tmp00_77_3;
	wire [WIDTH*2-1+0:0] tmp00_77_4;
	wire [WIDTH*2-1+0:0] tmp00_77_5;
	wire [WIDTH*2-1+0:0] tmp00_77_6;
	wire [WIDTH*2-1+0:0] tmp00_77_7;
	wire [WIDTH*2-1+0:0] tmp00_77_8;
	wire [WIDTH*2-1+0:0] tmp00_77_9;
	wire [WIDTH*2-1+0:0] tmp00_78_0;
	wire [WIDTH*2-1+0:0] tmp00_78_1;
	wire [WIDTH*2-1+0:0] tmp00_78_2;
	wire [WIDTH*2-1+0:0] tmp00_78_3;
	wire [WIDTH*2-1+0:0] tmp00_78_4;
	wire [WIDTH*2-1+0:0] tmp00_78_5;
	wire [WIDTH*2-1+0:0] tmp00_78_6;
	wire [WIDTH*2-1+0:0] tmp00_78_7;
	wire [WIDTH*2-1+0:0] tmp00_78_8;
	wire [WIDTH*2-1+0:0] tmp00_78_9;
	wire [WIDTH*2-1+0:0] tmp00_79_0;
	wire [WIDTH*2-1+0:0] tmp00_79_1;
	wire [WIDTH*2-1+0:0] tmp00_79_2;
	wire [WIDTH*2-1+0:0] tmp00_79_3;
	wire [WIDTH*2-1+0:0] tmp00_79_4;
	wire [WIDTH*2-1+0:0] tmp00_79_5;
	wire [WIDTH*2-1+0:0] tmp00_79_6;
	wire [WIDTH*2-1+0:0] tmp00_79_7;
	wire [WIDTH*2-1+0:0] tmp00_79_8;
	wire [WIDTH*2-1+0:0] tmp00_79_9;
	wire [WIDTH*2-1+0:0] tmp00_80_0;
	wire [WIDTH*2-1+0:0] tmp00_80_1;
	wire [WIDTH*2-1+0:0] tmp00_80_2;
	wire [WIDTH*2-1+0:0] tmp00_80_3;
	wire [WIDTH*2-1+0:0] tmp00_80_4;
	wire [WIDTH*2-1+0:0] tmp00_80_5;
	wire [WIDTH*2-1+0:0] tmp00_80_6;
	wire [WIDTH*2-1+0:0] tmp00_80_7;
	wire [WIDTH*2-1+0:0] tmp00_80_8;
	wire [WIDTH*2-1+0:0] tmp00_80_9;
	wire [WIDTH*2-1+0:0] tmp00_81_0;
	wire [WIDTH*2-1+0:0] tmp00_81_1;
	wire [WIDTH*2-1+0:0] tmp00_81_2;
	wire [WIDTH*2-1+0:0] tmp00_81_3;
	wire [WIDTH*2-1+0:0] tmp00_81_4;
	wire [WIDTH*2-1+0:0] tmp00_81_5;
	wire [WIDTH*2-1+0:0] tmp00_81_6;
	wire [WIDTH*2-1+0:0] tmp00_81_7;
	wire [WIDTH*2-1+0:0] tmp00_81_8;
	wire [WIDTH*2-1+0:0] tmp00_81_9;
	wire [WIDTH*2-1+0:0] tmp00_82_0;
	wire [WIDTH*2-1+0:0] tmp00_82_1;
	wire [WIDTH*2-1+0:0] tmp00_82_2;
	wire [WIDTH*2-1+0:0] tmp00_82_3;
	wire [WIDTH*2-1+0:0] tmp00_82_4;
	wire [WIDTH*2-1+0:0] tmp00_82_5;
	wire [WIDTH*2-1+0:0] tmp00_82_6;
	wire [WIDTH*2-1+0:0] tmp00_82_7;
	wire [WIDTH*2-1+0:0] tmp00_82_8;
	wire [WIDTH*2-1+0:0] tmp00_82_9;
	wire [WIDTH*2-1+0:0] tmp00_83_0;
	wire [WIDTH*2-1+0:0] tmp00_83_1;
	wire [WIDTH*2-1+0:0] tmp00_83_2;
	wire [WIDTH*2-1+0:0] tmp00_83_3;
	wire [WIDTH*2-1+0:0] tmp00_83_4;
	wire [WIDTH*2-1+0:0] tmp00_83_5;
	wire [WIDTH*2-1+0:0] tmp00_83_6;
	wire [WIDTH*2-1+0:0] tmp00_83_7;
	wire [WIDTH*2-1+0:0] tmp00_83_8;
	wire [WIDTH*2-1+0:0] tmp00_83_9;
	wire [WIDTH*2-1+1:0] tmp01_0_0;
	wire [WIDTH*2-1+1:0] tmp01_0_1;
	wire [WIDTH*2-1+1:0] tmp01_0_2;
	wire [WIDTH*2-1+1:0] tmp01_0_3;
	wire [WIDTH*2-1+1:0] tmp01_0_4;
	wire [WIDTH*2-1+1:0] tmp01_0_5;
	wire [WIDTH*2-1+1:0] tmp01_0_6;
	wire [WIDTH*2-1+1:0] tmp01_0_7;
	wire [WIDTH*2-1+1:0] tmp01_0_8;
	wire [WIDTH*2-1+1:0] tmp01_0_9;
	wire [WIDTH*2-1+1:0] tmp01_1_0;
	wire [WIDTH*2-1+1:0] tmp01_1_1;
	wire [WIDTH*2-1+1:0] tmp01_1_2;
	wire [WIDTH*2-1+1:0] tmp01_1_3;
	wire [WIDTH*2-1+1:0] tmp01_1_4;
	wire [WIDTH*2-1+1:0] tmp01_1_5;
	wire [WIDTH*2-1+1:0] tmp01_1_6;
	wire [WIDTH*2-1+1:0] tmp01_1_7;
	wire [WIDTH*2-1+1:0] tmp01_1_8;
	wire [WIDTH*2-1+1:0] tmp01_1_9;
	wire [WIDTH*2-1+1:0] tmp01_2_0;
	wire [WIDTH*2-1+1:0] tmp01_2_1;
	wire [WIDTH*2-1+1:0] tmp01_2_2;
	wire [WIDTH*2-1+1:0] tmp01_2_3;
	wire [WIDTH*2-1+1:0] tmp01_2_4;
	wire [WIDTH*2-1+1:0] tmp01_2_5;
	wire [WIDTH*2-1+1:0] tmp01_2_6;
	wire [WIDTH*2-1+1:0] tmp01_2_7;
	wire [WIDTH*2-1+1:0] tmp01_2_8;
	wire [WIDTH*2-1+1:0] tmp01_2_9;
	wire [WIDTH*2-1+1:0] tmp01_3_0;
	wire [WIDTH*2-1+1:0] tmp01_3_1;
	wire [WIDTH*2-1+1:0] tmp01_3_2;
	wire [WIDTH*2-1+1:0] tmp01_3_3;
	wire [WIDTH*2-1+1:0] tmp01_3_4;
	wire [WIDTH*2-1+1:0] tmp01_3_5;
	wire [WIDTH*2-1+1:0] tmp01_3_6;
	wire [WIDTH*2-1+1:0] tmp01_3_7;
	wire [WIDTH*2-1+1:0] tmp01_3_8;
	wire [WIDTH*2-1+1:0] tmp01_3_9;
	wire [WIDTH*2-1+1:0] tmp01_4_0;
	wire [WIDTH*2-1+1:0] tmp01_4_1;
	wire [WIDTH*2-1+1:0] tmp01_4_2;
	wire [WIDTH*2-1+1:0] tmp01_4_3;
	wire [WIDTH*2-1+1:0] tmp01_4_4;
	wire [WIDTH*2-1+1:0] tmp01_4_5;
	wire [WIDTH*2-1+1:0] tmp01_4_6;
	wire [WIDTH*2-1+1:0] tmp01_4_7;
	wire [WIDTH*2-1+1:0] tmp01_4_8;
	wire [WIDTH*2-1+1:0] tmp01_4_9;
	wire [WIDTH*2-1+1:0] tmp01_5_0;
	wire [WIDTH*2-1+1:0] tmp01_5_1;
	wire [WIDTH*2-1+1:0] tmp01_5_2;
	wire [WIDTH*2-1+1:0] tmp01_5_3;
	wire [WIDTH*2-1+1:0] tmp01_5_4;
	wire [WIDTH*2-1+1:0] tmp01_5_5;
	wire [WIDTH*2-1+1:0] tmp01_5_6;
	wire [WIDTH*2-1+1:0] tmp01_5_7;
	wire [WIDTH*2-1+1:0] tmp01_5_8;
	wire [WIDTH*2-1+1:0] tmp01_5_9;
	wire [WIDTH*2-1+1:0] tmp01_6_0;
	wire [WIDTH*2-1+1:0] tmp01_6_1;
	wire [WIDTH*2-1+1:0] tmp01_6_2;
	wire [WIDTH*2-1+1:0] tmp01_6_3;
	wire [WIDTH*2-1+1:0] tmp01_6_4;
	wire [WIDTH*2-1+1:0] tmp01_6_5;
	wire [WIDTH*2-1+1:0] tmp01_6_6;
	wire [WIDTH*2-1+1:0] tmp01_6_7;
	wire [WIDTH*2-1+1:0] tmp01_6_8;
	wire [WIDTH*2-1+1:0] tmp01_6_9;
	wire [WIDTH*2-1+1:0] tmp01_7_0;
	wire [WIDTH*2-1+1:0] tmp01_7_1;
	wire [WIDTH*2-1+1:0] tmp01_7_2;
	wire [WIDTH*2-1+1:0] tmp01_7_3;
	wire [WIDTH*2-1+1:0] tmp01_7_4;
	wire [WIDTH*2-1+1:0] tmp01_7_5;
	wire [WIDTH*2-1+1:0] tmp01_7_6;
	wire [WIDTH*2-1+1:0] tmp01_7_7;
	wire [WIDTH*2-1+1:0] tmp01_7_8;
	wire [WIDTH*2-1+1:0] tmp01_7_9;
	wire [WIDTH*2-1+1:0] tmp01_8_0;
	wire [WIDTH*2-1+1:0] tmp01_8_1;
	wire [WIDTH*2-1+1:0] tmp01_8_2;
	wire [WIDTH*2-1+1:0] tmp01_8_3;
	wire [WIDTH*2-1+1:0] tmp01_8_4;
	wire [WIDTH*2-1+1:0] tmp01_8_5;
	wire [WIDTH*2-1+1:0] tmp01_8_6;
	wire [WIDTH*2-1+1:0] tmp01_8_7;
	wire [WIDTH*2-1+1:0] tmp01_8_8;
	wire [WIDTH*2-1+1:0] tmp01_8_9;
	wire [WIDTH*2-1+1:0] tmp01_9_0;
	wire [WIDTH*2-1+1:0] tmp01_9_1;
	wire [WIDTH*2-1+1:0] tmp01_9_2;
	wire [WIDTH*2-1+1:0] tmp01_9_3;
	wire [WIDTH*2-1+1:0] tmp01_9_4;
	wire [WIDTH*2-1+1:0] tmp01_9_5;
	wire [WIDTH*2-1+1:0] tmp01_9_6;
	wire [WIDTH*2-1+1:0] tmp01_9_7;
	wire [WIDTH*2-1+1:0] tmp01_9_8;
	wire [WIDTH*2-1+1:0] tmp01_9_9;
	wire [WIDTH*2-1+1:0] tmp01_10_0;
	wire [WIDTH*2-1+1:0] tmp01_10_1;
	wire [WIDTH*2-1+1:0] tmp01_10_2;
	wire [WIDTH*2-1+1:0] tmp01_10_3;
	wire [WIDTH*2-1+1:0] tmp01_10_4;
	wire [WIDTH*2-1+1:0] tmp01_10_5;
	wire [WIDTH*2-1+1:0] tmp01_10_6;
	wire [WIDTH*2-1+1:0] tmp01_10_7;
	wire [WIDTH*2-1+1:0] tmp01_10_8;
	wire [WIDTH*2-1+1:0] tmp01_10_9;
	wire [WIDTH*2-1+1:0] tmp01_11_0;
	wire [WIDTH*2-1+1:0] tmp01_11_1;
	wire [WIDTH*2-1+1:0] tmp01_11_2;
	wire [WIDTH*2-1+1:0] tmp01_11_3;
	wire [WIDTH*2-1+1:0] tmp01_11_4;
	wire [WIDTH*2-1+1:0] tmp01_11_5;
	wire [WIDTH*2-1+1:0] tmp01_11_6;
	wire [WIDTH*2-1+1:0] tmp01_11_7;
	wire [WIDTH*2-1+1:0] tmp01_11_8;
	wire [WIDTH*2-1+1:0] tmp01_11_9;
	wire [WIDTH*2-1+1:0] tmp01_12_0;
	wire [WIDTH*2-1+1:0] tmp01_12_1;
	wire [WIDTH*2-1+1:0] tmp01_12_2;
	wire [WIDTH*2-1+1:0] tmp01_12_3;
	wire [WIDTH*2-1+1:0] tmp01_12_4;
	wire [WIDTH*2-1+1:0] tmp01_12_5;
	wire [WIDTH*2-1+1:0] tmp01_12_6;
	wire [WIDTH*2-1+1:0] tmp01_12_7;
	wire [WIDTH*2-1+1:0] tmp01_12_8;
	wire [WIDTH*2-1+1:0] tmp01_12_9;
	wire [WIDTH*2-1+1:0] tmp01_13_0;
	wire [WIDTH*2-1+1:0] tmp01_13_1;
	wire [WIDTH*2-1+1:0] tmp01_13_2;
	wire [WIDTH*2-1+1:0] tmp01_13_3;
	wire [WIDTH*2-1+1:0] tmp01_13_4;
	wire [WIDTH*2-1+1:0] tmp01_13_5;
	wire [WIDTH*2-1+1:0] tmp01_13_6;
	wire [WIDTH*2-1+1:0] tmp01_13_7;
	wire [WIDTH*2-1+1:0] tmp01_13_8;
	wire [WIDTH*2-1+1:0] tmp01_13_9;
	wire [WIDTH*2-1+1:0] tmp01_14_0;
	wire [WIDTH*2-1+1:0] tmp01_14_1;
	wire [WIDTH*2-1+1:0] tmp01_14_2;
	wire [WIDTH*2-1+1:0] tmp01_14_3;
	wire [WIDTH*2-1+1:0] tmp01_14_4;
	wire [WIDTH*2-1+1:0] tmp01_14_5;
	wire [WIDTH*2-1+1:0] tmp01_14_6;
	wire [WIDTH*2-1+1:0] tmp01_14_7;
	wire [WIDTH*2-1+1:0] tmp01_14_8;
	wire [WIDTH*2-1+1:0] tmp01_14_9;
	wire [WIDTH*2-1+1:0] tmp01_15_0;
	wire [WIDTH*2-1+1:0] tmp01_15_1;
	wire [WIDTH*2-1+1:0] tmp01_15_2;
	wire [WIDTH*2-1+1:0] tmp01_15_3;
	wire [WIDTH*2-1+1:0] tmp01_15_4;
	wire [WIDTH*2-1+1:0] tmp01_15_5;
	wire [WIDTH*2-1+1:0] tmp01_15_6;
	wire [WIDTH*2-1+1:0] tmp01_15_7;
	wire [WIDTH*2-1+1:0] tmp01_15_8;
	wire [WIDTH*2-1+1:0] tmp01_15_9;
	wire [WIDTH*2-1+1:0] tmp01_16_0;
	wire [WIDTH*2-1+1:0] tmp01_16_1;
	wire [WIDTH*2-1+1:0] tmp01_16_2;
	wire [WIDTH*2-1+1:0] tmp01_16_3;
	wire [WIDTH*2-1+1:0] tmp01_16_4;
	wire [WIDTH*2-1+1:0] tmp01_16_5;
	wire [WIDTH*2-1+1:0] tmp01_16_6;
	wire [WIDTH*2-1+1:0] tmp01_16_7;
	wire [WIDTH*2-1+1:0] tmp01_16_8;
	wire [WIDTH*2-1+1:0] tmp01_16_9;
	wire [WIDTH*2-1+1:0] tmp01_17_0;
	wire [WIDTH*2-1+1:0] tmp01_17_1;
	wire [WIDTH*2-1+1:0] tmp01_17_2;
	wire [WIDTH*2-1+1:0] tmp01_17_3;
	wire [WIDTH*2-1+1:0] tmp01_17_4;
	wire [WIDTH*2-1+1:0] tmp01_17_5;
	wire [WIDTH*2-1+1:0] tmp01_17_6;
	wire [WIDTH*2-1+1:0] tmp01_17_7;
	wire [WIDTH*2-1+1:0] tmp01_17_8;
	wire [WIDTH*2-1+1:0] tmp01_17_9;
	wire [WIDTH*2-1+1:0] tmp01_18_0;
	wire [WIDTH*2-1+1:0] tmp01_18_1;
	wire [WIDTH*2-1+1:0] tmp01_18_2;
	wire [WIDTH*2-1+1:0] tmp01_18_3;
	wire [WIDTH*2-1+1:0] tmp01_18_4;
	wire [WIDTH*2-1+1:0] tmp01_18_5;
	wire [WIDTH*2-1+1:0] tmp01_18_6;
	wire [WIDTH*2-1+1:0] tmp01_18_7;
	wire [WIDTH*2-1+1:0] tmp01_18_8;
	wire [WIDTH*2-1+1:0] tmp01_18_9;
	wire [WIDTH*2-1+1:0] tmp01_19_0;
	wire [WIDTH*2-1+1:0] tmp01_19_1;
	wire [WIDTH*2-1+1:0] tmp01_19_2;
	wire [WIDTH*2-1+1:0] tmp01_19_3;
	wire [WIDTH*2-1+1:0] tmp01_19_4;
	wire [WIDTH*2-1+1:0] tmp01_19_5;
	wire [WIDTH*2-1+1:0] tmp01_19_6;
	wire [WIDTH*2-1+1:0] tmp01_19_7;
	wire [WIDTH*2-1+1:0] tmp01_19_8;
	wire [WIDTH*2-1+1:0] tmp01_19_9;
	wire [WIDTH*2-1+1:0] tmp01_20_0;
	wire [WIDTH*2-1+1:0] tmp01_20_1;
	wire [WIDTH*2-1+1:0] tmp01_20_2;
	wire [WIDTH*2-1+1:0] tmp01_20_3;
	wire [WIDTH*2-1+1:0] tmp01_20_4;
	wire [WIDTH*2-1+1:0] tmp01_20_5;
	wire [WIDTH*2-1+1:0] tmp01_20_6;
	wire [WIDTH*2-1+1:0] tmp01_20_7;
	wire [WIDTH*2-1+1:0] tmp01_20_8;
	wire [WIDTH*2-1+1:0] tmp01_20_9;
	wire [WIDTH*2-1+1:0] tmp01_21_0;
	wire [WIDTH*2-1+1:0] tmp01_21_1;
	wire [WIDTH*2-1+1:0] tmp01_21_2;
	wire [WIDTH*2-1+1:0] tmp01_21_3;
	wire [WIDTH*2-1+1:0] tmp01_21_4;
	wire [WIDTH*2-1+1:0] tmp01_21_5;
	wire [WIDTH*2-1+1:0] tmp01_21_6;
	wire [WIDTH*2-1+1:0] tmp01_21_7;
	wire [WIDTH*2-1+1:0] tmp01_21_8;
	wire [WIDTH*2-1+1:0] tmp01_21_9;
	wire [WIDTH*2-1+1:0] tmp01_22_0;
	wire [WIDTH*2-1+1:0] tmp01_22_1;
	wire [WIDTH*2-1+1:0] tmp01_22_2;
	wire [WIDTH*2-1+1:0] tmp01_22_3;
	wire [WIDTH*2-1+1:0] tmp01_22_4;
	wire [WIDTH*2-1+1:0] tmp01_22_5;
	wire [WIDTH*2-1+1:0] tmp01_22_6;
	wire [WIDTH*2-1+1:0] tmp01_22_7;
	wire [WIDTH*2-1+1:0] tmp01_22_8;
	wire [WIDTH*2-1+1:0] tmp01_22_9;
	wire [WIDTH*2-1+1:0] tmp01_23_0;
	wire [WIDTH*2-1+1:0] tmp01_23_1;
	wire [WIDTH*2-1+1:0] tmp01_23_2;
	wire [WIDTH*2-1+1:0] tmp01_23_3;
	wire [WIDTH*2-1+1:0] tmp01_23_4;
	wire [WIDTH*2-1+1:0] tmp01_23_5;
	wire [WIDTH*2-1+1:0] tmp01_23_6;
	wire [WIDTH*2-1+1:0] tmp01_23_7;
	wire [WIDTH*2-1+1:0] tmp01_23_8;
	wire [WIDTH*2-1+1:0] tmp01_23_9;
	wire [WIDTH*2-1+1:0] tmp01_24_0;
	wire [WIDTH*2-1+1:0] tmp01_24_1;
	wire [WIDTH*2-1+1:0] tmp01_24_2;
	wire [WIDTH*2-1+1:0] tmp01_24_3;
	wire [WIDTH*2-1+1:0] tmp01_24_4;
	wire [WIDTH*2-1+1:0] tmp01_24_5;
	wire [WIDTH*2-1+1:0] tmp01_24_6;
	wire [WIDTH*2-1+1:0] tmp01_24_7;
	wire [WIDTH*2-1+1:0] tmp01_24_8;
	wire [WIDTH*2-1+1:0] tmp01_24_9;
	wire [WIDTH*2-1+1:0] tmp01_25_0;
	wire [WIDTH*2-1+1:0] tmp01_25_1;
	wire [WIDTH*2-1+1:0] tmp01_25_2;
	wire [WIDTH*2-1+1:0] tmp01_25_3;
	wire [WIDTH*2-1+1:0] tmp01_25_4;
	wire [WIDTH*2-1+1:0] tmp01_25_5;
	wire [WIDTH*2-1+1:0] tmp01_25_6;
	wire [WIDTH*2-1+1:0] tmp01_25_7;
	wire [WIDTH*2-1+1:0] tmp01_25_8;
	wire [WIDTH*2-1+1:0] tmp01_25_9;
	wire [WIDTH*2-1+1:0] tmp01_26_0;
	wire [WIDTH*2-1+1:0] tmp01_26_1;
	wire [WIDTH*2-1+1:0] tmp01_26_2;
	wire [WIDTH*2-1+1:0] tmp01_26_3;
	wire [WIDTH*2-1+1:0] tmp01_26_4;
	wire [WIDTH*2-1+1:0] tmp01_26_5;
	wire [WIDTH*2-1+1:0] tmp01_26_6;
	wire [WIDTH*2-1+1:0] tmp01_26_7;
	wire [WIDTH*2-1+1:0] tmp01_26_8;
	wire [WIDTH*2-1+1:0] tmp01_26_9;
	wire [WIDTH*2-1+1:0] tmp01_27_0;
	wire [WIDTH*2-1+1:0] tmp01_27_1;
	wire [WIDTH*2-1+1:0] tmp01_27_2;
	wire [WIDTH*2-1+1:0] tmp01_27_3;
	wire [WIDTH*2-1+1:0] tmp01_27_4;
	wire [WIDTH*2-1+1:0] tmp01_27_5;
	wire [WIDTH*2-1+1:0] tmp01_27_6;
	wire [WIDTH*2-1+1:0] tmp01_27_7;
	wire [WIDTH*2-1+1:0] tmp01_27_8;
	wire [WIDTH*2-1+1:0] tmp01_27_9;
	wire [WIDTH*2-1+1:0] tmp01_28_0;
	wire [WIDTH*2-1+1:0] tmp01_28_1;
	wire [WIDTH*2-1+1:0] tmp01_28_2;
	wire [WIDTH*2-1+1:0] tmp01_28_3;
	wire [WIDTH*2-1+1:0] tmp01_28_4;
	wire [WIDTH*2-1+1:0] tmp01_28_5;
	wire [WIDTH*2-1+1:0] tmp01_28_6;
	wire [WIDTH*2-1+1:0] tmp01_28_7;
	wire [WIDTH*2-1+1:0] tmp01_28_8;
	wire [WIDTH*2-1+1:0] tmp01_28_9;
	wire [WIDTH*2-1+1:0] tmp01_29_0;
	wire [WIDTH*2-1+1:0] tmp01_29_1;
	wire [WIDTH*2-1+1:0] tmp01_29_2;
	wire [WIDTH*2-1+1:0] tmp01_29_3;
	wire [WIDTH*2-1+1:0] tmp01_29_4;
	wire [WIDTH*2-1+1:0] tmp01_29_5;
	wire [WIDTH*2-1+1:0] tmp01_29_6;
	wire [WIDTH*2-1+1:0] tmp01_29_7;
	wire [WIDTH*2-1+1:0] tmp01_29_8;
	wire [WIDTH*2-1+1:0] tmp01_29_9;
	wire [WIDTH*2-1+1:0] tmp01_30_0;
	wire [WIDTH*2-1+1:0] tmp01_30_1;
	wire [WIDTH*2-1+1:0] tmp01_30_2;
	wire [WIDTH*2-1+1:0] tmp01_30_3;
	wire [WIDTH*2-1+1:0] tmp01_30_4;
	wire [WIDTH*2-1+1:0] tmp01_30_5;
	wire [WIDTH*2-1+1:0] tmp01_30_6;
	wire [WIDTH*2-1+1:0] tmp01_30_7;
	wire [WIDTH*2-1+1:0] tmp01_30_8;
	wire [WIDTH*2-1+1:0] tmp01_30_9;
	wire [WIDTH*2-1+1:0] tmp01_31_0;
	wire [WIDTH*2-1+1:0] tmp01_31_1;
	wire [WIDTH*2-1+1:0] tmp01_31_2;
	wire [WIDTH*2-1+1:0] tmp01_31_3;
	wire [WIDTH*2-1+1:0] tmp01_31_4;
	wire [WIDTH*2-1+1:0] tmp01_31_5;
	wire [WIDTH*2-1+1:0] tmp01_31_6;
	wire [WIDTH*2-1+1:0] tmp01_31_7;
	wire [WIDTH*2-1+1:0] tmp01_31_8;
	wire [WIDTH*2-1+1:0] tmp01_31_9;
	wire [WIDTH*2-1+1:0] tmp01_32_0;
	wire [WIDTH*2-1+1:0] tmp01_32_1;
	wire [WIDTH*2-1+1:0] tmp01_32_2;
	wire [WIDTH*2-1+1:0] tmp01_32_3;
	wire [WIDTH*2-1+1:0] tmp01_32_4;
	wire [WIDTH*2-1+1:0] tmp01_32_5;
	wire [WIDTH*2-1+1:0] tmp01_32_6;
	wire [WIDTH*2-1+1:0] tmp01_32_7;
	wire [WIDTH*2-1+1:0] tmp01_32_8;
	wire [WIDTH*2-1+1:0] tmp01_32_9;
	wire [WIDTH*2-1+1:0] tmp01_33_0;
	wire [WIDTH*2-1+1:0] tmp01_33_1;
	wire [WIDTH*2-1+1:0] tmp01_33_2;
	wire [WIDTH*2-1+1:0] tmp01_33_3;
	wire [WIDTH*2-1+1:0] tmp01_33_4;
	wire [WIDTH*2-1+1:0] tmp01_33_5;
	wire [WIDTH*2-1+1:0] tmp01_33_6;
	wire [WIDTH*2-1+1:0] tmp01_33_7;
	wire [WIDTH*2-1+1:0] tmp01_33_8;
	wire [WIDTH*2-1+1:0] tmp01_33_9;
	wire [WIDTH*2-1+1:0] tmp01_34_0;
	wire [WIDTH*2-1+1:0] tmp01_34_1;
	wire [WIDTH*2-1+1:0] tmp01_34_2;
	wire [WIDTH*2-1+1:0] tmp01_34_3;
	wire [WIDTH*2-1+1:0] tmp01_34_4;
	wire [WIDTH*2-1+1:0] tmp01_34_5;
	wire [WIDTH*2-1+1:0] tmp01_34_6;
	wire [WIDTH*2-1+1:0] tmp01_34_7;
	wire [WIDTH*2-1+1:0] tmp01_34_8;
	wire [WIDTH*2-1+1:0] tmp01_34_9;
	wire [WIDTH*2-1+1:0] tmp01_35_0;
	wire [WIDTH*2-1+1:0] tmp01_35_1;
	wire [WIDTH*2-1+1:0] tmp01_35_2;
	wire [WIDTH*2-1+1:0] tmp01_35_3;
	wire [WIDTH*2-1+1:0] tmp01_35_4;
	wire [WIDTH*2-1+1:0] tmp01_35_5;
	wire [WIDTH*2-1+1:0] tmp01_35_6;
	wire [WIDTH*2-1+1:0] tmp01_35_7;
	wire [WIDTH*2-1+1:0] tmp01_35_8;
	wire [WIDTH*2-1+1:0] tmp01_35_9;
	wire [WIDTH*2-1+1:0] tmp01_36_0;
	wire [WIDTH*2-1+1:0] tmp01_36_1;
	wire [WIDTH*2-1+1:0] tmp01_36_2;
	wire [WIDTH*2-1+1:0] tmp01_36_3;
	wire [WIDTH*2-1+1:0] tmp01_36_4;
	wire [WIDTH*2-1+1:0] tmp01_36_5;
	wire [WIDTH*2-1+1:0] tmp01_36_6;
	wire [WIDTH*2-1+1:0] tmp01_36_7;
	wire [WIDTH*2-1+1:0] tmp01_36_8;
	wire [WIDTH*2-1+1:0] tmp01_36_9;
	wire [WIDTH*2-1+1:0] tmp01_37_0;
	wire [WIDTH*2-1+1:0] tmp01_37_1;
	wire [WIDTH*2-1+1:0] tmp01_37_2;
	wire [WIDTH*2-1+1:0] tmp01_37_3;
	wire [WIDTH*2-1+1:0] tmp01_37_4;
	wire [WIDTH*2-1+1:0] tmp01_37_5;
	wire [WIDTH*2-1+1:0] tmp01_37_6;
	wire [WIDTH*2-1+1:0] tmp01_37_7;
	wire [WIDTH*2-1+1:0] tmp01_37_8;
	wire [WIDTH*2-1+1:0] tmp01_37_9;
	wire [WIDTH*2-1+1:0] tmp01_38_0;
	wire [WIDTH*2-1+1:0] tmp01_38_1;
	wire [WIDTH*2-1+1:0] tmp01_38_2;
	wire [WIDTH*2-1+1:0] tmp01_38_3;
	wire [WIDTH*2-1+1:0] tmp01_38_4;
	wire [WIDTH*2-1+1:0] tmp01_38_5;
	wire [WIDTH*2-1+1:0] tmp01_38_6;
	wire [WIDTH*2-1+1:0] tmp01_38_7;
	wire [WIDTH*2-1+1:0] tmp01_38_8;
	wire [WIDTH*2-1+1:0] tmp01_38_9;
	wire [WIDTH*2-1+1:0] tmp01_39_0;
	wire [WIDTH*2-1+1:0] tmp01_39_1;
	wire [WIDTH*2-1+1:0] tmp01_39_2;
	wire [WIDTH*2-1+1:0] tmp01_39_3;
	wire [WIDTH*2-1+1:0] tmp01_39_4;
	wire [WIDTH*2-1+1:0] tmp01_39_5;
	wire [WIDTH*2-1+1:0] tmp01_39_6;
	wire [WIDTH*2-1+1:0] tmp01_39_7;
	wire [WIDTH*2-1+1:0] tmp01_39_8;
	wire [WIDTH*2-1+1:0] tmp01_39_9;
	wire [WIDTH*2-1+1:0] tmp01_40_0;
	wire [WIDTH*2-1+1:0] tmp01_40_1;
	wire [WIDTH*2-1+1:0] tmp01_40_2;
	wire [WIDTH*2-1+1:0] tmp01_40_3;
	wire [WIDTH*2-1+1:0] tmp01_40_4;
	wire [WIDTH*2-1+1:0] tmp01_40_5;
	wire [WIDTH*2-1+1:0] tmp01_40_6;
	wire [WIDTH*2-1+1:0] tmp01_40_7;
	wire [WIDTH*2-1+1:0] tmp01_40_8;
	wire [WIDTH*2-1+1:0] tmp01_40_9;
	wire [WIDTH*2-1+1:0] tmp01_41_0;
	wire [WIDTH*2-1+1:0] tmp01_41_1;
	wire [WIDTH*2-1+1:0] tmp01_41_2;
	wire [WIDTH*2-1+1:0] tmp01_41_3;
	wire [WIDTH*2-1+1:0] tmp01_41_4;
	wire [WIDTH*2-1+1:0] tmp01_41_5;
	wire [WIDTH*2-1+1:0] tmp01_41_6;
	wire [WIDTH*2-1+1:0] tmp01_41_7;
	wire [WIDTH*2-1+1:0] tmp01_41_8;
	wire [WIDTH*2-1+1:0] tmp01_41_9;
	wire [WIDTH*2-1+2:0] tmp02_0_0;
	wire [WIDTH*2-1+2:0] tmp02_0_1;
	wire [WIDTH*2-1+2:0] tmp02_0_2;
	wire [WIDTH*2-1+2:0] tmp02_0_3;
	wire [WIDTH*2-1+2:0] tmp02_0_4;
	wire [WIDTH*2-1+2:0] tmp02_0_5;
	wire [WIDTH*2-1+2:0] tmp02_0_6;
	wire [WIDTH*2-1+2:0] tmp02_0_7;
	wire [WIDTH*2-1+2:0] tmp02_0_8;
	wire [WIDTH*2-1+2:0] tmp02_0_9;
	wire [WIDTH*2-1+2:0] tmp02_1_0;
	wire [WIDTH*2-1+2:0] tmp02_1_1;
	wire [WIDTH*2-1+2:0] tmp02_1_2;
	wire [WIDTH*2-1+2:0] tmp02_1_3;
	wire [WIDTH*2-1+2:0] tmp02_1_4;
	wire [WIDTH*2-1+2:0] tmp02_1_5;
	wire [WIDTH*2-1+2:0] tmp02_1_6;
	wire [WIDTH*2-1+2:0] tmp02_1_7;
	wire [WIDTH*2-1+2:0] tmp02_1_8;
	wire [WIDTH*2-1+2:0] tmp02_1_9;
	wire [WIDTH*2-1+2:0] tmp02_2_0;
	wire [WIDTH*2-1+2:0] tmp02_2_1;
	wire [WIDTH*2-1+2:0] tmp02_2_2;
	wire [WIDTH*2-1+2:0] tmp02_2_3;
	wire [WIDTH*2-1+2:0] tmp02_2_4;
	wire [WIDTH*2-1+2:0] tmp02_2_5;
	wire [WIDTH*2-1+2:0] tmp02_2_6;
	wire [WIDTH*2-1+2:0] tmp02_2_7;
	wire [WIDTH*2-1+2:0] tmp02_2_8;
	wire [WIDTH*2-1+2:0] tmp02_2_9;
	wire [WIDTH*2-1+2:0] tmp02_3_0;
	wire [WIDTH*2-1+2:0] tmp02_3_1;
	wire [WIDTH*2-1+2:0] tmp02_3_2;
	wire [WIDTH*2-1+2:0] tmp02_3_3;
	wire [WIDTH*2-1+2:0] tmp02_3_4;
	wire [WIDTH*2-1+2:0] tmp02_3_5;
	wire [WIDTH*2-1+2:0] tmp02_3_6;
	wire [WIDTH*2-1+2:0] tmp02_3_7;
	wire [WIDTH*2-1+2:0] tmp02_3_8;
	wire [WIDTH*2-1+2:0] tmp02_3_9;
	wire [WIDTH*2-1+2:0] tmp02_4_0;
	wire [WIDTH*2-1+2:0] tmp02_4_1;
	wire [WIDTH*2-1+2:0] tmp02_4_2;
	wire [WIDTH*2-1+2:0] tmp02_4_3;
	wire [WIDTH*2-1+2:0] tmp02_4_4;
	wire [WIDTH*2-1+2:0] tmp02_4_5;
	wire [WIDTH*2-1+2:0] tmp02_4_6;
	wire [WIDTH*2-1+2:0] tmp02_4_7;
	wire [WIDTH*2-1+2:0] tmp02_4_8;
	wire [WIDTH*2-1+2:0] tmp02_4_9;
	wire [WIDTH*2-1+2:0] tmp02_5_0;
	wire [WIDTH*2-1+2:0] tmp02_5_1;
	wire [WIDTH*2-1+2:0] tmp02_5_2;
	wire [WIDTH*2-1+2:0] tmp02_5_3;
	wire [WIDTH*2-1+2:0] tmp02_5_4;
	wire [WIDTH*2-1+2:0] tmp02_5_5;
	wire [WIDTH*2-1+2:0] tmp02_5_6;
	wire [WIDTH*2-1+2:0] tmp02_5_7;
	wire [WIDTH*2-1+2:0] tmp02_5_8;
	wire [WIDTH*2-1+2:0] tmp02_5_9;
	wire [WIDTH*2-1+2:0] tmp02_6_0;
	wire [WIDTH*2-1+2:0] tmp02_6_1;
	wire [WIDTH*2-1+2:0] tmp02_6_2;
	wire [WIDTH*2-1+2:0] tmp02_6_3;
	wire [WIDTH*2-1+2:0] tmp02_6_4;
	wire [WIDTH*2-1+2:0] tmp02_6_5;
	wire [WIDTH*2-1+2:0] tmp02_6_6;
	wire [WIDTH*2-1+2:0] tmp02_6_7;
	wire [WIDTH*2-1+2:0] tmp02_6_8;
	wire [WIDTH*2-1+2:0] tmp02_6_9;
	wire [WIDTH*2-1+2:0] tmp02_7_0;
	wire [WIDTH*2-1+2:0] tmp02_7_1;
	wire [WIDTH*2-1+2:0] tmp02_7_2;
	wire [WIDTH*2-1+2:0] tmp02_7_3;
	wire [WIDTH*2-1+2:0] tmp02_7_4;
	wire [WIDTH*2-1+2:0] tmp02_7_5;
	wire [WIDTH*2-1+2:0] tmp02_7_6;
	wire [WIDTH*2-1+2:0] tmp02_7_7;
	wire [WIDTH*2-1+2:0] tmp02_7_8;
	wire [WIDTH*2-1+2:0] tmp02_7_9;
	wire [WIDTH*2-1+2:0] tmp02_8_0;
	wire [WIDTH*2-1+2:0] tmp02_8_1;
	wire [WIDTH*2-1+2:0] tmp02_8_2;
	wire [WIDTH*2-1+2:0] tmp02_8_3;
	wire [WIDTH*2-1+2:0] tmp02_8_4;
	wire [WIDTH*2-1+2:0] tmp02_8_5;
	wire [WIDTH*2-1+2:0] tmp02_8_6;
	wire [WIDTH*2-1+2:0] tmp02_8_7;
	wire [WIDTH*2-1+2:0] tmp02_8_8;
	wire [WIDTH*2-1+2:0] tmp02_8_9;
	wire [WIDTH*2-1+2:0] tmp02_9_0;
	wire [WIDTH*2-1+2:0] tmp02_9_1;
	wire [WIDTH*2-1+2:0] tmp02_9_2;
	wire [WIDTH*2-1+2:0] tmp02_9_3;
	wire [WIDTH*2-1+2:0] tmp02_9_4;
	wire [WIDTH*2-1+2:0] tmp02_9_5;
	wire [WIDTH*2-1+2:0] tmp02_9_6;
	wire [WIDTH*2-1+2:0] tmp02_9_7;
	wire [WIDTH*2-1+2:0] tmp02_9_8;
	wire [WIDTH*2-1+2:0] tmp02_9_9;
	wire [WIDTH*2-1+2:0] tmp02_10_0;
	wire [WIDTH*2-1+2:0] tmp02_10_1;
	wire [WIDTH*2-1+2:0] tmp02_10_2;
	wire [WIDTH*2-1+2:0] tmp02_10_3;
	wire [WIDTH*2-1+2:0] tmp02_10_4;
	wire [WIDTH*2-1+2:0] tmp02_10_5;
	wire [WIDTH*2-1+2:0] tmp02_10_6;
	wire [WIDTH*2-1+2:0] tmp02_10_7;
	wire [WIDTH*2-1+2:0] tmp02_10_8;
	wire [WIDTH*2-1+2:0] tmp02_10_9;
	wire [WIDTH*2-1+2:0] tmp02_11_0;
	wire [WIDTH*2-1+2:0] tmp02_11_1;
	wire [WIDTH*2-1+2:0] tmp02_11_2;
	wire [WIDTH*2-1+2:0] tmp02_11_3;
	wire [WIDTH*2-1+2:0] tmp02_11_4;
	wire [WIDTH*2-1+2:0] tmp02_11_5;
	wire [WIDTH*2-1+2:0] tmp02_11_6;
	wire [WIDTH*2-1+2:0] tmp02_11_7;
	wire [WIDTH*2-1+2:0] tmp02_11_8;
	wire [WIDTH*2-1+2:0] tmp02_11_9;
	wire [WIDTH*2-1+2:0] tmp02_12_0;
	wire [WIDTH*2-1+2:0] tmp02_12_1;
	wire [WIDTH*2-1+2:0] tmp02_12_2;
	wire [WIDTH*2-1+2:0] tmp02_12_3;
	wire [WIDTH*2-1+2:0] tmp02_12_4;
	wire [WIDTH*2-1+2:0] tmp02_12_5;
	wire [WIDTH*2-1+2:0] tmp02_12_6;
	wire [WIDTH*2-1+2:0] tmp02_12_7;
	wire [WIDTH*2-1+2:0] tmp02_12_8;
	wire [WIDTH*2-1+2:0] tmp02_12_9;
	wire [WIDTH*2-1+2:0] tmp02_13_0;
	wire [WIDTH*2-1+2:0] tmp02_13_1;
	wire [WIDTH*2-1+2:0] tmp02_13_2;
	wire [WIDTH*2-1+2:0] tmp02_13_3;
	wire [WIDTH*2-1+2:0] tmp02_13_4;
	wire [WIDTH*2-1+2:0] tmp02_13_5;
	wire [WIDTH*2-1+2:0] tmp02_13_6;
	wire [WIDTH*2-1+2:0] tmp02_13_7;
	wire [WIDTH*2-1+2:0] tmp02_13_8;
	wire [WIDTH*2-1+2:0] tmp02_13_9;
	wire [WIDTH*2-1+2:0] tmp02_14_0;
	wire [WIDTH*2-1+2:0] tmp02_14_1;
	wire [WIDTH*2-1+2:0] tmp02_14_2;
	wire [WIDTH*2-1+2:0] tmp02_14_3;
	wire [WIDTH*2-1+2:0] tmp02_14_4;
	wire [WIDTH*2-1+2:0] tmp02_14_5;
	wire [WIDTH*2-1+2:0] tmp02_14_6;
	wire [WIDTH*2-1+2:0] tmp02_14_7;
	wire [WIDTH*2-1+2:0] tmp02_14_8;
	wire [WIDTH*2-1+2:0] tmp02_14_9;
	wire [WIDTH*2-1+2:0] tmp02_15_0;
	wire [WIDTH*2-1+2:0] tmp02_15_1;
	wire [WIDTH*2-1+2:0] tmp02_15_2;
	wire [WIDTH*2-1+2:0] tmp02_15_3;
	wire [WIDTH*2-1+2:0] tmp02_15_4;
	wire [WIDTH*2-1+2:0] tmp02_15_5;
	wire [WIDTH*2-1+2:0] tmp02_15_6;
	wire [WIDTH*2-1+2:0] tmp02_15_7;
	wire [WIDTH*2-1+2:0] tmp02_15_8;
	wire [WIDTH*2-1+2:0] tmp02_15_9;
	wire [WIDTH*2-1+2:0] tmp02_16_0;
	wire [WIDTH*2-1+2:0] tmp02_16_1;
	wire [WIDTH*2-1+2:0] tmp02_16_2;
	wire [WIDTH*2-1+2:0] tmp02_16_3;
	wire [WIDTH*2-1+2:0] tmp02_16_4;
	wire [WIDTH*2-1+2:0] tmp02_16_5;
	wire [WIDTH*2-1+2:0] tmp02_16_6;
	wire [WIDTH*2-1+2:0] tmp02_16_7;
	wire [WIDTH*2-1+2:0] tmp02_16_8;
	wire [WIDTH*2-1+2:0] tmp02_16_9;
	wire [WIDTH*2-1+2:0] tmp02_17_0;
	wire [WIDTH*2-1+2:0] tmp02_17_1;
	wire [WIDTH*2-1+2:0] tmp02_17_2;
	wire [WIDTH*2-1+2:0] tmp02_17_3;
	wire [WIDTH*2-1+2:0] tmp02_17_4;
	wire [WIDTH*2-1+2:0] tmp02_17_5;
	wire [WIDTH*2-1+2:0] tmp02_17_6;
	wire [WIDTH*2-1+2:0] tmp02_17_7;
	wire [WIDTH*2-1+2:0] tmp02_17_8;
	wire [WIDTH*2-1+2:0] tmp02_17_9;
	wire [WIDTH*2-1+2:0] tmp02_18_0;
	wire [WIDTH*2-1+2:0] tmp02_18_1;
	wire [WIDTH*2-1+2:0] tmp02_18_2;
	wire [WIDTH*2-1+2:0] tmp02_18_3;
	wire [WIDTH*2-1+2:0] tmp02_18_4;
	wire [WIDTH*2-1+2:0] tmp02_18_5;
	wire [WIDTH*2-1+2:0] tmp02_18_6;
	wire [WIDTH*2-1+2:0] tmp02_18_7;
	wire [WIDTH*2-1+2:0] tmp02_18_8;
	wire [WIDTH*2-1+2:0] tmp02_18_9;
	wire [WIDTH*2-1+2:0] tmp02_19_0;
	wire [WIDTH*2-1+2:0] tmp02_19_1;
	wire [WIDTH*2-1+2:0] tmp02_19_2;
	wire [WIDTH*2-1+2:0] tmp02_19_3;
	wire [WIDTH*2-1+2:0] tmp02_19_4;
	wire [WIDTH*2-1+2:0] tmp02_19_5;
	wire [WIDTH*2-1+2:0] tmp02_19_6;
	wire [WIDTH*2-1+2:0] tmp02_19_7;
	wire [WIDTH*2-1+2:0] tmp02_19_8;
	wire [WIDTH*2-1+2:0] tmp02_19_9;
	wire [WIDTH*2-1+2:0] tmp02_20_0;
	wire [WIDTH*2-1+2:0] tmp02_20_1;
	wire [WIDTH*2-1+2:0] tmp02_20_2;
	wire [WIDTH*2-1+2:0] tmp02_20_3;
	wire [WIDTH*2-1+2:0] tmp02_20_4;
	wire [WIDTH*2-1+2:0] tmp02_20_5;
	wire [WIDTH*2-1+2:0] tmp02_20_6;
	wire [WIDTH*2-1+2:0] tmp02_20_7;
	wire [WIDTH*2-1+2:0] tmp02_20_8;
	wire [WIDTH*2-1+2:0] tmp02_20_9;
	wire [WIDTH*2-1+3:0] tmp03_0_0;
	wire [WIDTH*2-1+3:0] tmp03_0_1;
	wire [WIDTH*2-1+3:0] tmp03_0_2;
	wire [WIDTH*2-1+3:0] tmp03_0_3;
	wire [WIDTH*2-1+3:0] tmp03_0_4;
	wire [WIDTH*2-1+3:0] tmp03_0_5;
	wire [WIDTH*2-1+3:0] tmp03_0_6;
	wire [WIDTH*2-1+3:0] tmp03_0_7;
	wire [WIDTH*2-1+3:0] tmp03_0_8;
	wire [WIDTH*2-1+3:0] tmp03_0_9;
	wire [WIDTH*2-1+3:0] tmp03_1_0;
	wire [WIDTH*2-1+3:0] tmp03_1_1;
	wire [WIDTH*2-1+3:0] tmp03_1_2;
	wire [WIDTH*2-1+3:0] tmp03_1_3;
	wire [WIDTH*2-1+3:0] tmp03_1_4;
	wire [WIDTH*2-1+3:0] tmp03_1_5;
	wire [WIDTH*2-1+3:0] tmp03_1_6;
	wire [WIDTH*2-1+3:0] tmp03_1_7;
	wire [WIDTH*2-1+3:0] tmp03_1_8;
	wire [WIDTH*2-1+3:0] tmp03_1_9;
	wire [WIDTH*2-1+3:0] tmp03_2_0;
	wire [WIDTH*2-1+3:0] tmp03_2_1;
	wire [WIDTH*2-1+3:0] tmp03_2_2;
	wire [WIDTH*2-1+3:0] tmp03_2_3;
	wire [WIDTH*2-1+3:0] tmp03_2_4;
	wire [WIDTH*2-1+3:0] tmp03_2_5;
	wire [WIDTH*2-1+3:0] tmp03_2_6;
	wire [WIDTH*2-1+3:0] tmp03_2_7;
	wire [WIDTH*2-1+3:0] tmp03_2_8;
	wire [WIDTH*2-1+3:0] tmp03_2_9;
	wire [WIDTH*2-1+3:0] tmp03_3_0;
	wire [WIDTH*2-1+3:0] tmp03_3_1;
	wire [WIDTH*2-1+3:0] tmp03_3_2;
	wire [WIDTH*2-1+3:0] tmp03_3_3;
	wire [WIDTH*2-1+3:0] tmp03_3_4;
	wire [WIDTH*2-1+3:0] tmp03_3_5;
	wire [WIDTH*2-1+3:0] tmp03_3_6;
	wire [WIDTH*2-1+3:0] tmp03_3_7;
	wire [WIDTH*2-1+3:0] tmp03_3_8;
	wire [WIDTH*2-1+3:0] tmp03_3_9;
	wire [WIDTH*2-1+3:0] tmp03_4_0;
	wire [WIDTH*2-1+3:0] tmp03_4_1;
	wire [WIDTH*2-1+3:0] tmp03_4_2;
	wire [WIDTH*2-1+3:0] tmp03_4_3;
	wire [WIDTH*2-1+3:0] tmp03_4_4;
	wire [WIDTH*2-1+3:0] tmp03_4_5;
	wire [WIDTH*2-1+3:0] tmp03_4_6;
	wire [WIDTH*2-1+3:0] tmp03_4_7;
	wire [WIDTH*2-1+3:0] tmp03_4_8;
	wire [WIDTH*2-1+3:0] tmp03_4_9;
	wire [WIDTH*2-1+3:0] tmp03_5_0;
	wire [WIDTH*2-1+3:0] tmp03_5_1;
	wire [WIDTH*2-1+3:0] tmp03_5_2;
	wire [WIDTH*2-1+3:0] tmp03_5_3;
	wire [WIDTH*2-1+3:0] tmp03_5_4;
	wire [WIDTH*2-1+3:0] tmp03_5_5;
	wire [WIDTH*2-1+3:0] tmp03_5_6;
	wire [WIDTH*2-1+3:0] tmp03_5_7;
	wire [WIDTH*2-1+3:0] tmp03_5_8;
	wire [WIDTH*2-1+3:0] tmp03_5_9;
	wire [WIDTH*2-1+3:0] tmp03_6_0;
	wire [WIDTH*2-1+3:0] tmp03_6_1;
	wire [WIDTH*2-1+3:0] tmp03_6_2;
	wire [WIDTH*2-1+3:0] tmp03_6_3;
	wire [WIDTH*2-1+3:0] tmp03_6_4;
	wire [WIDTH*2-1+3:0] tmp03_6_5;
	wire [WIDTH*2-1+3:0] tmp03_6_6;
	wire [WIDTH*2-1+3:0] tmp03_6_7;
	wire [WIDTH*2-1+3:0] tmp03_6_8;
	wire [WIDTH*2-1+3:0] tmp03_6_9;
	wire [WIDTH*2-1+3:0] tmp03_7_0;
	wire [WIDTH*2-1+3:0] tmp03_7_1;
	wire [WIDTH*2-1+3:0] tmp03_7_2;
	wire [WIDTH*2-1+3:0] tmp03_7_3;
	wire [WIDTH*2-1+3:0] tmp03_7_4;
	wire [WIDTH*2-1+3:0] tmp03_7_5;
	wire [WIDTH*2-1+3:0] tmp03_7_6;
	wire [WIDTH*2-1+3:0] tmp03_7_7;
	wire [WIDTH*2-1+3:0] tmp03_7_8;
	wire [WIDTH*2-1+3:0] tmp03_7_9;
	wire [WIDTH*2-1+3:0] tmp03_8_0;
	wire [WIDTH*2-1+3:0] tmp03_8_1;
	wire [WIDTH*2-1+3:0] tmp03_8_2;
	wire [WIDTH*2-1+3:0] tmp03_8_3;
	wire [WIDTH*2-1+3:0] tmp03_8_4;
	wire [WIDTH*2-1+3:0] tmp03_8_5;
	wire [WIDTH*2-1+3:0] tmp03_8_6;
	wire [WIDTH*2-1+3:0] tmp03_8_7;
	wire [WIDTH*2-1+3:0] tmp03_8_8;
	wire [WIDTH*2-1+3:0] tmp03_8_9;
	wire [WIDTH*2-1+3:0] tmp03_9_0;
	wire [WIDTH*2-1+3:0] tmp03_9_1;
	wire [WIDTH*2-1+3:0] tmp03_9_2;
	wire [WIDTH*2-1+3:0] tmp03_9_3;
	wire [WIDTH*2-1+3:0] tmp03_9_4;
	wire [WIDTH*2-1+3:0] tmp03_9_5;
	wire [WIDTH*2-1+3:0] tmp03_9_6;
	wire [WIDTH*2-1+3:0] tmp03_9_7;
	wire [WIDTH*2-1+3:0] tmp03_9_8;
	wire [WIDTH*2-1+3:0] tmp03_9_9;
	wire [WIDTH*2-1+3:0] tmp03_10_0;
	wire [WIDTH*2-1+3:0] tmp03_10_1;
	wire [WIDTH*2-1+3:0] tmp03_10_2;
	wire [WIDTH*2-1+3:0] tmp03_10_3;
	wire [WIDTH*2-1+3:0] tmp03_10_4;
	wire [WIDTH*2-1+3:0] tmp03_10_5;
	wire [WIDTH*2-1+3:0] tmp03_10_6;
	wire [WIDTH*2-1+3:0] tmp03_10_7;
	wire [WIDTH*2-1+3:0] tmp03_10_8;
	wire [WIDTH*2-1+3:0] tmp03_10_9;
	wire [WIDTH*2-1+4:0] tmp04_0_0;
	wire [WIDTH*2-1+4:0] tmp04_0_1;
	wire [WIDTH*2-1+4:0] tmp04_0_2;
	wire [WIDTH*2-1+4:0] tmp04_0_3;
	wire [WIDTH*2-1+4:0] tmp04_0_4;
	wire [WIDTH*2-1+4:0] tmp04_0_5;
	wire [WIDTH*2-1+4:0] tmp04_0_6;
	wire [WIDTH*2-1+4:0] tmp04_0_7;
	wire [WIDTH*2-1+4:0] tmp04_0_8;
	wire [WIDTH*2-1+4:0] tmp04_0_9;
	wire [WIDTH*2-1+4:0] tmp04_1_0;
	wire [WIDTH*2-1+4:0] tmp04_1_1;
	wire [WIDTH*2-1+4:0] tmp04_1_2;
	wire [WIDTH*2-1+4:0] tmp04_1_3;
	wire [WIDTH*2-1+4:0] tmp04_1_4;
	wire [WIDTH*2-1+4:0] tmp04_1_5;
	wire [WIDTH*2-1+4:0] tmp04_1_6;
	wire [WIDTH*2-1+4:0] tmp04_1_7;
	wire [WIDTH*2-1+4:0] tmp04_1_8;
	wire [WIDTH*2-1+4:0] tmp04_1_9;
	wire [WIDTH*2-1+4:0] tmp04_2_0;
	wire [WIDTH*2-1+4:0] tmp04_2_1;
	wire [WIDTH*2-1+4:0] tmp04_2_2;
	wire [WIDTH*2-1+4:0] tmp04_2_3;
	wire [WIDTH*2-1+4:0] tmp04_2_4;
	wire [WIDTH*2-1+4:0] tmp04_2_5;
	wire [WIDTH*2-1+4:0] tmp04_2_6;
	wire [WIDTH*2-1+4:0] tmp04_2_7;
	wire [WIDTH*2-1+4:0] tmp04_2_8;
	wire [WIDTH*2-1+4:0] tmp04_2_9;
	wire [WIDTH*2-1+4:0] tmp04_3_0;
	wire [WIDTH*2-1+4:0] tmp04_3_1;
	wire [WIDTH*2-1+4:0] tmp04_3_2;
	wire [WIDTH*2-1+4:0] tmp04_3_3;
	wire [WIDTH*2-1+4:0] tmp04_3_4;
	wire [WIDTH*2-1+4:0] tmp04_3_5;
	wire [WIDTH*2-1+4:0] tmp04_3_6;
	wire [WIDTH*2-1+4:0] tmp04_3_7;
	wire [WIDTH*2-1+4:0] tmp04_3_8;
	wire [WIDTH*2-1+4:0] tmp04_3_9;
	wire [WIDTH*2-1+4:0] tmp04_4_0;
	wire [WIDTH*2-1+4:0] tmp04_4_1;
	wire [WIDTH*2-1+4:0] tmp04_4_2;
	wire [WIDTH*2-1+4:0] tmp04_4_3;
	wire [WIDTH*2-1+4:0] tmp04_4_4;
	wire [WIDTH*2-1+4:0] tmp04_4_5;
	wire [WIDTH*2-1+4:0] tmp04_4_6;
	wire [WIDTH*2-1+4:0] tmp04_4_7;
	wire [WIDTH*2-1+4:0] tmp04_4_8;
	wire [WIDTH*2-1+4:0] tmp04_4_9;
	wire [WIDTH*2-1+4:0] tmp04_5_0;
	wire [WIDTH*2-1+4:0] tmp04_5_1;
	wire [WIDTH*2-1+4:0] tmp04_5_2;
	wire [WIDTH*2-1+4:0] tmp04_5_3;
	wire [WIDTH*2-1+4:0] tmp04_5_4;
	wire [WIDTH*2-1+4:0] tmp04_5_5;
	wire [WIDTH*2-1+4:0] tmp04_5_6;
	wire [WIDTH*2-1+4:0] tmp04_5_7;
	wire [WIDTH*2-1+4:0] tmp04_5_8;
	wire [WIDTH*2-1+4:0] tmp04_5_9;
	wire [WIDTH*2-1+5:0] tmp05_0_0;
	wire [WIDTH*2-1+5:0] tmp05_0_1;
	wire [WIDTH*2-1+5:0] tmp05_0_2;
	wire [WIDTH*2-1+5:0] tmp05_0_3;
	wire [WIDTH*2-1+5:0] tmp05_0_4;
	wire [WIDTH*2-1+5:0] tmp05_0_5;
	wire [WIDTH*2-1+5:0] tmp05_0_6;
	wire [WIDTH*2-1+5:0] tmp05_0_7;
	wire [WIDTH*2-1+5:0] tmp05_0_8;
	wire [WIDTH*2-1+5:0] tmp05_0_9;
	wire [WIDTH*2-1+5:0] tmp05_1_0;
	wire [WIDTH*2-1+5:0] tmp05_1_1;
	wire [WIDTH*2-1+5:0] tmp05_1_2;
	wire [WIDTH*2-1+5:0] tmp05_1_3;
	wire [WIDTH*2-1+5:0] tmp05_1_4;
	wire [WIDTH*2-1+5:0] tmp05_1_5;
	wire [WIDTH*2-1+5:0] tmp05_1_6;
	wire [WIDTH*2-1+5:0] tmp05_1_7;
	wire [WIDTH*2-1+5:0] tmp05_1_8;
	wire [WIDTH*2-1+5:0] tmp05_1_9;
	wire [WIDTH*2-1+5:0] tmp05_2_0;
	wire [WIDTH*2-1+5:0] tmp05_2_1;
	wire [WIDTH*2-1+5:0] tmp05_2_2;
	wire [WIDTH*2-1+5:0] tmp05_2_3;
	wire [WIDTH*2-1+5:0] tmp05_2_4;
	wire [WIDTH*2-1+5:0] tmp05_2_5;
	wire [WIDTH*2-1+5:0] tmp05_2_6;
	wire [WIDTH*2-1+5:0] tmp05_2_7;
	wire [WIDTH*2-1+5:0] tmp05_2_8;
	wire [WIDTH*2-1+5:0] tmp05_2_9;
	wire [WIDTH*2-1+6:0] tmp06_0_0;
	wire [WIDTH*2-1+6:0] tmp06_0_1;
	wire [WIDTH*2-1+6:0] tmp06_0_2;
	wire [WIDTH*2-1+6:0] tmp06_0_3;
	wire [WIDTH*2-1+6:0] tmp06_0_4;
	wire [WIDTH*2-1+6:0] tmp06_0_5;
	wire [WIDTH*2-1+6:0] tmp06_0_6;
	wire [WIDTH*2-1+6:0] tmp06_0_7;
	wire [WIDTH*2-1+6:0] tmp06_0_8;
	wire [WIDTH*2-1+6:0] tmp06_0_9;
	wire [WIDTH*2-1+6:0] tmp06_1_0;
	wire [WIDTH*2-1+6:0] tmp06_1_1;
	wire [WIDTH*2-1+6:0] tmp06_1_2;
	wire [WIDTH*2-1+6:0] tmp06_1_3;
	wire [WIDTH*2-1+6:0] tmp06_1_4;
	wire [WIDTH*2-1+6:0] tmp06_1_5;
	wire [WIDTH*2-1+6:0] tmp06_1_6;
	wire [WIDTH*2-1+6:0] tmp06_1_7;
	wire [WIDTH*2-1+6:0] tmp06_1_8;
	wire [WIDTH*2-1+6:0] tmp06_1_9;
	wire [WIDTH*2-1+7:0] tmp07_0_0;
	wire [WIDTH*2-1+7:0] tmp07_0_1;
	wire [WIDTH*2-1+7:0] tmp07_0_2;
	wire [WIDTH*2-1+7:0] tmp07_0_3;
	wire [WIDTH*2-1+7:0] tmp07_0_4;
	wire [WIDTH*2-1+7:0] tmp07_0_5;
	wire [WIDTH*2-1+7:0] tmp07_0_6;
	wire [WIDTH*2-1+7:0] tmp07_0_7;
	wire [WIDTH*2-1+7:0] tmp07_0_8;
	wire [WIDTH*2-1+7:0] tmp07_0_9;

	booth__006 #(.WIDTH(WIDTH)) mul00000000(.x(x_0), .z(tmp00_0_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000001(.x(x_1), .z(tmp00_1_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000002(.x(x_2), .z(tmp00_2_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000003(.x(x_3), .z(tmp00_3_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000004(.x(x_4), .z(tmp00_4_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000005(.x(x_5), .z(tmp00_5_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000006(.x(x_6), .z(tmp00_6_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000007(.x(x_7), .z(tmp00_7_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000008(.x(x_8), .z(tmp00_8_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000009(.x(x_9), .z(tmp00_9_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000010(.x(x_10), .z(tmp00_10_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000011(.x(x_11), .z(tmp00_11_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000012(.x(x_12), .z(tmp00_12_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000013(.x(x_13), .z(tmp00_13_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000014(.x(x_14), .z(tmp00_14_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000015(.x(x_15), .z(tmp00_15_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000016(.x(x_16), .z(tmp00_16_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000017(.x(x_17), .z(tmp00_17_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000018(.x(x_18), .z(tmp00_18_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000019(.x(x_19), .z(tmp00_19_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000020(.x(x_20), .z(tmp00_20_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000021(.x(x_21), .z(tmp00_21_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000022(.x(x_22), .z(tmp00_22_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000023(.x(x_23), .z(tmp00_23_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000024(.x(x_24), .z(tmp00_24_0));
	booth__008 #(.WIDTH(WIDTH)) mul00000025(.x(x_25), .z(tmp00_25_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000026(.x(x_26), .z(tmp00_26_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000027(.x(x_27), .z(tmp00_27_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000028(.x(x_28), .z(tmp00_28_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000029(.x(x_29), .z(tmp00_29_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000030(.x(x_30), .z(tmp00_30_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000031(.x(x_31), .z(tmp00_31_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000032(.x(x_32), .z(tmp00_32_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000033(.x(x_33), .z(tmp00_33_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000034(.x(x_34), .z(tmp00_34_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000035(.x(x_35), .z(tmp00_35_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000036(.x(x_36), .z(tmp00_36_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000037(.x(x_37), .z(tmp00_37_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000038(.x(x_38), .z(tmp00_38_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000039(.x(x_39), .z(tmp00_39_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000040(.x(x_40), .z(tmp00_40_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000041(.x(x_41), .z(tmp00_41_0));
	booth__002 #(.WIDTH(WIDTH)) mul00000042(.x(x_42), .z(tmp00_42_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000043(.x(x_43), .z(tmp00_43_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000044(.x(x_44), .z(tmp00_44_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000045(.x(x_45), .z(tmp00_45_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000046(.x(x_46), .z(tmp00_46_0));
	booth__006 #(.WIDTH(WIDTH)) mul00000047(.x(x_47), .z(tmp00_47_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000048(.x(x_48), .z(tmp00_48_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000049(.x(x_49), .z(tmp00_49_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000050(.x(x_50), .z(tmp00_50_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000051(.x(x_51), .z(tmp00_51_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000052(.x(x_52), .z(tmp00_52_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000053(.x(x_53), .z(tmp00_53_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000054(.x(x_54), .z(tmp00_54_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000055(.x(x_55), .z(tmp00_55_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000056(.x(x_56), .z(tmp00_56_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000057(.x(x_57), .z(tmp00_57_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000058(.x(x_58), .z(tmp00_58_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000059(.x(x_59), .z(tmp00_59_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000060(.x(x_60), .z(tmp00_60_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000061(.x(x_61), .z(tmp00_61_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000062(.x(x_62), .z(tmp00_62_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000063(.x(x_63), .z(tmp00_63_0));
	booth__006 #(.WIDTH(WIDTH)) mul00000064(.x(x_64), .z(tmp00_64_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000065(.x(x_65), .z(tmp00_65_0));
	booth_0006 #(.WIDTH(WIDTH)) mul00000066(.x(x_66), .z(tmp00_66_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000067(.x(x_67), .z(tmp00_67_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000068(.x(x_68), .z(tmp00_68_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000069(.x(x_69), .z(tmp00_69_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000070(.x(x_70), .z(tmp00_70_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000071(.x(x_71), .z(tmp00_71_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000072(.x(x_72), .z(tmp00_72_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000073(.x(x_73), .z(tmp00_73_0));
	booth__002 #(.WIDTH(WIDTH)) mul00000074(.x(x_74), .z(tmp00_74_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000075(.x(x_75), .z(tmp00_75_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000076(.x(x_76), .z(tmp00_76_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000077(.x(x_77), .z(tmp00_77_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000078(.x(x_78), .z(tmp00_78_0));
	booth_0004 #(.WIDTH(WIDTH)) mul00000079(.x(x_79), .z(tmp00_79_0));
	booth__004 #(.WIDTH(WIDTH)) mul00000080(.x(x_80), .z(tmp00_80_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00000081(.x(x_81), .z(tmp00_81_0));
	booth__006 #(.WIDTH(WIDTH)) mul00000082(.x(x_82), .z(tmp00_82_0));
	booth_0008 #(.WIDTH(WIDTH)) mul00000083(.x(x_83), .z(tmp00_83_0));
	booth_0000 #(.WIDTH(WIDTH)) mul00010000(.x(x_0), .z(tmp00_0_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010001(.x(x_1), .z(tmp00_1_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010002(.x(x_2), .z(tmp00_2_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010003(.x(x_3), .z(tmp00_3_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010004(.x(x_4), .z(tmp00_4_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010005(.x(x_5), .z(tmp00_5_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010006(.x(x_6), .z(tmp00_6_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010007(.x(x_7), .z(tmp00_7_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010008(.x(x_8), .z(tmp00_8_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010009(.x(x_9), .z(tmp00_9_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010010(.x(x_10), .z(tmp00_10_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010011(.x(x_11), .z(tmp00_11_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010012(.x(x_12), .z(tmp00_12_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010013(.x(x_13), .z(tmp00_13_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010014(.x(x_14), .z(tmp00_14_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010015(.x(x_15), .z(tmp00_15_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010016(.x(x_16), .z(tmp00_16_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010017(.x(x_17), .z(tmp00_17_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010018(.x(x_18), .z(tmp00_18_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010019(.x(x_19), .z(tmp00_19_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010020(.x(x_20), .z(tmp00_20_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010021(.x(x_21), .z(tmp00_21_1));
	booth__002 #(.WIDTH(WIDTH)) mul00010022(.x(x_22), .z(tmp00_22_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010023(.x(x_23), .z(tmp00_23_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010024(.x(x_24), .z(tmp00_24_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010025(.x(x_25), .z(tmp00_25_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010026(.x(x_26), .z(tmp00_26_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010027(.x(x_27), .z(tmp00_27_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010028(.x(x_28), .z(tmp00_28_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010029(.x(x_29), .z(tmp00_29_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010030(.x(x_30), .z(tmp00_30_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010031(.x(x_31), .z(tmp00_31_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010032(.x(x_32), .z(tmp00_32_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010033(.x(x_33), .z(tmp00_33_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010034(.x(x_34), .z(tmp00_34_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010035(.x(x_35), .z(tmp00_35_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010036(.x(x_36), .z(tmp00_36_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010037(.x(x_37), .z(tmp00_37_1));
	booth__008 #(.WIDTH(WIDTH)) mul00010038(.x(x_38), .z(tmp00_38_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010039(.x(x_39), .z(tmp00_39_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010040(.x(x_40), .z(tmp00_40_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010041(.x(x_41), .z(tmp00_41_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010042(.x(x_42), .z(tmp00_42_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010043(.x(x_43), .z(tmp00_43_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010044(.x(x_44), .z(tmp00_44_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010045(.x(x_45), .z(tmp00_45_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010046(.x(x_46), .z(tmp00_46_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010047(.x(x_47), .z(tmp00_47_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010048(.x(x_48), .z(tmp00_48_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010049(.x(x_49), .z(tmp00_49_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010050(.x(x_50), .z(tmp00_50_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010051(.x(x_51), .z(tmp00_51_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010052(.x(x_52), .z(tmp00_52_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010053(.x(x_53), .z(tmp00_53_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010054(.x(x_54), .z(tmp00_54_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010055(.x(x_55), .z(tmp00_55_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010056(.x(x_56), .z(tmp00_56_1));
	booth_0006 #(.WIDTH(WIDTH)) mul00010057(.x(x_57), .z(tmp00_57_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010058(.x(x_58), .z(tmp00_58_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010059(.x(x_59), .z(tmp00_59_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010060(.x(x_60), .z(tmp00_60_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010061(.x(x_61), .z(tmp00_61_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010062(.x(x_62), .z(tmp00_62_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010063(.x(x_63), .z(tmp00_63_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010064(.x(x_64), .z(tmp00_64_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010065(.x(x_65), .z(tmp00_65_1));
	booth_0004 #(.WIDTH(WIDTH)) mul00010066(.x(x_66), .z(tmp00_66_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010067(.x(x_67), .z(tmp00_67_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010068(.x(x_68), .z(tmp00_68_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010069(.x(x_69), .z(tmp00_69_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010070(.x(x_70), .z(tmp00_70_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010071(.x(x_71), .z(tmp00_71_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010072(.x(x_72), .z(tmp00_72_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010073(.x(x_73), .z(tmp00_73_1));
	booth_0008 #(.WIDTH(WIDTH)) mul00010074(.x(x_74), .z(tmp00_74_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010075(.x(x_75), .z(tmp00_75_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010076(.x(x_76), .z(tmp00_76_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010077(.x(x_77), .z(tmp00_77_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010078(.x(x_78), .z(tmp00_78_1));
	booth_0002 #(.WIDTH(WIDTH)) mul00010079(.x(x_79), .z(tmp00_79_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010080(.x(x_80), .z(tmp00_80_1));
	booth__004 #(.WIDTH(WIDTH)) mul00010081(.x(x_81), .z(tmp00_81_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010082(.x(x_82), .z(tmp00_82_1));
	booth_0000 #(.WIDTH(WIDTH)) mul00010083(.x(x_83), .z(tmp00_83_1));
	booth__006 #(.WIDTH(WIDTH)) mul00020000(.x(x_0), .z(tmp00_0_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020001(.x(x_1), .z(tmp00_1_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020002(.x(x_2), .z(tmp00_2_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020003(.x(x_3), .z(tmp00_3_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020004(.x(x_4), .z(tmp00_4_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020005(.x(x_5), .z(tmp00_5_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020006(.x(x_6), .z(tmp00_6_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020007(.x(x_7), .z(tmp00_7_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020008(.x(x_8), .z(tmp00_8_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020009(.x(x_9), .z(tmp00_9_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020010(.x(x_10), .z(tmp00_10_2));
	booth_0002 #(.WIDTH(WIDTH)) mul00020011(.x(x_11), .z(tmp00_11_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020012(.x(x_12), .z(tmp00_12_2));
	booth_0002 #(.WIDTH(WIDTH)) mul00020013(.x(x_13), .z(tmp00_13_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020014(.x(x_14), .z(tmp00_14_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020015(.x(x_15), .z(tmp00_15_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020016(.x(x_16), .z(tmp00_16_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020017(.x(x_17), .z(tmp00_17_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020018(.x(x_18), .z(tmp00_18_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020019(.x(x_19), .z(tmp00_19_2));
	booth__006 #(.WIDTH(WIDTH)) mul00020020(.x(x_20), .z(tmp00_20_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020021(.x(x_21), .z(tmp00_21_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020022(.x(x_22), .z(tmp00_22_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020023(.x(x_23), .z(tmp00_23_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020024(.x(x_24), .z(tmp00_24_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020025(.x(x_25), .z(tmp00_25_2));
	booth_0006 #(.WIDTH(WIDTH)) mul00020026(.x(x_26), .z(tmp00_26_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020027(.x(x_27), .z(tmp00_27_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020028(.x(x_28), .z(tmp00_28_2));
	booth_0006 #(.WIDTH(WIDTH)) mul00020029(.x(x_29), .z(tmp00_29_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020030(.x(x_30), .z(tmp00_30_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020031(.x(x_31), .z(tmp00_31_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020032(.x(x_32), .z(tmp00_32_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020033(.x(x_33), .z(tmp00_33_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020034(.x(x_34), .z(tmp00_34_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020035(.x(x_35), .z(tmp00_35_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020036(.x(x_36), .z(tmp00_36_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020037(.x(x_37), .z(tmp00_37_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020038(.x(x_38), .z(tmp00_38_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020039(.x(x_39), .z(tmp00_39_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020040(.x(x_40), .z(tmp00_40_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020041(.x(x_41), .z(tmp00_41_2));
	booth_0006 #(.WIDTH(WIDTH)) mul00020042(.x(x_42), .z(tmp00_42_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020043(.x(x_43), .z(tmp00_43_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020044(.x(x_44), .z(tmp00_44_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020045(.x(x_45), .z(tmp00_45_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020046(.x(x_46), .z(tmp00_46_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020047(.x(x_47), .z(tmp00_47_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020048(.x(x_48), .z(tmp00_48_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020049(.x(x_49), .z(tmp00_49_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020050(.x(x_50), .z(tmp00_50_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020051(.x(x_51), .z(tmp00_51_2));
	booth__002 #(.WIDTH(WIDTH)) mul00020052(.x(x_52), .z(tmp00_52_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020053(.x(x_53), .z(tmp00_53_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020054(.x(x_54), .z(tmp00_54_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020055(.x(x_55), .z(tmp00_55_2));
	booth_0002 #(.WIDTH(WIDTH)) mul00020056(.x(x_56), .z(tmp00_56_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020057(.x(x_57), .z(tmp00_57_2));
	booth_0002 #(.WIDTH(WIDTH)) mul00020058(.x(x_58), .z(tmp00_58_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020059(.x(x_59), .z(tmp00_59_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020060(.x(x_60), .z(tmp00_60_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020061(.x(x_61), .z(tmp00_61_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020062(.x(x_62), .z(tmp00_62_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020063(.x(x_63), .z(tmp00_63_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020064(.x(x_64), .z(tmp00_64_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00020065(.x(x_65), .z(tmp00_65_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020066(.x(x_66), .z(tmp00_66_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020067(.x(x_67), .z(tmp00_67_2));
	booth__006 #(.WIDTH(WIDTH)) mul00020068(.x(x_68), .z(tmp00_68_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020069(.x(x_69), .z(tmp00_69_2));
	booth__006 #(.WIDTH(WIDTH)) mul00020070(.x(x_70), .z(tmp00_70_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020071(.x(x_71), .z(tmp00_71_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020072(.x(x_72), .z(tmp00_72_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020073(.x(x_73), .z(tmp00_73_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020074(.x(x_74), .z(tmp00_74_2));
	booth__006 #(.WIDTH(WIDTH)) mul00020075(.x(x_75), .z(tmp00_75_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020076(.x(x_76), .z(tmp00_76_2));
	booth__006 #(.WIDTH(WIDTH)) mul00020077(.x(x_77), .z(tmp00_77_2));
	booth__004 #(.WIDTH(WIDTH)) mul00020078(.x(x_78), .z(tmp00_78_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020079(.x(x_79), .z(tmp00_79_2));
	booth__006 #(.WIDTH(WIDTH)) mul00020080(.x(x_80), .z(tmp00_80_2));
	booth_0004 #(.WIDTH(WIDTH)) mul00020081(.x(x_81), .z(tmp00_81_2));
	booth_0000 #(.WIDTH(WIDTH)) mul00020082(.x(x_82), .z(tmp00_82_2));
	booth__008 #(.WIDTH(WIDTH)) mul00020083(.x(x_83), .z(tmp00_83_2));
	booth_0008 #(.WIDTH(WIDTH)) mul00030000(.x(x_0), .z(tmp00_0_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030001(.x(x_1), .z(tmp00_1_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030002(.x(x_2), .z(tmp00_2_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030003(.x(x_3), .z(tmp00_3_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030004(.x(x_4), .z(tmp00_4_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030005(.x(x_5), .z(tmp00_5_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030006(.x(x_6), .z(tmp00_6_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030007(.x(x_7), .z(tmp00_7_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030008(.x(x_8), .z(tmp00_8_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030009(.x(x_9), .z(tmp00_9_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030010(.x(x_10), .z(tmp00_10_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030011(.x(x_11), .z(tmp00_11_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030012(.x(x_12), .z(tmp00_12_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030013(.x(x_13), .z(tmp00_13_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030014(.x(x_14), .z(tmp00_14_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030015(.x(x_15), .z(tmp00_15_3));
	booth_0002 #(.WIDTH(WIDTH)) mul00030016(.x(x_16), .z(tmp00_16_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030017(.x(x_17), .z(tmp00_17_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030018(.x(x_18), .z(tmp00_18_3));
	booth_0002 #(.WIDTH(WIDTH)) mul00030019(.x(x_19), .z(tmp00_19_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030020(.x(x_20), .z(tmp00_20_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030021(.x(x_21), .z(tmp00_21_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030022(.x(x_22), .z(tmp00_22_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030023(.x(x_23), .z(tmp00_23_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030024(.x(x_24), .z(tmp00_24_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030025(.x(x_25), .z(tmp00_25_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030026(.x(x_26), .z(tmp00_26_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030027(.x(x_27), .z(tmp00_27_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030028(.x(x_28), .z(tmp00_28_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030029(.x(x_29), .z(tmp00_29_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030030(.x(x_30), .z(tmp00_30_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030031(.x(x_31), .z(tmp00_31_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030032(.x(x_32), .z(tmp00_32_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030033(.x(x_33), .z(tmp00_33_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030034(.x(x_34), .z(tmp00_34_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030035(.x(x_35), .z(tmp00_35_3));
	booth_0002 #(.WIDTH(WIDTH)) mul00030036(.x(x_36), .z(tmp00_36_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030037(.x(x_37), .z(tmp00_37_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030038(.x(x_38), .z(tmp00_38_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030039(.x(x_39), .z(tmp00_39_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030040(.x(x_40), .z(tmp00_40_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030041(.x(x_41), .z(tmp00_41_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030042(.x(x_42), .z(tmp00_42_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030043(.x(x_43), .z(tmp00_43_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030044(.x(x_44), .z(tmp00_44_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030045(.x(x_45), .z(tmp00_45_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030046(.x(x_46), .z(tmp00_46_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030047(.x(x_47), .z(tmp00_47_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030048(.x(x_48), .z(tmp00_48_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030049(.x(x_49), .z(tmp00_49_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030050(.x(x_50), .z(tmp00_50_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030051(.x(x_51), .z(tmp00_51_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030052(.x(x_52), .z(tmp00_52_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030053(.x(x_53), .z(tmp00_53_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030054(.x(x_54), .z(tmp00_54_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030055(.x(x_55), .z(tmp00_55_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030056(.x(x_56), .z(tmp00_56_3));
	booth_0008 #(.WIDTH(WIDTH)) mul00030057(.x(x_57), .z(tmp00_57_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030058(.x(x_58), .z(tmp00_58_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030059(.x(x_59), .z(tmp00_59_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030060(.x(x_60), .z(tmp00_60_3));
	booth_0006 #(.WIDTH(WIDTH)) mul00030061(.x(x_61), .z(tmp00_61_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030062(.x(x_62), .z(tmp00_62_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030063(.x(x_63), .z(tmp00_63_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030064(.x(x_64), .z(tmp00_64_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030065(.x(x_65), .z(tmp00_65_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030066(.x(x_66), .z(tmp00_66_3));
	booth__002 #(.WIDTH(WIDTH)) mul00030067(.x(x_67), .z(tmp00_67_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030068(.x(x_68), .z(tmp00_68_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030069(.x(x_69), .z(tmp00_69_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030070(.x(x_70), .z(tmp00_70_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030071(.x(x_71), .z(tmp00_71_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030072(.x(x_72), .z(tmp00_72_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030073(.x(x_73), .z(tmp00_73_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030074(.x(x_74), .z(tmp00_74_3));
	booth__004 #(.WIDTH(WIDTH)) mul00030075(.x(x_75), .z(tmp00_75_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030076(.x(x_76), .z(tmp00_76_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030077(.x(x_77), .z(tmp00_77_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030078(.x(x_78), .z(tmp00_78_3));
	booth__006 #(.WIDTH(WIDTH)) mul00030079(.x(x_79), .z(tmp00_79_3));
	booth__008 #(.WIDTH(WIDTH)) mul00030080(.x(x_80), .z(tmp00_80_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030081(.x(x_81), .z(tmp00_81_3));
	booth_0000 #(.WIDTH(WIDTH)) mul00030082(.x(x_82), .z(tmp00_82_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00030083(.x(x_83), .z(tmp00_83_3));
	booth_0004 #(.WIDTH(WIDTH)) mul00040000(.x(x_0), .z(tmp00_0_4));
	booth_0002 #(.WIDTH(WIDTH)) mul00040001(.x(x_1), .z(tmp00_1_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040002(.x(x_2), .z(tmp00_2_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040003(.x(x_3), .z(tmp00_3_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040004(.x(x_4), .z(tmp00_4_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040005(.x(x_5), .z(tmp00_5_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040006(.x(x_6), .z(tmp00_6_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040007(.x(x_7), .z(tmp00_7_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040008(.x(x_8), .z(tmp00_8_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040009(.x(x_9), .z(tmp00_9_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040010(.x(x_10), .z(tmp00_10_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040011(.x(x_11), .z(tmp00_11_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040012(.x(x_12), .z(tmp00_12_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040013(.x(x_13), .z(tmp00_13_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040014(.x(x_14), .z(tmp00_14_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040015(.x(x_15), .z(tmp00_15_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040016(.x(x_16), .z(tmp00_16_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040017(.x(x_17), .z(tmp00_17_4));
	booth_0002 #(.WIDTH(WIDTH)) mul00040018(.x(x_18), .z(tmp00_18_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040019(.x(x_19), .z(tmp00_19_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040020(.x(x_20), .z(tmp00_20_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040021(.x(x_21), .z(tmp00_21_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040022(.x(x_22), .z(tmp00_22_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040023(.x(x_23), .z(tmp00_23_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040024(.x(x_24), .z(tmp00_24_4));
	booth_0006 #(.WIDTH(WIDTH)) mul00040025(.x(x_25), .z(tmp00_25_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040026(.x(x_26), .z(tmp00_26_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040027(.x(x_27), .z(tmp00_27_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040028(.x(x_28), .z(tmp00_28_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040029(.x(x_29), .z(tmp00_29_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040030(.x(x_30), .z(tmp00_30_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040031(.x(x_31), .z(tmp00_31_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040032(.x(x_32), .z(tmp00_32_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040033(.x(x_33), .z(tmp00_33_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040034(.x(x_34), .z(tmp00_34_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040035(.x(x_35), .z(tmp00_35_4));
	booth_0006 #(.WIDTH(WIDTH)) mul00040036(.x(x_36), .z(tmp00_36_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040037(.x(x_37), .z(tmp00_37_4));
	booth_0006 #(.WIDTH(WIDTH)) mul00040038(.x(x_38), .z(tmp00_38_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040039(.x(x_39), .z(tmp00_39_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040040(.x(x_40), .z(tmp00_40_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040041(.x(x_41), .z(tmp00_41_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040042(.x(x_42), .z(tmp00_42_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040043(.x(x_43), .z(tmp00_43_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040044(.x(x_44), .z(tmp00_44_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040045(.x(x_45), .z(tmp00_45_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040046(.x(x_46), .z(tmp00_46_4));
	booth__016 #(.WIDTH(WIDTH)) mul00040047(.x(x_47), .z(tmp00_47_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040048(.x(x_48), .z(tmp00_48_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040049(.x(x_49), .z(tmp00_49_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040050(.x(x_50), .z(tmp00_50_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040051(.x(x_51), .z(tmp00_51_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040052(.x(x_52), .z(tmp00_52_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040053(.x(x_53), .z(tmp00_53_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040054(.x(x_54), .z(tmp00_54_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040055(.x(x_55), .z(tmp00_55_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040056(.x(x_56), .z(tmp00_56_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040057(.x(x_57), .z(tmp00_57_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040058(.x(x_58), .z(tmp00_58_4));
	booth__004 #(.WIDTH(WIDTH)) mul00040059(.x(x_59), .z(tmp00_59_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040060(.x(x_60), .z(tmp00_60_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040061(.x(x_61), .z(tmp00_61_4));
	booth_0002 #(.WIDTH(WIDTH)) mul00040062(.x(x_62), .z(tmp00_62_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040063(.x(x_63), .z(tmp00_63_4));
	booth_0002 #(.WIDTH(WIDTH)) mul00040064(.x(x_64), .z(tmp00_64_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040065(.x(x_65), .z(tmp00_65_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040066(.x(x_66), .z(tmp00_66_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040067(.x(x_67), .z(tmp00_67_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040068(.x(x_68), .z(tmp00_68_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040069(.x(x_69), .z(tmp00_69_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040070(.x(x_70), .z(tmp00_70_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040071(.x(x_71), .z(tmp00_71_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040072(.x(x_72), .z(tmp00_72_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040073(.x(x_73), .z(tmp00_73_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040074(.x(x_74), .z(tmp00_74_4));
	booth__002 #(.WIDTH(WIDTH)) mul00040075(.x(x_75), .z(tmp00_75_4));
	booth__008 #(.WIDTH(WIDTH)) mul00040076(.x(x_76), .z(tmp00_76_4));
	booth_0012 #(.WIDTH(WIDTH)) mul00040077(.x(x_77), .z(tmp00_77_4));
	booth_0002 #(.WIDTH(WIDTH)) mul00040078(.x(x_78), .z(tmp00_78_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040079(.x(x_79), .z(tmp00_79_4));
	booth_0004 #(.WIDTH(WIDTH)) mul00040080(.x(x_80), .z(tmp00_80_4));
	booth_0008 #(.WIDTH(WIDTH)) mul00040081(.x(x_81), .z(tmp00_81_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040082(.x(x_82), .z(tmp00_82_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00040083(.x(x_83), .z(tmp00_83_4));
	booth_0000 #(.WIDTH(WIDTH)) mul00050000(.x(x_0), .z(tmp00_0_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050001(.x(x_1), .z(tmp00_1_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050002(.x(x_2), .z(tmp00_2_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050003(.x(x_3), .z(tmp00_3_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050004(.x(x_4), .z(tmp00_4_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050005(.x(x_5), .z(tmp00_5_5));
	booth__002 #(.WIDTH(WIDTH)) mul00050006(.x(x_6), .z(tmp00_6_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050007(.x(x_7), .z(tmp00_7_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050008(.x(x_8), .z(tmp00_8_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050009(.x(x_9), .z(tmp00_9_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050010(.x(x_10), .z(tmp00_10_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050011(.x(x_11), .z(tmp00_11_5));
	booth_0006 #(.WIDTH(WIDTH)) mul00050012(.x(x_12), .z(tmp00_12_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050013(.x(x_13), .z(tmp00_13_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050014(.x(x_14), .z(tmp00_14_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050015(.x(x_15), .z(tmp00_15_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050016(.x(x_16), .z(tmp00_16_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050017(.x(x_17), .z(tmp00_17_5));
	booth__002 #(.WIDTH(WIDTH)) mul00050018(.x(x_18), .z(tmp00_18_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050019(.x(x_19), .z(tmp00_19_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050020(.x(x_20), .z(tmp00_20_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050021(.x(x_21), .z(tmp00_21_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050022(.x(x_22), .z(tmp00_22_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050023(.x(x_23), .z(tmp00_23_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050024(.x(x_24), .z(tmp00_24_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050025(.x(x_25), .z(tmp00_25_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050026(.x(x_26), .z(tmp00_26_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050027(.x(x_27), .z(tmp00_27_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050028(.x(x_28), .z(tmp00_28_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050029(.x(x_29), .z(tmp00_29_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050030(.x(x_30), .z(tmp00_30_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050031(.x(x_31), .z(tmp00_31_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050032(.x(x_32), .z(tmp00_32_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050033(.x(x_33), .z(tmp00_33_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050034(.x(x_34), .z(tmp00_34_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050035(.x(x_35), .z(tmp00_35_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050036(.x(x_36), .z(tmp00_36_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050037(.x(x_37), .z(tmp00_37_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050038(.x(x_38), .z(tmp00_38_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050039(.x(x_39), .z(tmp00_39_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050040(.x(x_40), .z(tmp00_40_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050041(.x(x_41), .z(tmp00_41_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050042(.x(x_42), .z(tmp00_42_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050043(.x(x_43), .z(tmp00_43_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050044(.x(x_44), .z(tmp00_44_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050045(.x(x_45), .z(tmp00_45_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050046(.x(x_46), .z(tmp00_46_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050047(.x(x_47), .z(tmp00_47_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050048(.x(x_48), .z(tmp00_48_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050049(.x(x_49), .z(tmp00_49_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050050(.x(x_50), .z(tmp00_50_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050051(.x(x_51), .z(tmp00_51_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050052(.x(x_52), .z(tmp00_52_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050053(.x(x_53), .z(tmp00_53_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050054(.x(x_54), .z(tmp00_54_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050055(.x(x_55), .z(tmp00_55_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050056(.x(x_56), .z(tmp00_56_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050057(.x(x_57), .z(tmp00_57_5));
	booth_0006 #(.WIDTH(WIDTH)) mul00050058(.x(x_58), .z(tmp00_58_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050059(.x(x_59), .z(tmp00_59_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050060(.x(x_60), .z(tmp00_60_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050061(.x(x_61), .z(tmp00_61_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050062(.x(x_62), .z(tmp00_62_5));
	booth_0002 #(.WIDTH(WIDTH)) mul00050063(.x(x_63), .z(tmp00_63_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050064(.x(x_64), .z(tmp00_64_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050065(.x(x_65), .z(tmp00_65_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050066(.x(x_66), .z(tmp00_66_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050067(.x(x_67), .z(tmp00_67_5));
	booth_0008 #(.WIDTH(WIDTH)) mul00050068(.x(x_68), .z(tmp00_68_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050069(.x(x_69), .z(tmp00_69_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050070(.x(x_70), .z(tmp00_70_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050071(.x(x_71), .z(tmp00_71_5));
	booth__004 #(.WIDTH(WIDTH)) mul00050072(.x(x_72), .z(tmp00_72_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050073(.x(x_73), .z(tmp00_73_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050074(.x(x_74), .z(tmp00_74_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050075(.x(x_75), .z(tmp00_75_5));
	booth_0004 #(.WIDTH(WIDTH)) mul00050076(.x(x_76), .z(tmp00_76_5));
	booth__002 #(.WIDTH(WIDTH)) mul00050077(.x(x_77), .z(tmp00_77_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050078(.x(x_78), .z(tmp00_78_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050079(.x(x_79), .z(tmp00_79_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050080(.x(x_80), .z(tmp00_80_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050081(.x(x_81), .z(tmp00_81_5));
	booth__006 #(.WIDTH(WIDTH)) mul00050082(.x(x_82), .z(tmp00_82_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00050083(.x(x_83), .z(tmp00_83_5));
	booth_0000 #(.WIDTH(WIDTH)) mul00060000(.x(x_0), .z(tmp00_0_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060001(.x(x_1), .z(tmp00_1_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060002(.x(x_2), .z(tmp00_2_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060003(.x(x_3), .z(tmp00_3_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060004(.x(x_4), .z(tmp00_4_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060005(.x(x_5), .z(tmp00_5_6));
	booth__006 #(.WIDTH(WIDTH)) mul00060006(.x(x_6), .z(tmp00_6_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060007(.x(x_7), .z(tmp00_7_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060008(.x(x_8), .z(tmp00_8_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060009(.x(x_9), .z(tmp00_9_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060010(.x(x_10), .z(tmp00_10_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060011(.x(x_11), .z(tmp00_11_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060012(.x(x_12), .z(tmp00_12_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060013(.x(x_13), .z(tmp00_13_6));
	booth__006 #(.WIDTH(WIDTH)) mul00060014(.x(x_14), .z(tmp00_14_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060015(.x(x_15), .z(tmp00_15_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060016(.x(x_16), .z(tmp00_16_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060017(.x(x_17), .z(tmp00_17_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060018(.x(x_18), .z(tmp00_18_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060019(.x(x_19), .z(tmp00_19_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060020(.x(x_20), .z(tmp00_20_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060021(.x(x_21), .z(tmp00_21_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060022(.x(x_22), .z(tmp00_22_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060023(.x(x_23), .z(tmp00_23_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060024(.x(x_24), .z(tmp00_24_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060025(.x(x_25), .z(tmp00_25_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060026(.x(x_26), .z(tmp00_26_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060027(.x(x_27), .z(tmp00_27_6));
	booth_0008 #(.WIDTH(WIDTH)) mul00060028(.x(x_28), .z(tmp00_28_6));
	booth__002 #(.WIDTH(WIDTH)) mul00060029(.x(x_29), .z(tmp00_29_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060030(.x(x_30), .z(tmp00_30_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060031(.x(x_31), .z(tmp00_31_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060032(.x(x_32), .z(tmp00_32_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060033(.x(x_33), .z(tmp00_33_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060034(.x(x_34), .z(tmp00_34_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060035(.x(x_35), .z(tmp00_35_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060036(.x(x_36), .z(tmp00_36_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060037(.x(x_37), .z(tmp00_37_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060038(.x(x_38), .z(tmp00_38_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060039(.x(x_39), .z(tmp00_39_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060040(.x(x_40), .z(tmp00_40_6));
	booth__002 #(.WIDTH(WIDTH)) mul00060041(.x(x_41), .z(tmp00_41_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060042(.x(x_42), .z(tmp00_42_6));
	booth_0006 #(.WIDTH(WIDTH)) mul00060043(.x(x_43), .z(tmp00_43_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060044(.x(x_44), .z(tmp00_44_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060045(.x(x_45), .z(tmp00_45_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060046(.x(x_46), .z(tmp00_46_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060047(.x(x_47), .z(tmp00_47_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060048(.x(x_48), .z(tmp00_48_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060049(.x(x_49), .z(tmp00_49_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060050(.x(x_50), .z(tmp00_50_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060051(.x(x_51), .z(tmp00_51_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060052(.x(x_52), .z(tmp00_52_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060053(.x(x_53), .z(tmp00_53_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060054(.x(x_54), .z(tmp00_54_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060055(.x(x_55), .z(tmp00_55_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060056(.x(x_56), .z(tmp00_56_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060057(.x(x_57), .z(tmp00_57_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060058(.x(x_58), .z(tmp00_58_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060059(.x(x_59), .z(tmp00_59_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060060(.x(x_60), .z(tmp00_60_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060061(.x(x_61), .z(tmp00_61_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060062(.x(x_62), .z(tmp00_62_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060063(.x(x_63), .z(tmp00_63_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060064(.x(x_64), .z(tmp00_64_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060065(.x(x_65), .z(tmp00_65_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060066(.x(x_66), .z(tmp00_66_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060067(.x(x_67), .z(tmp00_67_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060068(.x(x_68), .z(tmp00_68_6));
	booth_0002 #(.WIDTH(WIDTH)) mul00060069(.x(x_69), .z(tmp00_69_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060070(.x(x_70), .z(tmp00_70_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060071(.x(x_71), .z(tmp00_71_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060072(.x(x_72), .z(tmp00_72_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060073(.x(x_73), .z(tmp00_73_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060074(.x(x_74), .z(tmp00_74_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060075(.x(x_75), .z(tmp00_75_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060076(.x(x_76), .z(tmp00_76_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060077(.x(x_77), .z(tmp00_77_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060078(.x(x_78), .z(tmp00_78_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060079(.x(x_79), .z(tmp00_79_6));
	booth__004 #(.WIDTH(WIDTH)) mul00060080(.x(x_80), .z(tmp00_80_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060081(.x(x_81), .z(tmp00_81_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00060082(.x(x_82), .z(tmp00_82_6));
	booth_0004 #(.WIDTH(WIDTH)) mul00060083(.x(x_83), .z(tmp00_83_6));
	booth_0000 #(.WIDTH(WIDTH)) mul00070000(.x(x_0), .z(tmp00_0_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070001(.x(x_1), .z(tmp00_1_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070002(.x(x_2), .z(tmp00_2_7));
	booth__002 #(.WIDTH(WIDTH)) mul00070003(.x(x_3), .z(tmp00_3_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070004(.x(x_4), .z(tmp00_4_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070005(.x(x_5), .z(tmp00_5_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070006(.x(x_6), .z(tmp00_6_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070007(.x(x_7), .z(tmp00_7_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070008(.x(x_8), .z(tmp00_8_7));
	booth__006 #(.WIDTH(WIDTH)) mul00070009(.x(x_9), .z(tmp00_9_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070010(.x(x_10), .z(tmp00_10_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070011(.x(x_11), .z(tmp00_11_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070012(.x(x_12), .z(tmp00_12_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070013(.x(x_13), .z(tmp00_13_7));
	booth__002 #(.WIDTH(WIDTH)) mul00070014(.x(x_14), .z(tmp00_14_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070015(.x(x_15), .z(tmp00_15_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070016(.x(x_16), .z(tmp00_16_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070017(.x(x_17), .z(tmp00_17_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070018(.x(x_18), .z(tmp00_18_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070019(.x(x_19), .z(tmp00_19_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070020(.x(x_20), .z(tmp00_20_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070021(.x(x_21), .z(tmp00_21_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070022(.x(x_22), .z(tmp00_22_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070023(.x(x_23), .z(tmp00_23_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070024(.x(x_24), .z(tmp00_24_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070025(.x(x_25), .z(tmp00_25_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070026(.x(x_26), .z(tmp00_26_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070027(.x(x_27), .z(tmp00_27_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070028(.x(x_28), .z(tmp00_28_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070029(.x(x_29), .z(tmp00_29_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070030(.x(x_30), .z(tmp00_30_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070031(.x(x_31), .z(tmp00_31_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070032(.x(x_32), .z(tmp00_32_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070033(.x(x_33), .z(tmp00_33_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070034(.x(x_34), .z(tmp00_34_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070035(.x(x_35), .z(tmp00_35_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070036(.x(x_36), .z(tmp00_36_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070037(.x(x_37), .z(tmp00_37_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070038(.x(x_38), .z(tmp00_38_7));
	booth_0002 #(.WIDTH(WIDTH)) mul00070039(.x(x_39), .z(tmp00_39_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070040(.x(x_40), .z(tmp00_40_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070041(.x(x_41), .z(tmp00_41_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070042(.x(x_42), .z(tmp00_42_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070043(.x(x_43), .z(tmp00_43_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070044(.x(x_44), .z(tmp00_44_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070045(.x(x_45), .z(tmp00_45_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070046(.x(x_46), .z(tmp00_46_7));
	booth_0002 #(.WIDTH(WIDTH)) mul00070047(.x(x_47), .z(tmp00_47_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070048(.x(x_48), .z(tmp00_48_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070049(.x(x_49), .z(tmp00_49_7));
	booth__006 #(.WIDTH(WIDTH)) mul00070050(.x(x_50), .z(tmp00_50_7));
	booth__006 #(.WIDTH(WIDTH)) mul00070051(.x(x_51), .z(tmp00_51_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070052(.x(x_52), .z(tmp00_52_7));
	booth__002 #(.WIDTH(WIDTH)) mul00070053(.x(x_53), .z(tmp00_53_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070054(.x(x_54), .z(tmp00_54_7));
	booth_0006 #(.WIDTH(WIDTH)) mul00070055(.x(x_55), .z(tmp00_55_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070056(.x(x_56), .z(tmp00_56_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070057(.x(x_57), .z(tmp00_57_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070058(.x(x_58), .z(tmp00_58_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070059(.x(x_59), .z(tmp00_59_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070060(.x(x_60), .z(tmp00_60_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070061(.x(x_61), .z(tmp00_61_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070062(.x(x_62), .z(tmp00_62_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070063(.x(x_63), .z(tmp00_63_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070064(.x(x_64), .z(tmp00_64_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070065(.x(x_65), .z(tmp00_65_7));
	booth__002 #(.WIDTH(WIDTH)) mul00070066(.x(x_66), .z(tmp00_66_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070067(.x(x_67), .z(tmp00_67_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070068(.x(x_68), .z(tmp00_68_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070069(.x(x_69), .z(tmp00_69_7));
	booth__004 #(.WIDTH(WIDTH)) mul00070070(.x(x_70), .z(tmp00_70_7));
	booth__010 #(.WIDTH(WIDTH)) mul00070071(.x(x_71), .z(tmp00_71_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070072(.x(x_72), .z(tmp00_72_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070073(.x(x_73), .z(tmp00_73_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070074(.x(x_74), .z(tmp00_74_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070075(.x(x_75), .z(tmp00_75_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070076(.x(x_76), .z(tmp00_76_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070077(.x(x_77), .z(tmp00_77_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070078(.x(x_78), .z(tmp00_78_7));
	booth_0004 #(.WIDTH(WIDTH)) mul00070079(.x(x_79), .z(tmp00_79_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070080(.x(x_80), .z(tmp00_80_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070081(.x(x_81), .z(tmp00_81_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070082(.x(x_82), .z(tmp00_82_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00070083(.x(x_83), .z(tmp00_83_7));
	booth_0000 #(.WIDTH(WIDTH)) mul00080000(.x(x_0), .z(tmp00_0_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080001(.x(x_1), .z(tmp00_1_8));
	booth__006 #(.WIDTH(WIDTH)) mul00080002(.x(x_2), .z(tmp00_2_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080003(.x(x_3), .z(tmp00_3_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080004(.x(x_4), .z(tmp00_4_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080005(.x(x_5), .z(tmp00_5_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080006(.x(x_6), .z(tmp00_6_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080007(.x(x_7), .z(tmp00_7_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080008(.x(x_8), .z(tmp00_8_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080009(.x(x_9), .z(tmp00_9_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080010(.x(x_10), .z(tmp00_10_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080011(.x(x_11), .z(tmp00_11_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080012(.x(x_12), .z(tmp00_12_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080013(.x(x_13), .z(tmp00_13_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080014(.x(x_14), .z(tmp00_14_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080015(.x(x_15), .z(tmp00_15_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080016(.x(x_16), .z(tmp00_16_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080017(.x(x_17), .z(tmp00_17_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080018(.x(x_18), .z(tmp00_18_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080019(.x(x_19), .z(tmp00_19_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080020(.x(x_20), .z(tmp00_20_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080021(.x(x_21), .z(tmp00_21_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080022(.x(x_22), .z(tmp00_22_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080023(.x(x_23), .z(tmp00_23_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080024(.x(x_24), .z(tmp00_24_8));
	booth__006 #(.WIDTH(WIDTH)) mul00080025(.x(x_25), .z(tmp00_25_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080026(.x(x_26), .z(tmp00_26_8));
	booth_0006 #(.WIDTH(WIDTH)) mul00080027(.x(x_27), .z(tmp00_27_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080028(.x(x_28), .z(tmp00_28_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080029(.x(x_29), .z(tmp00_29_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080030(.x(x_30), .z(tmp00_30_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080031(.x(x_31), .z(tmp00_31_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080032(.x(x_32), .z(tmp00_32_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080033(.x(x_33), .z(tmp00_33_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080034(.x(x_34), .z(tmp00_34_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080035(.x(x_35), .z(tmp00_35_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080036(.x(x_36), .z(tmp00_36_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080037(.x(x_37), .z(tmp00_37_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080038(.x(x_38), .z(tmp00_38_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080039(.x(x_39), .z(tmp00_39_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080040(.x(x_40), .z(tmp00_40_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080041(.x(x_41), .z(tmp00_41_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080042(.x(x_42), .z(tmp00_42_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080043(.x(x_43), .z(tmp00_43_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080044(.x(x_44), .z(tmp00_44_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080045(.x(x_45), .z(tmp00_45_8));
	booth__002 #(.WIDTH(WIDTH)) mul00080046(.x(x_46), .z(tmp00_46_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080047(.x(x_47), .z(tmp00_47_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080048(.x(x_48), .z(tmp00_48_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080049(.x(x_49), .z(tmp00_49_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080050(.x(x_50), .z(tmp00_50_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080051(.x(x_51), .z(tmp00_51_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080052(.x(x_52), .z(tmp00_52_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080053(.x(x_53), .z(tmp00_53_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080054(.x(x_54), .z(tmp00_54_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080055(.x(x_55), .z(tmp00_55_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080056(.x(x_56), .z(tmp00_56_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080057(.x(x_57), .z(tmp00_57_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080058(.x(x_58), .z(tmp00_58_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080059(.x(x_59), .z(tmp00_59_8));
	booth__006 #(.WIDTH(WIDTH)) mul00080060(.x(x_60), .z(tmp00_60_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080061(.x(x_61), .z(tmp00_61_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080062(.x(x_62), .z(tmp00_62_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080063(.x(x_63), .z(tmp00_63_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080064(.x(x_64), .z(tmp00_64_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080065(.x(x_65), .z(tmp00_65_8));
	booth_0008 #(.WIDTH(WIDTH)) mul00080066(.x(x_66), .z(tmp00_66_8));
	booth_0012 #(.WIDTH(WIDTH)) mul00080067(.x(x_67), .z(tmp00_67_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080068(.x(x_68), .z(tmp00_68_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080069(.x(x_69), .z(tmp00_69_8));
	booth_0004 #(.WIDTH(WIDTH)) mul00080070(.x(x_70), .z(tmp00_70_8));
	booth_0006 #(.WIDTH(WIDTH)) mul00080071(.x(x_71), .z(tmp00_71_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080072(.x(x_72), .z(tmp00_72_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080073(.x(x_73), .z(tmp00_73_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080074(.x(x_74), .z(tmp00_74_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080075(.x(x_75), .z(tmp00_75_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080076(.x(x_76), .z(tmp00_76_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080077(.x(x_77), .z(tmp00_77_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080078(.x(x_78), .z(tmp00_78_8));
	booth_0000 #(.WIDTH(WIDTH)) mul00080079(.x(x_79), .z(tmp00_79_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080080(.x(x_80), .z(tmp00_80_8));
	booth_0002 #(.WIDTH(WIDTH)) mul00080081(.x(x_81), .z(tmp00_81_8));
	booth__008 #(.WIDTH(WIDTH)) mul00080082(.x(x_82), .z(tmp00_82_8));
	booth__004 #(.WIDTH(WIDTH)) mul00080083(.x(x_83), .z(tmp00_83_8));
	booth__002 #(.WIDTH(WIDTH)) mul00090000(.x(x_0), .z(tmp00_0_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090001(.x(x_1), .z(tmp00_1_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090002(.x(x_2), .z(tmp00_2_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090003(.x(x_3), .z(tmp00_3_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090004(.x(x_4), .z(tmp00_4_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090005(.x(x_5), .z(tmp00_5_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090006(.x(x_6), .z(tmp00_6_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090007(.x(x_7), .z(tmp00_7_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090008(.x(x_8), .z(tmp00_8_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090009(.x(x_9), .z(tmp00_9_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090010(.x(x_10), .z(tmp00_10_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090011(.x(x_11), .z(tmp00_11_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090012(.x(x_12), .z(tmp00_12_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090013(.x(x_13), .z(tmp00_13_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090014(.x(x_14), .z(tmp00_14_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090015(.x(x_15), .z(tmp00_15_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090016(.x(x_16), .z(tmp00_16_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090017(.x(x_17), .z(tmp00_17_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090018(.x(x_18), .z(tmp00_18_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090019(.x(x_19), .z(tmp00_19_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090020(.x(x_20), .z(tmp00_20_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090021(.x(x_21), .z(tmp00_21_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090022(.x(x_22), .z(tmp00_22_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090023(.x(x_23), .z(tmp00_23_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090024(.x(x_24), .z(tmp00_24_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090025(.x(x_25), .z(tmp00_25_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090026(.x(x_26), .z(tmp00_26_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090027(.x(x_27), .z(tmp00_27_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090028(.x(x_28), .z(tmp00_28_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090029(.x(x_29), .z(tmp00_29_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090030(.x(x_30), .z(tmp00_30_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090031(.x(x_31), .z(tmp00_31_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090032(.x(x_32), .z(tmp00_32_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090033(.x(x_33), .z(tmp00_33_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090034(.x(x_34), .z(tmp00_34_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090035(.x(x_35), .z(tmp00_35_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090036(.x(x_36), .z(tmp00_36_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090037(.x(x_37), .z(tmp00_37_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090038(.x(x_38), .z(tmp00_38_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090039(.x(x_39), .z(tmp00_39_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090040(.x(x_40), .z(tmp00_40_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090041(.x(x_41), .z(tmp00_41_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090042(.x(x_42), .z(tmp00_42_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090043(.x(x_43), .z(tmp00_43_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090044(.x(x_44), .z(tmp00_44_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090045(.x(x_45), .z(tmp00_45_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090046(.x(x_46), .z(tmp00_46_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090047(.x(x_47), .z(tmp00_47_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090048(.x(x_48), .z(tmp00_48_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090049(.x(x_49), .z(tmp00_49_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090050(.x(x_50), .z(tmp00_50_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090051(.x(x_51), .z(tmp00_51_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090052(.x(x_52), .z(tmp00_52_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090053(.x(x_53), .z(tmp00_53_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090054(.x(x_54), .z(tmp00_54_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090055(.x(x_55), .z(tmp00_55_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090056(.x(x_56), .z(tmp00_56_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090057(.x(x_57), .z(tmp00_57_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090058(.x(x_58), .z(tmp00_58_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090059(.x(x_59), .z(tmp00_59_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090060(.x(x_60), .z(tmp00_60_9));
	booth__004 #(.WIDTH(WIDTH)) mul00090061(.x(x_61), .z(tmp00_61_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090062(.x(x_62), .z(tmp00_62_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090063(.x(x_63), .z(tmp00_63_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090064(.x(x_64), .z(tmp00_64_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090065(.x(x_65), .z(tmp00_65_9));
	booth_0008 #(.WIDTH(WIDTH)) mul00090066(.x(x_66), .z(tmp00_66_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090067(.x(x_67), .z(tmp00_67_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090068(.x(x_68), .z(tmp00_68_9));
	booth_0006 #(.WIDTH(WIDTH)) mul00090069(.x(x_69), .z(tmp00_69_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090070(.x(x_70), .z(tmp00_70_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090071(.x(x_71), .z(tmp00_71_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090072(.x(x_72), .z(tmp00_72_9));
	booth__008 #(.WIDTH(WIDTH)) mul00090073(.x(x_73), .z(tmp00_73_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090074(.x(x_74), .z(tmp00_74_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090075(.x(x_75), .z(tmp00_75_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090076(.x(x_76), .z(tmp00_76_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090077(.x(x_77), .z(tmp00_77_9));
	booth_0004 #(.WIDTH(WIDTH)) mul00090078(.x(x_78), .z(tmp00_78_9));
	booth__002 #(.WIDTH(WIDTH)) mul00090079(.x(x_79), .z(tmp00_79_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090080(.x(x_80), .z(tmp00_80_9));
	booth_0000 #(.WIDTH(WIDTH)) mul00090081(.x(x_81), .z(tmp00_81_9));
	booth_0002 #(.WIDTH(WIDTH)) mul00090082(.x(x_82), .z(tmp00_82_9));
	booth__006 #(.WIDTH(WIDTH)) mul00090083(.x(x_83), .z(tmp00_83_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000000(.in0(tmp00_0_0), .in1(tmp00_1_0), .out(tmp01_0_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000001(.in0(tmp00_2_0), .in1(tmp00_3_0), .out(tmp01_1_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000002(.in0(tmp00_4_0), .in1(tmp00_5_0), .out(tmp01_2_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000003(.in0(tmp00_6_0), .in1(tmp00_7_0), .out(tmp01_3_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000004(.in0(tmp00_8_0), .in1(tmp00_9_0), .out(tmp01_4_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000005(.in0(tmp00_10_0), .in1(tmp00_11_0), .out(tmp01_5_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000006(.in0(tmp00_12_0), .in1(tmp00_13_0), .out(tmp01_6_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000007(.in0(tmp00_14_0), .in1(tmp00_15_0), .out(tmp01_7_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000008(.in0(tmp00_16_0), .in1(tmp00_17_0), .out(tmp01_8_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000009(.in0(tmp00_18_0), .in1(tmp00_19_0), .out(tmp01_9_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000010(.in0(tmp00_20_0), .in1(tmp00_21_0), .out(tmp01_10_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000011(.in0(tmp00_22_0), .in1(tmp00_23_0), .out(tmp01_11_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000012(.in0(tmp00_24_0), .in1(tmp00_25_0), .out(tmp01_12_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000013(.in0(tmp00_26_0), .in1(tmp00_27_0), .out(tmp01_13_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000014(.in0(tmp00_28_0), .in1(tmp00_29_0), .out(tmp01_14_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000015(.in0(tmp00_30_0), .in1(tmp00_31_0), .out(tmp01_15_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000016(.in0(tmp00_32_0), .in1(tmp00_33_0), .out(tmp01_16_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000017(.in0(tmp00_34_0), .in1(tmp00_35_0), .out(tmp01_17_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000018(.in0(tmp00_36_0), .in1(tmp00_37_0), .out(tmp01_18_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000019(.in0(tmp00_38_0), .in1(tmp00_39_0), .out(tmp01_19_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000020(.in0(tmp00_40_0), .in1(tmp00_41_0), .out(tmp01_20_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000021(.in0(tmp00_42_0), .in1(tmp00_43_0), .out(tmp01_21_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000022(.in0(tmp00_44_0), .in1(tmp00_45_0), .out(tmp01_22_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000023(.in0(tmp00_46_0), .in1(tmp00_47_0), .out(tmp01_23_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000024(.in0(tmp00_48_0), .in1(tmp00_49_0), .out(tmp01_24_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000025(.in0(tmp00_50_0), .in1(tmp00_51_0), .out(tmp01_25_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000026(.in0(tmp00_52_0), .in1(tmp00_53_0), .out(tmp01_26_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000027(.in0(tmp00_54_0), .in1(tmp00_55_0), .out(tmp01_27_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000028(.in0(tmp00_56_0), .in1(tmp00_57_0), .out(tmp01_28_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000029(.in0(tmp00_58_0), .in1(tmp00_59_0), .out(tmp01_29_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000030(.in0(tmp00_60_0), .in1(tmp00_61_0), .out(tmp01_30_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000031(.in0(tmp00_62_0), .in1(tmp00_63_0), .out(tmp01_31_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000032(.in0(tmp00_64_0), .in1(tmp00_65_0), .out(tmp01_32_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000033(.in0(tmp00_66_0), .in1(tmp00_67_0), .out(tmp01_33_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000034(.in0(tmp00_68_0), .in1(tmp00_69_0), .out(tmp01_34_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000035(.in0(tmp00_70_0), .in1(tmp00_71_0), .out(tmp01_35_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000036(.in0(tmp00_72_0), .in1(tmp00_73_0), .out(tmp01_36_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000037(.in0(tmp00_74_0), .in1(tmp00_75_0), .out(tmp01_37_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000038(.in0(tmp00_76_0), .in1(tmp00_77_0), .out(tmp01_38_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000039(.in0(tmp00_78_0), .in1(tmp00_79_0), .out(tmp01_39_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000040(.in0(tmp00_80_0), .in1(tmp00_81_0), .out(tmp01_40_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000041(.in0(tmp00_82_0), .in1(tmp00_83_0), .out(tmp01_41_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000042(.in0(tmp01_0_0), .in1(tmp01_1_0), .out(tmp02_0_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000043(.in0(tmp01_2_0), .in1(tmp01_3_0), .out(tmp02_1_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000044(.in0(tmp01_4_0), .in1(tmp01_5_0), .out(tmp02_2_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000045(.in0(tmp01_6_0), .in1(tmp01_7_0), .out(tmp02_3_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000046(.in0(tmp01_8_0), .in1(tmp01_9_0), .out(tmp02_4_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000047(.in0(tmp01_10_0), .in1(tmp01_11_0), .out(tmp02_5_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000048(.in0(tmp01_12_0), .in1(tmp01_13_0), .out(tmp02_6_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000049(.in0(tmp01_14_0), .in1(tmp01_15_0), .out(tmp02_7_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000050(.in0(tmp01_16_0), .in1(tmp01_17_0), .out(tmp02_8_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000051(.in0(tmp01_18_0), .in1(tmp01_19_0), .out(tmp02_9_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000052(.in0(tmp01_20_0), .in1(tmp01_21_0), .out(tmp02_10_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000053(.in0(tmp01_22_0), .in1(tmp01_23_0), .out(tmp02_11_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000054(.in0(tmp01_24_0), .in1(tmp01_25_0), .out(tmp02_12_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000055(.in0(tmp01_26_0), .in1(tmp01_27_0), .out(tmp02_13_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000056(.in0(tmp01_28_0), .in1(tmp01_29_0), .out(tmp02_14_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000057(.in0(tmp01_30_0), .in1(tmp01_31_0), .out(tmp02_15_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000058(.in0(tmp01_32_0), .in1(tmp01_33_0), .out(tmp02_16_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000059(.in0(tmp01_34_0), .in1(tmp01_35_0), .out(tmp02_17_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000060(.in0(tmp01_36_0), .in1(tmp01_37_0), .out(tmp02_18_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000061(.in0(tmp01_38_0), .in1(tmp01_39_0), .out(tmp02_19_0));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000062(.in0(tmp01_40_0), .in1(tmp01_41_0), .out(tmp02_20_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000063(.in0(tmp02_0_0), .in1(tmp02_1_0), .out(tmp03_0_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000064(.in0(tmp02_2_0), .in1(tmp02_3_0), .out(tmp03_1_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000065(.in0(tmp02_4_0), .in1(tmp02_5_0), .out(tmp03_2_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000066(.in0(tmp02_6_0), .in1(tmp02_7_0), .out(tmp03_3_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000067(.in0(tmp02_8_0), .in1(tmp02_9_0), .out(tmp03_4_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000068(.in0(tmp02_10_0), .in1(tmp02_11_0), .out(tmp03_5_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000069(.in0(tmp02_12_0), .in1(tmp02_13_0), .out(tmp03_6_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000070(.in0(tmp02_14_0), .in1(tmp02_15_0), .out(tmp03_7_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000071(.in0(tmp02_16_0), .in1(tmp02_17_0), .out(tmp03_8_0));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000072(.in0(tmp02_18_0), .in1(tmp02_19_0), .out(tmp03_9_0));
	assign tmp03_10_0 = $signed(tmp02_20_0);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000073(.in0(tmp03_0_0), .in1(tmp03_1_0), .out(tmp04_0_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000074(.in0(tmp03_2_0), .in1(tmp03_3_0), .out(tmp04_1_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000075(.in0(tmp03_4_0), .in1(tmp03_5_0), .out(tmp04_2_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000076(.in0(tmp03_6_0), .in1(tmp03_7_0), .out(tmp04_3_0));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000077(.in0(tmp03_8_0), .in1(tmp03_9_0), .out(tmp04_4_0));
	assign tmp04_5_0 = $signed(tmp03_10_0);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000078(.in0(tmp04_0_0), .in1(tmp04_1_0), .out(tmp05_0_0));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000079(.in0(tmp04_2_0), .in1(tmp04_3_0), .out(tmp05_1_0));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000080(.in0(tmp04_4_0), .in1(tmp04_5_0), .out(tmp05_2_0));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000081(.in0(tmp05_0_0), .in1(tmp05_1_0), .out(tmp06_0_0));
	assign tmp06_1_0 = $signed(tmp05_2_0);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000082(.in0(tmp06_0_0), .in1(tmp06_1_0), .out(tmp07_0_0));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000083(.in0(tmp00_0_1), .in1(tmp00_1_1), .out(tmp01_0_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000084(.in0(tmp00_2_1), .in1(tmp00_3_1), .out(tmp01_1_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000085(.in0(tmp00_4_1), .in1(tmp00_5_1), .out(tmp01_2_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000086(.in0(tmp00_6_1), .in1(tmp00_7_1), .out(tmp01_3_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000087(.in0(tmp00_8_1), .in1(tmp00_9_1), .out(tmp01_4_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000088(.in0(tmp00_10_1), .in1(tmp00_11_1), .out(tmp01_5_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000089(.in0(tmp00_12_1), .in1(tmp00_13_1), .out(tmp01_6_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000090(.in0(tmp00_14_1), .in1(tmp00_15_1), .out(tmp01_7_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000091(.in0(tmp00_16_1), .in1(tmp00_17_1), .out(tmp01_8_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000092(.in0(tmp00_18_1), .in1(tmp00_19_1), .out(tmp01_9_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000093(.in0(tmp00_20_1), .in1(tmp00_21_1), .out(tmp01_10_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000094(.in0(tmp00_22_1), .in1(tmp00_23_1), .out(tmp01_11_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000095(.in0(tmp00_24_1), .in1(tmp00_25_1), .out(tmp01_12_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000096(.in0(tmp00_26_1), .in1(tmp00_27_1), .out(tmp01_13_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000097(.in0(tmp00_28_1), .in1(tmp00_29_1), .out(tmp01_14_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000098(.in0(tmp00_30_1), .in1(tmp00_31_1), .out(tmp01_15_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000099(.in0(tmp00_32_1), .in1(tmp00_33_1), .out(tmp01_16_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000100(.in0(tmp00_34_1), .in1(tmp00_35_1), .out(tmp01_17_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000101(.in0(tmp00_36_1), .in1(tmp00_37_1), .out(tmp01_18_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000102(.in0(tmp00_38_1), .in1(tmp00_39_1), .out(tmp01_19_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000103(.in0(tmp00_40_1), .in1(tmp00_41_1), .out(tmp01_20_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000104(.in0(tmp00_42_1), .in1(tmp00_43_1), .out(tmp01_21_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000105(.in0(tmp00_44_1), .in1(tmp00_45_1), .out(tmp01_22_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000106(.in0(tmp00_46_1), .in1(tmp00_47_1), .out(tmp01_23_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000107(.in0(tmp00_48_1), .in1(tmp00_49_1), .out(tmp01_24_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000108(.in0(tmp00_50_1), .in1(tmp00_51_1), .out(tmp01_25_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000109(.in0(tmp00_52_1), .in1(tmp00_53_1), .out(tmp01_26_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000110(.in0(tmp00_54_1), .in1(tmp00_55_1), .out(tmp01_27_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000111(.in0(tmp00_56_1), .in1(tmp00_57_1), .out(tmp01_28_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000112(.in0(tmp00_58_1), .in1(tmp00_59_1), .out(tmp01_29_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000113(.in0(tmp00_60_1), .in1(tmp00_61_1), .out(tmp01_30_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000114(.in0(tmp00_62_1), .in1(tmp00_63_1), .out(tmp01_31_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000115(.in0(tmp00_64_1), .in1(tmp00_65_1), .out(tmp01_32_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000116(.in0(tmp00_66_1), .in1(tmp00_67_1), .out(tmp01_33_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000117(.in0(tmp00_68_1), .in1(tmp00_69_1), .out(tmp01_34_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000118(.in0(tmp00_70_1), .in1(tmp00_71_1), .out(tmp01_35_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000119(.in0(tmp00_72_1), .in1(tmp00_73_1), .out(tmp01_36_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000120(.in0(tmp00_74_1), .in1(tmp00_75_1), .out(tmp01_37_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000121(.in0(tmp00_76_1), .in1(tmp00_77_1), .out(tmp01_38_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000122(.in0(tmp00_78_1), .in1(tmp00_79_1), .out(tmp01_39_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000123(.in0(tmp00_80_1), .in1(tmp00_81_1), .out(tmp01_40_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000124(.in0(tmp00_82_1), .in1(tmp00_83_1), .out(tmp01_41_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000125(.in0(tmp01_0_1), .in1(tmp01_1_1), .out(tmp02_0_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000126(.in0(tmp01_2_1), .in1(tmp01_3_1), .out(tmp02_1_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000127(.in0(tmp01_4_1), .in1(tmp01_5_1), .out(tmp02_2_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000128(.in0(tmp01_6_1), .in1(tmp01_7_1), .out(tmp02_3_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000129(.in0(tmp01_8_1), .in1(tmp01_9_1), .out(tmp02_4_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000130(.in0(tmp01_10_1), .in1(tmp01_11_1), .out(tmp02_5_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000131(.in0(tmp01_12_1), .in1(tmp01_13_1), .out(tmp02_6_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000132(.in0(tmp01_14_1), .in1(tmp01_15_1), .out(tmp02_7_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000133(.in0(tmp01_16_1), .in1(tmp01_17_1), .out(tmp02_8_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000134(.in0(tmp01_18_1), .in1(tmp01_19_1), .out(tmp02_9_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000135(.in0(tmp01_20_1), .in1(tmp01_21_1), .out(tmp02_10_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000136(.in0(tmp01_22_1), .in1(tmp01_23_1), .out(tmp02_11_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000137(.in0(tmp01_24_1), .in1(tmp01_25_1), .out(tmp02_12_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000138(.in0(tmp01_26_1), .in1(tmp01_27_1), .out(tmp02_13_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000139(.in0(tmp01_28_1), .in1(tmp01_29_1), .out(tmp02_14_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000140(.in0(tmp01_30_1), .in1(tmp01_31_1), .out(tmp02_15_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000141(.in0(tmp01_32_1), .in1(tmp01_33_1), .out(tmp02_16_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000142(.in0(tmp01_34_1), .in1(tmp01_35_1), .out(tmp02_17_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000143(.in0(tmp01_36_1), .in1(tmp01_37_1), .out(tmp02_18_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000144(.in0(tmp01_38_1), .in1(tmp01_39_1), .out(tmp02_19_1));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000145(.in0(tmp01_40_1), .in1(tmp01_41_1), .out(tmp02_20_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000146(.in0(tmp02_0_1), .in1(tmp02_1_1), .out(tmp03_0_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000147(.in0(tmp02_2_1), .in1(tmp02_3_1), .out(tmp03_1_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000148(.in0(tmp02_4_1), .in1(tmp02_5_1), .out(tmp03_2_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000149(.in0(tmp02_6_1), .in1(tmp02_7_1), .out(tmp03_3_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000150(.in0(tmp02_8_1), .in1(tmp02_9_1), .out(tmp03_4_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000151(.in0(tmp02_10_1), .in1(tmp02_11_1), .out(tmp03_5_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000152(.in0(tmp02_12_1), .in1(tmp02_13_1), .out(tmp03_6_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000153(.in0(tmp02_14_1), .in1(tmp02_15_1), .out(tmp03_7_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000154(.in0(tmp02_16_1), .in1(tmp02_17_1), .out(tmp03_8_1));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000155(.in0(tmp02_18_1), .in1(tmp02_19_1), .out(tmp03_9_1));
	assign tmp03_10_1 = $signed(tmp02_20_1);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000156(.in0(tmp03_0_1), .in1(tmp03_1_1), .out(tmp04_0_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000157(.in0(tmp03_2_1), .in1(tmp03_3_1), .out(tmp04_1_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000158(.in0(tmp03_4_1), .in1(tmp03_5_1), .out(tmp04_2_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000159(.in0(tmp03_6_1), .in1(tmp03_7_1), .out(tmp04_3_1));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000160(.in0(tmp03_8_1), .in1(tmp03_9_1), .out(tmp04_4_1));
	assign tmp04_5_1 = $signed(tmp03_10_1);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000161(.in0(tmp04_0_1), .in1(tmp04_1_1), .out(tmp05_0_1));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000162(.in0(tmp04_2_1), .in1(tmp04_3_1), .out(tmp05_1_1));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000163(.in0(tmp04_4_1), .in1(tmp04_5_1), .out(tmp05_2_1));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000164(.in0(tmp05_0_1), .in1(tmp05_1_1), .out(tmp06_0_1));
	assign tmp06_1_1 = $signed(tmp05_2_1);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000165(.in0(tmp06_0_1), .in1(tmp06_1_1), .out(tmp07_0_1));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000166(.in0(tmp00_0_2), .in1(tmp00_1_2), .out(tmp01_0_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000167(.in0(tmp00_2_2), .in1(tmp00_3_2), .out(tmp01_1_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000168(.in0(tmp00_4_2), .in1(tmp00_5_2), .out(tmp01_2_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000169(.in0(tmp00_6_2), .in1(tmp00_7_2), .out(tmp01_3_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000170(.in0(tmp00_8_2), .in1(tmp00_9_2), .out(tmp01_4_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000171(.in0(tmp00_10_2), .in1(tmp00_11_2), .out(tmp01_5_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000172(.in0(tmp00_12_2), .in1(tmp00_13_2), .out(tmp01_6_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000173(.in0(tmp00_14_2), .in1(tmp00_15_2), .out(tmp01_7_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000174(.in0(tmp00_16_2), .in1(tmp00_17_2), .out(tmp01_8_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000175(.in0(tmp00_18_2), .in1(tmp00_19_2), .out(tmp01_9_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000176(.in0(tmp00_20_2), .in1(tmp00_21_2), .out(tmp01_10_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000177(.in0(tmp00_22_2), .in1(tmp00_23_2), .out(tmp01_11_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000178(.in0(tmp00_24_2), .in1(tmp00_25_2), .out(tmp01_12_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000179(.in0(tmp00_26_2), .in1(tmp00_27_2), .out(tmp01_13_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000180(.in0(tmp00_28_2), .in1(tmp00_29_2), .out(tmp01_14_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000181(.in0(tmp00_30_2), .in1(tmp00_31_2), .out(tmp01_15_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000182(.in0(tmp00_32_2), .in1(tmp00_33_2), .out(tmp01_16_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000183(.in0(tmp00_34_2), .in1(tmp00_35_2), .out(tmp01_17_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000184(.in0(tmp00_36_2), .in1(tmp00_37_2), .out(tmp01_18_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000185(.in0(tmp00_38_2), .in1(tmp00_39_2), .out(tmp01_19_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000186(.in0(tmp00_40_2), .in1(tmp00_41_2), .out(tmp01_20_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000187(.in0(tmp00_42_2), .in1(tmp00_43_2), .out(tmp01_21_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000188(.in0(tmp00_44_2), .in1(tmp00_45_2), .out(tmp01_22_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000189(.in0(tmp00_46_2), .in1(tmp00_47_2), .out(tmp01_23_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000190(.in0(tmp00_48_2), .in1(tmp00_49_2), .out(tmp01_24_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000191(.in0(tmp00_50_2), .in1(tmp00_51_2), .out(tmp01_25_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000192(.in0(tmp00_52_2), .in1(tmp00_53_2), .out(tmp01_26_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000193(.in0(tmp00_54_2), .in1(tmp00_55_2), .out(tmp01_27_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000194(.in0(tmp00_56_2), .in1(tmp00_57_2), .out(tmp01_28_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000195(.in0(tmp00_58_2), .in1(tmp00_59_2), .out(tmp01_29_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000196(.in0(tmp00_60_2), .in1(tmp00_61_2), .out(tmp01_30_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000197(.in0(tmp00_62_2), .in1(tmp00_63_2), .out(tmp01_31_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000198(.in0(tmp00_64_2), .in1(tmp00_65_2), .out(tmp01_32_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000199(.in0(tmp00_66_2), .in1(tmp00_67_2), .out(tmp01_33_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000200(.in0(tmp00_68_2), .in1(tmp00_69_2), .out(tmp01_34_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000201(.in0(tmp00_70_2), .in1(tmp00_71_2), .out(tmp01_35_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000202(.in0(tmp00_72_2), .in1(tmp00_73_2), .out(tmp01_36_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000203(.in0(tmp00_74_2), .in1(tmp00_75_2), .out(tmp01_37_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000204(.in0(tmp00_76_2), .in1(tmp00_77_2), .out(tmp01_38_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000205(.in0(tmp00_78_2), .in1(tmp00_79_2), .out(tmp01_39_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000206(.in0(tmp00_80_2), .in1(tmp00_81_2), .out(tmp01_40_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000207(.in0(tmp00_82_2), .in1(tmp00_83_2), .out(tmp01_41_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000208(.in0(tmp01_0_2), .in1(tmp01_1_2), .out(tmp02_0_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000209(.in0(tmp01_2_2), .in1(tmp01_3_2), .out(tmp02_1_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000210(.in0(tmp01_4_2), .in1(tmp01_5_2), .out(tmp02_2_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000211(.in0(tmp01_6_2), .in1(tmp01_7_2), .out(tmp02_3_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000212(.in0(tmp01_8_2), .in1(tmp01_9_2), .out(tmp02_4_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000213(.in0(tmp01_10_2), .in1(tmp01_11_2), .out(tmp02_5_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000214(.in0(tmp01_12_2), .in1(tmp01_13_2), .out(tmp02_6_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000215(.in0(tmp01_14_2), .in1(tmp01_15_2), .out(tmp02_7_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000216(.in0(tmp01_16_2), .in1(tmp01_17_2), .out(tmp02_8_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000217(.in0(tmp01_18_2), .in1(tmp01_19_2), .out(tmp02_9_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000218(.in0(tmp01_20_2), .in1(tmp01_21_2), .out(tmp02_10_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000219(.in0(tmp01_22_2), .in1(tmp01_23_2), .out(tmp02_11_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000220(.in0(tmp01_24_2), .in1(tmp01_25_2), .out(tmp02_12_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000221(.in0(tmp01_26_2), .in1(tmp01_27_2), .out(tmp02_13_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000222(.in0(tmp01_28_2), .in1(tmp01_29_2), .out(tmp02_14_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000223(.in0(tmp01_30_2), .in1(tmp01_31_2), .out(tmp02_15_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000224(.in0(tmp01_32_2), .in1(tmp01_33_2), .out(tmp02_16_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000225(.in0(tmp01_34_2), .in1(tmp01_35_2), .out(tmp02_17_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000226(.in0(tmp01_36_2), .in1(tmp01_37_2), .out(tmp02_18_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000227(.in0(tmp01_38_2), .in1(tmp01_39_2), .out(tmp02_19_2));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000228(.in0(tmp01_40_2), .in1(tmp01_41_2), .out(tmp02_20_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000229(.in0(tmp02_0_2), .in1(tmp02_1_2), .out(tmp03_0_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000230(.in0(tmp02_2_2), .in1(tmp02_3_2), .out(tmp03_1_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000231(.in0(tmp02_4_2), .in1(tmp02_5_2), .out(tmp03_2_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000232(.in0(tmp02_6_2), .in1(tmp02_7_2), .out(tmp03_3_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000233(.in0(tmp02_8_2), .in1(tmp02_9_2), .out(tmp03_4_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000234(.in0(tmp02_10_2), .in1(tmp02_11_2), .out(tmp03_5_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000235(.in0(tmp02_12_2), .in1(tmp02_13_2), .out(tmp03_6_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000236(.in0(tmp02_14_2), .in1(tmp02_15_2), .out(tmp03_7_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000237(.in0(tmp02_16_2), .in1(tmp02_17_2), .out(tmp03_8_2));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000238(.in0(tmp02_18_2), .in1(tmp02_19_2), .out(tmp03_9_2));
	assign tmp03_10_2 = $signed(tmp02_20_2);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000239(.in0(tmp03_0_2), .in1(tmp03_1_2), .out(tmp04_0_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000240(.in0(tmp03_2_2), .in1(tmp03_3_2), .out(tmp04_1_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000241(.in0(tmp03_4_2), .in1(tmp03_5_2), .out(tmp04_2_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000242(.in0(tmp03_6_2), .in1(tmp03_7_2), .out(tmp04_3_2));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000243(.in0(tmp03_8_2), .in1(tmp03_9_2), .out(tmp04_4_2));
	assign tmp04_5_2 = $signed(tmp03_10_2);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000244(.in0(tmp04_0_2), .in1(tmp04_1_2), .out(tmp05_0_2));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000245(.in0(tmp04_2_2), .in1(tmp04_3_2), .out(tmp05_1_2));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000246(.in0(tmp04_4_2), .in1(tmp04_5_2), .out(tmp05_2_2));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000247(.in0(tmp05_0_2), .in1(tmp05_1_2), .out(tmp06_0_2));
	assign tmp06_1_2 = $signed(tmp05_2_2);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000248(.in0(tmp06_0_2), .in1(tmp06_1_2), .out(tmp07_0_2));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000249(.in0(tmp00_0_3), .in1(tmp00_1_3), .out(tmp01_0_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000250(.in0(tmp00_2_3), .in1(tmp00_3_3), .out(tmp01_1_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000251(.in0(tmp00_4_3), .in1(tmp00_5_3), .out(tmp01_2_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000252(.in0(tmp00_6_3), .in1(tmp00_7_3), .out(tmp01_3_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000253(.in0(tmp00_8_3), .in1(tmp00_9_3), .out(tmp01_4_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000254(.in0(tmp00_10_3), .in1(tmp00_11_3), .out(tmp01_5_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000255(.in0(tmp00_12_3), .in1(tmp00_13_3), .out(tmp01_6_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000256(.in0(tmp00_14_3), .in1(tmp00_15_3), .out(tmp01_7_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000257(.in0(tmp00_16_3), .in1(tmp00_17_3), .out(tmp01_8_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000258(.in0(tmp00_18_3), .in1(tmp00_19_3), .out(tmp01_9_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000259(.in0(tmp00_20_3), .in1(tmp00_21_3), .out(tmp01_10_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000260(.in0(tmp00_22_3), .in1(tmp00_23_3), .out(tmp01_11_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000261(.in0(tmp00_24_3), .in1(tmp00_25_3), .out(tmp01_12_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000262(.in0(tmp00_26_3), .in1(tmp00_27_3), .out(tmp01_13_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000263(.in0(tmp00_28_3), .in1(tmp00_29_3), .out(tmp01_14_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000264(.in0(tmp00_30_3), .in1(tmp00_31_3), .out(tmp01_15_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000265(.in0(tmp00_32_3), .in1(tmp00_33_3), .out(tmp01_16_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000266(.in0(tmp00_34_3), .in1(tmp00_35_3), .out(tmp01_17_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000267(.in0(tmp00_36_3), .in1(tmp00_37_3), .out(tmp01_18_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000268(.in0(tmp00_38_3), .in1(tmp00_39_3), .out(tmp01_19_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000269(.in0(tmp00_40_3), .in1(tmp00_41_3), .out(tmp01_20_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000270(.in0(tmp00_42_3), .in1(tmp00_43_3), .out(tmp01_21_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000271(.in0(tmp00_44_3), .in1(tmp00_45_3), .out(tmp01_22_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000272(.in0(tmp00_46_3), .in1(tmp00_47_3), .out(tmp01_23_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000273(.in0(tmp00_48_3), .in1(tmp00_49_3), .out(tmp01_24_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000274(.in0(tmp00_50_3), .in1(tmp00_51_3), .out(tmp01_25_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000275(.in0(tmp00_52_3), .in1(tmp00_53_3), .out(tmp01_26_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000276(.in0(tmp00_54_3), .in1(tmp00_55_3), .out(tmp01_27_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000277(.in0(tmp00_56_3), .in1(tmp00_57_3), .out(tmp01_28_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000278(.in0(tmp00_58_3), .in1(tmp00_59_3), .out(tmp01_29_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000279(.in0(tmp00_60_3), .in1(tmp00_61_3), .out(tmp01_30_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000280(.in0(tmp00_62_3), .in1(tmp00_63_3), .out(tmp01_31_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000281(.in0(tmp00_64_3), .in1(tmp00_65_3), .out(tmp01_32_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000282(.in0(tmp00_66_3), .in1(tmp00_67_3), .out(tmp01_33_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000283(.in0(tmp00_68_3), .in1(tmp00_69_3), .out(tmp01_34_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000284(.in0(tmp00_70_3), .in1(tmp00_71_3), .out(tmp01_35_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000285(.in0(tmp00_72_3), .in1(tmp00_73_3), .out(tmp01_36_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000286(.in0(tmp00_74_3), .in1(tmp00_75_3), .out(tmp01_37_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000287(.in0(tmp00_76_3), .in1(tmp00_77_3), .out(tmp01_38_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000288(.in0(tmp00_78_3), .in1(tmp00_79_3), .out(tmp01_39_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000289(.in0(tmp00_80_3), .in1(tmp00_81_3), .out(tmp01_40_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000290(.in0(tmp00_82_3), .in1(tmp00_83_3), .out(tmp01_41_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000291(.in0(tmp01_0_3), .in1(tmp01_1_3), .out(tmp02_0_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000292(.in0(tmp01_2_3), .in1(tmp01_3_3), .out(tmp02_1_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000293(.in0(tmp01_4_3), .in1(tmp01_5_3), .out(tmp02_2_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000294(.in0(tmp01_6_3), .in1(tmp01_7_3), .out(tmp02_3_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000295(.in0(tmp01_8_3), .in1(tmp01_9_3), .out(tmp02_4_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000296(.in0(tmp01_10_3), .in1(tmp01_11_3), .out(tmp02_5_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000297(.in0(tmp01_12_3), .in1(tmp01_13_3), .out(tmp02_6_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000298(.in0(tmp01_14_3), .in1(tmp01_15_3), .out(tmp02_7_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000299(.in0(tmp01_16_3), .in1(tmp01_17_3), .out(tmp02_8_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000300(.in0(tmp01_18_3), .in1(tmp01_19_3), .out(tmp02_9_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000301(.in0(tmp01_20_3), .in1(tmp01_21_3), .out(tmp02_10_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000302(.in0(tmp01_22_3), .in1(tmp01_23_3), .out(tmp02_11_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000303(.in0(tmp01_24_3), .in1(tmp01_25_3), .out(tmp02_12_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000304(.in0(tmp01_26_3), .in1(tmp01_27_3), .out(tmp02_13_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000305(.in0(tmp01_28_3), .in1(tmp01_29_3), .out(tmp02_14_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000306(.in0(tmp01_30_3), .in1(tmp01_31_3), .out(tmp02_15_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000307(.in0(tmp01_32_3), .in1(tmp01_33_3), .out(tmp02_16_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000308(.in0(tmp01_34_3), .in1(tmp01_35_3), .out(tmp02_17_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000309(.in0(tmp01_36_3), .in1(tmp01_37_3), .out(tmp02_18_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000310(.in0(tmp01_38_3), .in1(tmp01_39_3), .out(tmp02_19_3));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000311(.in0(tmp01_40_3), .in1(tmp01_41_3), .out(tmp02_20_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000312(.in0(tmp02_0_3), .in1(tmp02_1_3), .out(tmp03_0_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000313(.in0(tmp02_2_3), .in1(tmp02_3_3), .out(tmp03_1_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000314(.in0(tmp02_4_3), .in1(tmp02_5_3), .out(tmp03_2_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000315(.in0(tmp02_6_3), .in1(tmp02_7_3), .out(tmp03_3_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000316(.in0(tmp02_8_3), .in1(tmp02_9_3), .out(tmp03_4_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000317(.in0(tmp02_10_3), .in1(tmp02_11_3), .out(tmp03_5_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000318(.in0(tmp02_12_3), .in1(tmp02_13_3), .out(tmp03_6_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000319(.in0(tmp02_14_3), .in1(tmp02_15_3), .out(tmp03_7_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000320(.in0(tmp02_16_3), .in1(tmp02_17_3), .out(tmp03_8_3));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000321(.in0(tmp02_18_3), .in1(tmp02_19_3), .out(tmp03_9_3));
	assign tmp03_10_3 = $signed(tmp02_20_3);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000322(.in0(tmp03_0_3), .in1(tmp03_1_3), .out(tmp04_0_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000323(.in0(tmp03_2_3), .in1(tmp03_3_3), .out(tmp04_1_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000324(.in0(tmp03_4_3), .in1(tmp03_5_3), .out(tmp04_2_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000325(.in0(tmp03_6_3), .in1(tmp03_7_3), .out(tmp04_3_3));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000326(.in0(tmp03_8_3), .in1(tmp03_9_3), .out(tmp04_4_3));
	assign tmp04_5_3 = $signed(tmp03_10_3);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000327(.in0(tmp04_0_3), .in1(tmp04_1_3), .out(tmp05_0_3));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000328(.in0(tmp04_2_3), .in1(tmp04_3_3), .out(tmp05_1_3));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000329(.in0(tmp04_4_3), .in1(tmp04_5_3), .out(tmp05_2_3));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000330(.in0(tmp05_0_3), .in1(tmp05_1_3), .out(tmp06_0_3));
	assign tmp06_1_3 = $signed(tmp05_2_3);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000331(.in0(tmp06_0_3), .in1(tmp06_1_3), .out(tmp07_0_3));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000332(.in0(tmp00_0_4), .in1(tmp00_1_4), .out(tmp01_0_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000333(.in0(tmp00_2_4), .in1(tmp00_3_4), .out(tmp01_1_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000334(.in0(tmp00_4_4), .in1(tmp00_5_4), .out(tmp01_2_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000335(.in0(tmp00_6_4), .in1(tmp00_7_4), .out(tmp01_3_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000336(.in0(tmp00_8_4), .in1(tmp00_9_4), .out(tmp01_4_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000337(.in0(tmp00_10_4), .in1(tmp00_11_4), .out(tmp01_5_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000338(.in0(tmp00_12_4), .in1(tmp00_13_4), .out(tmp01_6_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000339(.in0(tmp00_14_4), .in1(tmp00_15_4), .out(tmp01_7_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000340(.in0(tmp00_16_4), .in1(tmp00_17_4), .out(tmp01_8_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000341(.in0(tmp00_18_4), .in1(tmp00_19_4), .out(tmp01_9_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000342(.in0(tmp00_20_4), .in1(tmp00_21_4), .out(tmp01_10_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000343(.in0(tmp00_22_4), .in1(tmp00_23_4), .out(tmp01_11_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000344(.in0(tmp00_24_4), .in1(tmp00_25_4), .out(tmp01_12_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000345(.in0(tmp00_26_4), .in1(tmp00_27_4), .out(tmp01_13_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000346(.in0(tmp00_28_4), .in1(tmp00_29_4), .out(tmp01_14_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000347(.in0(tmp00_30_4), .in1(tmp00_31_4), .out(tmp01_15_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000348(.in0(tmp00_32_4), .in1(tmp00_33_4), .out(tmp01_16_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000349(.in0(tmp00_34_4), .in1(tmp00_35_4), .out(tmp01_17_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000350(.in0(tmp00_36_4), .in1(tmp00_37_4), .out(tmp01_18_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000351(.in0(tmp00_38_4), .in1(tmp00_39_4), .out(tmp01_19_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000352(.in0(tmp00_40_4), .in1(tmp00_41_4), .out(tmp01_20_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000353(.in0(tmp00_42_4), .in1(tmp00_43_4), .out(tmp01_21_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000354(.in0(tmp00_44_4), .in1(tmp00_45_4), .out(tmp01_22_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000355(.in0(tmp00_46_4), .in1(tmp00_47_4), .out(tmp01_23_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000356(.in0(tmp00_48_4), .in1(tmp00_49_4), .out(tmp01_24_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000357(.in0(tmp00_50_4), .in1(tmp00_51_4), .out(tmp01_25_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000358(.in0(tmp00_52_4), .in1(tmp00_53_4), .out(tmp01_26_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000359(.in0(tmp00_54_4), .in1(tmp00_55_4), .out(tmp01_27_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000360(.in0(tmp00_56_4), .in1(tmp00_57_4), .out(tmp01_28_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000361(.in0(tmp00_58_4), .in1(tmp00_59_4), .out(tmp01_29_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000362(.in0(tmp00_60_4), .in1(tmp00_61_4), .out(tmp01_30_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000363(.in0(tmp00_62_4), .in1(tmp00_63_4), .out(tmp01_31_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000364(.in0(tmp00_64_4), .in1(tmp00_65_4), .out(tmp01_32_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000365(.in0(tmp00_66_4), .in1(tmp00_67_4), .out(tmp01_33_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000366(.in0(tmp00_68_4), .in1(tmp00_69_4), .out(tmp01_34_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000367(.in0(tmp00_70_4), .in1(tmp00_71_4), .out(tmp01_35_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000368(.in0(tmp00_72_4), .in1(tmp00_73_4), .out(tmp01_36_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000369(.in0(tmp00_74_4), .in1(tmp00_75_4), .out(tmp01_37_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000370(.in0(tmp00_76_4), .in1(tmp00_77_4), .out(tmp01_38_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000371(.in0(tmp00_78_4), .in1(tmp00_79_4), .out(tmp01_39_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000372(.in0(tmp00_80_4), .in1(tmp00_81_4), .out(tmp01_40_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000373(.in0(tmp00_82_4), .in1(tmp00_83_4), .out(tmp01_41_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000374(.in0(tmp01_0_4), .in1(tmp01_1_4), .out(tmp02_0_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000375(.in0(tmp01_2_4), .in1(tmp01_3_4), .out(tmp02_1_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000376(.in0(tmp01_4_4), .in1(tmp01_5_4), .out(tmp02_2_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000377(.in0(tmp01_6_4), .in1(tmp01_7_4), .out(tmp02_3_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000378(.in0(tmp01_8_4), .in1(tmp01_9_4), .out(tmp02_4_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000379(.in0(tmp01_10_4), .in1(tmp01_11_4), .out(tmp02_5_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000380(.in0(tmp01_12_4), .in1(tmp01_13_4), .out(tmp02_6_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000381(.in0(tmp01_14_4), .in1(tmp01_15_4), .out(tmp02_7_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000382(.in0(tmp01_16_4), .in1(tmp01_17_4), .out(tmp02_8_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000383(.in0(tmp01_18_4), .in1(tmp01_19_4), .out(tmp02_9_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000384(.in0(tmp01_20_4), .in1(tmp01_21_4), .out(tmp02_10_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000385(.in0(tmp01_22_4), .in1(tmp01_23_4), .out(tmp02_11_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000386(.in0(tmp01_24_4), .in1(tmp01_25_4), .out(tmp02_12_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000387(.in0(tmp01_26_4), .in1(tmp01_27_4), .out(tmp02_13_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000388(.in0(tmp01_28_4), .in1(tmp01_29_4), .out(tmp02_14_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000389(.in0(tmp01_30_4), .in1(tmp01_31_4), .out(tmp02_15_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000390(.in0(tmp01_32_4), .in1(tmp01_33_4), .out(tmp02_16_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000391(.in0(tmp01_34_4), .in1(tmp01_35_4), .out(tmp02_17_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000392(.in0(tmp01_36_4), .in1(tmp01_37_4), .out(tmp02_18_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000393(.in0(tmp01_38_4), .in1(tmp01_39_4), .out(tmp02_19_4));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000394(.in0(tmp01_40_4), .in1(tmp01_41_4), .out(tmp02_20_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000395(.in0(tmp02_0_4), .in1(tmp02_1_4), .out(tmp03_0_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000396(.in0(tmp02_2_4), .in1(tmp02_3_4), .out(tmp03_1_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000397(.in0(tmp02_4_4), .in1(tmp02_5_4), .out(tmp03_2_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000398(.in0(tmp02_6_4), .in1(tmp02_7_4), .out(tmp03_3_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000399(.in0(tmp02_8_4), .in1(tmp02_9_4), .out(tmp03_4_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000400(.in0(tmp02_10_4), .in1(tmp02_11_4), .out(tmp03_5_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000401(.in0(tmp02_12_4), .in1(tmp02_13_4), .out(tmp03_6_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000402(.in0(tmp02_14_4), .in1(tmp02_15_4), .out(tmp03_7_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000403(.in0(tmp02_16_4), .in1(tmp02_17_4), .out(tmp03_8_4));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000404(.in0(tmp02_18_4), .in1(tmp02_19_4), .out(tmp03_9_4));
	assign tmp03_10_4 = $signed(tmp02_20_4);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000405(.in0(tmp03_0_4), .in1(tmp03_1_4), .out(tmp04_0_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000406(.in0(tmp03_2_4), .in1(tmp03_3_4), .out(tmp04_1_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000407(.in0(tmp03_4_4), .in1(tmp03_5_4), .out(tmp04_2_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000408(.in0(tmp03_6_4), .in1(tmp03_7_4), .out(tmp04_3_4));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000409(.in0(tmp03_8_4), .in1(tmp03_9_4), .out(tmp04_4_4));
	assign tmp04_5_4 = $signed(tmp03_10_4);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000410(.in0(tmp04_0_4), .in1(tmp04_1_4), .out(tmp05_0_4));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000411(.in0(tmp04_2_4), .in1(tmp04_3_4), .out(tmp05_1_4));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000412(.in0(tmp04_4_4), .in1(tmp04_5_4), .out(tmp05_2_4));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000413(.in0(tmp05_0_4), .in1(tmp05_1_4), .out(tmp06_0_4));
	assign tmp06_1_4 = $signed(tmp05_2_4);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000414(.in0(tmp06_0_4), .in1(tmp06_1_4), .out(tmp07_0_4));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000415(.in0(tmp00_0_5), .in1(tmp00_1_5), .out(tmp01_0_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000416(.in0(tmp00_2_5), .in1(tmp00_3_5), .out(tmp01_1_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000417(.in0(tmp00_4_5), .in1(tmp00_5_5), .out(tmp01_2_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000418(.in0(tmp00_6_5), .in1(tmp00_7_5), .out(tmp01_3_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000419(.in0(tmp00_8_5), .in1(tmp00_9_5), .out(tmp01_4_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000420(.in0(tmp00_10_5), .in1(tmp00_11_5), .out(tmp01_5_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000421(.in0(tmp00_12_5), .in1(tmp00_13_5), .out(tmp01_6_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000422(.in0(tmp00_14_5), .in1(tmp00_15_5), .out(tmp01_7_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000423(.in0(tmp00_16_5), .in1(tmp00_17_5), .out(tmp01_8_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000424(.in0(tmp00_18_5), .in1(tmp00_19_5), .out(tmp01_9_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000425(.in0(tmp00_20_5), .in1(tmp00_21_5), .out(tmp01_10_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000426(.in0(tmp00_22_5), .in1(tmp00_23_5), .out(tmp01_11_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000427(.in0(tmp00_24_5), .in1(tmp00_25_5), .out(tmp01_12_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000428(.in0(tmp00_26_5), .in1(tmp00_27_5), .out(tmp01_13_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000429(.in0(tmp00_28_5), .in1(tmp00_29_5), .out(tmp01_14_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000430(.in0(tmp00_30_5), .in1(tmp00_31_5), .out(tmp01_15_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000431(.in0(tmp00_32_5), .in1(tmp00_33_5), .out(tmp01_16_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000432(.in0(tmp00_34_5), .in1(tmp00_35_5), .out(tmp01_17_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000433(.in0(tmp00_36_5), .in1(tmp00_37_5), .out(tmp01_18_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000434(.in0(tmp00_38_5), .in1(tmp00_39_5), .out(tmp01_19_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000435(.in0(tmp00_40_5), .in1(tmp00_41_5), .out(tmp01_20_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000436(.in0(tmp00_42_5), .in1(tmp00_43_5), .out(tmp01_21_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000437(.in0(tmp00_44_5), .in1(tmp00_45_5), .out(tmp01_22_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000438(.in0(tmp00_46_5), .in1(tmp00_47_5), .out(tmp01_23_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000439(.in0(tmp00_48_5), .in1(tmp00_49_5), .out(tmp01_24_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000440(.in0(tmp00_50_5), .in1(tmp00_51_5), .out(tmp01_25_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000441(.in0(tmp00_52_5), .in1(tmp00_53_5), .out(tmp01_26_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000442(.in0(tmp00_54_5), .in1(tmp00_55_5), .out(tmp01_27_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000443(.in0(tmp00_56_5), .in1(tmp00_57_5), .out(tmp01_28_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000444(.in0(tmp00_58_5), .in1(tmp00_59_5), .out(tmp01_29_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000445(.in0(tmp00_60_5), .in1(tmp00_61_5), .out(tmp01_30_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000446(.in0(tmp00_62_5), .in1(tmp00_63_5), .out(tmp01_31_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000447(.in0(tmp00_64_5), .in1(tmp00_65_5), .out(tmp01_32_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000448(.in0(tmp00_66_5), .in1(tmp00_67_5), .out(tmp01_33_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000449(.in0(tmp00_68_5), .in1(tmp00_69_5), .out(tmp01_34_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000450(.in0(tmp00_70_5), .in1(tmp00_71_5), .out(tmp01_35_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000451(.in0(tmp00_72_5), .in1(tmp00_73_5), .out(tmp01_36_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000452(.in0(tmp00_74_5), .in1(tmp00_75_5), .out(tmp01_37_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000453(.in0(tmp00_76_5), .in1(tmp00_77_5), .out(tmp01_38_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000454(.in0(tmp00_78_5), .in1(tmp00_79_5), .out(tmp01_39_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000455(.in0(tmp00_80_5), .in1(tmp00_81_5), .out(tmp01_40_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000456(.in0(tmp00_82_5), .in1(tmp00_83_5), .out(tmp01_41_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000457(.in0(tmp01_0_5), .in1(tmp01_1_5), .out(tmp02_0_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000458(.in0(tmp01_2_5), .in1(tmp01_3_5), .out(tmp02_1_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000459(.in0(tmp01_4_5), .in1(tmp01_5_5), .out(tmp02_2_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000460(.in0(tmp01_6_5), .in1(tmp01_7_5), .out(tmp02_3_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000461(.in0(tmp01_8_5), .in1(tmp01_9_5), .out(tmp02_4_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000462(.in0(tmp01_10_5), .in1(tmp01_11_5), .out(tmp02_5_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000463(.in0(tmp01_12_5), .in1(tmp01_13_5), .out(tmp02_6_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000464(.in0(tmp01_14_5), .in1(tmp01_15_5), .out(tmp02_7_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000465(.in0(tmp01_16_5), .in1(tmp01_17_5), .out(tmp02_8_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000466(.in0(tmp01_18_5), .in1(tmp01_19_5), .out(tmp02_9_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000467(.in0(tmp01_20_5), .in1(tmp01_21_5), .out(tmp02_10_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000468(.in0(tmp01_22_5), .in1(tmp01_23_5), .out(tmp02_11_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000469(.in0(tmp01_24_5), .in1(tmp01_25_5), .out(tmp02_12_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000470(.in0(tmp01_26_5), .in1(tmp01_27_5), .out(tmp02_13_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000471(.in0(tmp01_28_5), .in1(tmp01_29_5), .out(tmp02_14_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000472(.in0(tmp01_30_5), .in1(tmp01_31_5), .out(tmp02_15_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000473(.in0(tmp01_32_5), .in1(tmp01_33_5), .out(tmp02_16_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000474(.in0(tmp01_34_5), .in1(tmp01_35_5), .out(tmp02_17_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000475(.in0(tmp01_36_5), .in1(tmp01_37_5), .out(tmp02_18_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000476(.in0(tmp01_38_5), .in1(tmp01_39_5), .out(tmp02_19_5));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000477(.in0(tmp01_40_5), .in1(tmp01_41_5), .out(tmp02_20_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000478(.in0(tmp02_0_5), .in1(tmp02_1_5), .out(tmp03_0_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000479(.in0(tmp02_2_5), .in1(tmp02_3_5), .out(tmp03_1_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000480(.in0(tmp02_4_5), .in1(tmp02_5_5), .out(tmp03_2_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000481(.in0(tmp02_6_5), .in1(tmp02_7_5), .out(tmp03_3_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000482(.in0(tmp02_8_5), .in1(tmp02_9_5), .out(tmp03_4_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000483(.in0(tmp02_10_5), .in1(tmp02_11_5), .out(tmp03_5_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000484(.in0(tmp02_12_5), .in1(tmp02_13_5), .out(tmp03_6_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000485(.in0(tmp02_14_5), .in1(tmp02_15_5), .out(tmp03_7_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000486(.in0(tmp02_16_5), .in1(tmp02_17_5), .out(tmp03_8_5));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000487(.in0(tmp02_18_5), .in1(tmp02_19_5), .out(tmp03_9_5));
	assign tmp03_10_5 = $signed(tmp02_20_5);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000488(.in0(tmp03_0_5), .in1(tmp03_1_5), .out(tmp04_0_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000489(.in0(tmp03_2_5), .in1(tmp03_3_5), .out(tmp04_1_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000490(.in0(tmp03_4_5), .in1(tmp03_5_5), .out(tmp04_2_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000491(.in0(tmp03_6_5), .in1(tmp03_7_5), .out(tmp04_3_5));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000492(.in0(tmp03_8_5), .in1(tmp03_9_5), .out(tmp04_4_5));
	assign tmp04_5_5 = $signed(tmp03_10_5);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000493(.in0(tmp04_0_5), .in1(tmp04_1_5), .out(tmp05_0_5));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000494(.in0(tmp04_2_5), .in1(tmp04_3_5), .out(tmp05_1_5));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000495(.in0(tmp04_4_5), .in1(tmp04_5_5), .out(tmp05_2_5));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000496(.in0(tmp05_0_5), .in1(tmp05_1_5), .out(tmp06_0_5));
	assign tmp06_1_5 = $signed(tmp05_2_5);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000497(.in0(tmp06_0_5), .in1(tmp06_1_5), .out(tmp07_0_5));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000498(.in0(tmp00_0_6), .in1(tmp00_1_6), .out(tmp01_0_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000499(.in0(tmp00_2_6), .in1(tmp00_3_6), .out(tmp01_1_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000500(.in0(tmp00_4_6), .in1(tmp00_5_6), .out(tmp01_2_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000501(.in0(tmp00_6_6), .in1(tmp00_7_6), .out(tmp01_3_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000502(.in0(tmp00_8_6), .in1(tmp00_9_6), .out(tmp01_4_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000503(.in0(tmp00_10_6), .in1(tmp00_11_6), .out(tmp01_5_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000504(.in0(tmp00_12_6), .in1(tmp00_13_6), .out(tmp01_6_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000505(.in0(tmp00_14_6), .in1(tmp00_15_6), .out(tmp01_7_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000506(.in0(tmp00_16_6), .in1(tmp00_17_6), .out(tmp01_8_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000507(.in0(tmp00_18_6), .in1(tmp00_19_6), .out(tmp01_9_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000508(.in0(tmp00_20_6), .in1(tmp00_21_6), .out(tmp01_10_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000509(.in0(tmp00_22_6), .in1(tmp00_23_6), .out(tmp01_11_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000510(.in0(tmp00_24_6), .in1(tmp00_25_6), .out(tmp01_12_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000511(.in0(tmp00_26_6), .in1(tmp00_27_6), .out(tmp01_13_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000512(.in0(tmp00_28_6), .in1(tmp00_29_6), .out(tmp01_14_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000513(.in0(tmp00_30_6), .in1(tmp00_31_6), .out(tmp01_15_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000514(.in0(tmp00_32_6), .in1(tmp00_33_6), .out(tmp01_16_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000515(.in0(tmp00_34_6), .in1(tmp00_35_6), .out(tmp01_17_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000516(.in0(tmp00_36_6), .in1(tmp00_37_6), .out(tmp01_18_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000517(.in0(tmp00_38_6), .in1(tmp00_39_6), .out(tmp01_19_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000518(.in0(tmp00_40_6), .in1(tmp00_41_6), .out(tmp01_20_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000519(.in0(tmp00_42_6), .in1(tmp00_43_6), .out(tmp01_21_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000520(.in0(tmp00_44_6), .in1(tmp00_45_6), .out(tmp01_22_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000521(.in0(tmp00_46_6), .in1(tmp00_47_6), .out(tmp01_23_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000522(.in0(tmp00_48_6), .in1(tmp00_49_6), .out(tmp01_24_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000523(.in0(tmp00_50_6), .in1(tmp00_51_6), .out(tmp01_25_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000524(.in0(tmp00_52_6), .in1(tmp00_53_6), .out(tmp01_26_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000525(.in0(tmp00_54_6), .in1(tmp00_55_6), .out(tmp01_27_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000526(.in0(tmp00_56_6), .in1(tmp00_57_6), .out(tmp01_28_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000527(.in0(tmp00_58_6), .in1(tmp00_59_6), .out(tmp01_29_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000528(.in0(tmp00_60_6), .in1(tmp00_61_6), .out(tmp01_30_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000529(.in0(tmp00_62_6), .in1(tmp00_63_6), .out(tmp01_31_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000530(.in0(tmp00_64_6), .in1(tmp00_65_6), .out(tmp01_32_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000531(.in0(tmp00_66_6), .in1(tmp00_67_6), .out(tmp01_33_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000532(.in0(tmp00_68_6), .in1(tmp00_69_6), .out(tmp01_34_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000533(.in0(tmp00_70_6), .in1(tmp00_71_6), .out(tmp01_35_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000534(.in0(tmp00_72_6), .in1(tmp00_73_6), .out(tmp01_36_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000535(.in0(tmp00_74_6), .in1(tmp00_75_6), .out(tmp01_37_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000536(.in0(tmp00_76_6), .in1(tmp00_77_6), .out(tmp01_38_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000537(.in0(tmp00_78_6), .in1(tmp00_79_6), .out(tmp01_39_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000538(.in0(tmp00_80_6), .in1(tmp00_81_6), .out(tmp01_40_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000539(.in0(tmp00_82_6), .in1(tmp00_83_6), .out(tmp01_41_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000540(.in0(tmp01_0_6), .in1(tmp01_1_6), .out(tmp02_0_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000541(.in0(tmp01_2_6), .in1(tmp01_3_6), .out(tmp02_1_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000542(.in0(tmp01_4_6), .in1(tmp01_5_6), .out(tmp02_2_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000543(.in0(tmp01_6_6), .in1(tmp01_7_6), .out(tmp02_3_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000544(.in0(tmp01_8_6), .in1(tmp01_9_6), .out(tmp02_4_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000545(.in0(tmp01_10_6), .in1(tmp01_11_6), .out(tmp02_5_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000546(.in0(tmp01_12_6), .in1(tmp01_13_6), .out(tmp02_6_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000547(.in0(tmp01_14_6), .in1(tmp01_15_6), .out(tmp02_7_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000548(.in0(tmp01_16_6), .in1(tmp01_17_6), .out(tmp02_8_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000549(.in0(tmp01_18_6), .in1(tmp01_19_6), .out(tmp02_9_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000550(.in0(tmp01_20_6), .in1(tmp01_21_6), .out(tmp02_10_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000551(.in0(tmp01_22_6), .in1(tmp01_23_6), .out(tmp02_11_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000552(.in0(tmp01_24_6), .in1(tmp01_25_6), .out(tmp02_12_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000553(.in0(tmp01_26_6), .in1(tmp01_27_6), .out(tmp02_13_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000554(.in0(tmp01_28_6), .in1(tmp01_29_6), .out(tmp02_14_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000555(.in0(tmp01_30_6), .in1(tmp01_31_6), .out(tmp02_15_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000556(.in0(tmp01_32_6), .in1(tmp01_33_6), .out(tmp02_16_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000557(.in0(tmp01_34_6), .in1(tmp01_35_6), .out(tmp02_17_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000558(.in0(tmp01_36_6), .in1(tmp01_37_6), .out(tmp02_18_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000559(.in0(tmp01_38_6), .in1(tmp01_39_6), .out(tmp02_19_6));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000560(.in0(tmp01_40_6), .in1(tmp01_41_6), .out(tmp02_20_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000561(.in0(tmp02_0_6), .in1(tmp02_1_6), .out(tmp03_0_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000562(.in0(tmp02_2_6), .in1(tmp02_3_6), .out(tmp03_1_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000563(.in0(tmp02_4_6), .in1(tmp02_5_6), .out(tmp03_2_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000564(.in0(tmp02_6_6), .in1(tmp02_7_6), .out(tmp03_3_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000565(.in0(tmp02_8_6), .in1(tmp02_9_6), .out(tmp03_4_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000566(.in0(tmp02_10_6), .in1(tmp02_11_6), .out(tmp03_5_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000567(.in0(tmp02_12_6), .in1(tmp02_13_6), .out(tmp03_6_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000568(.in0(tmp02_14_6), .in1(tmp02_15_6), .out(tmp03_7_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000569(.in0(tmp02_16_6), .in1(tmp02_17_6), .out(tmp03_8_6));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000570(.in0(tmp02_18_6), .in1(tmp02_19_6), .out(tmp03_9_6));
	assign tmp03_10_6 = $signed(tmp02_20_6);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000571(.in0(tmp03_0_6), .in1(tmp03_1_6), .out(tmp04_0_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000572(.in0(tmp03_2_6), .in1(tmp03_3_6), .out(tmp04_1_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000573(.in0(tmp03_4_6), .in1(tmp03_5_6), .out(tmp04_2_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000574(.in0(tmp03_6_6), .in1(tmp03_7_6), .out(tmp04_3_6));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000575(.in0(tmp03_8_6), .in1(tmp03_9_6), .out(tmp04_4_6));
	assign tmp04_5_6 = $signed(tmp03_10_6);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000576(.in0(tmp04_0_6), .in1(tmp04_1_6), .out(tmp05_0_6));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000577(.in0(tmp04_2_6), .in1(tmp04_3_6), .out(tmp05_1_6));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000578(.in0(tmp04_4_6), .in1(tmp04_5_6), .out(tmp05_2_6));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000579(.in0(tmp05_0_6), .in1(tmp05_1_6), .out(tmp06_0_6));
	assign tmp06_1_6 = $signed(tmp05_2_6);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000580(.in0(tmp06_0_6), .in1(tmp06_1_6), .out(tmp07_0_6));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000581(.in0(tmp00_0_7), .in1(tmp00_1_7), .out(tmp01_0_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000582(.in0(tmp00_2_7), .in1(tmp00_3_7), .out(tmp01_1_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000583(.in0(tmp00_4_7), .in1(tmp00_5_7), .out(tmp01_2_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000584(.in0(tmp00_6_7), .in1(tmp00_7_7), .out(tmp01_3_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000585(.in0(tmp00_8_7), .in1(tmp00_9_7), .out(tmp01_4_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000586(.in0(tmp00_10_7), .in1(tmp00_11_7), .out(tmp01_5_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000587(.in0(tmp00_12_7), .in1(tmp00_13_7), .out(tmp01_6_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000588(.in0(tmp00_14_7), .in1(tmp00_15_7), .out(tmp01_7_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000589(.in0(tmp00_16_7), .in1(tmp00_17_7), .out(tmp01_8_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000590(.in0(tmp00_18_7), .in1(tmp00_19_7), .out(tmp01_9_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000591(.in0(tmp00_20_7), .in1(tmp00_21_7), .out(tmp01_10_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000592(.in0(tmp00_22_7), .in1(tmp00_23_7), .out(tmp01_11_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000593(.in0(tmp00_24_7), .in1(tmp00_25_7), .out(tmp01_12_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000594(.in0(tmp00_26_7), .in1(tmp00_27_7), .out(tmp01_13_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000595(.in0(tmp00_28_7), .in1(tmp00_29_7), .out(tmp01_14_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000596(.in0(tmp00_30_7), .in1(tmp00_31_7), .out(tmp01_15_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000597(.in0(tmp00_32_7), .in1(tmp00_33_7), .out(tmp01_16_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000598(.in0(tmp00_34_7), .in1(tmp00_35_7), .out(tmp01_17_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000599(.in0(tmp00_36_7), .in1(tmp00_37_7), .out(tmp01_18_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000600(.in0(tmp00_38_7), .in1(tmp00_39_7), .out(tmp01_19_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000601(.in0(tmp00_40_7), .in1(tmp00_41_7), .out(tmp01_20_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000602(.in0(tmp00_42_7), .in1(tmp00_43_7), .out(tmp01_21_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000603(.in0(tmp00_44_7), .in1(tmp00_45_7), .out(tmp01_22_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000604(.in0(tmp00_46_7), .in1(tmp00_47_7), .out(tmp01_23_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000605(.in0(tmp00_48_7), .in1(tmp00_49_7), .out(tmp01_24_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000606(.in0(tmp00_50_7), .in1(tmp00_51_7), .out(tmp01_25_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000607(.in0(tmp00_52_7), .in1(tmp00_53_7), .out(tmp01_26_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000608(.in0(tmp00_54_7), .in1(tmp00_55_7), .out(tmp01_27_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000609(.in0(tmp00_56_7), .in1(tmp00_57_7), .out(tmp01_28_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000610(.in0(tmp00_58_7), .in1(tmp00_59_7), .out(tmp01_29_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000611(.in0(tmp00_60_7), .in1(tmp00_61_7), .out(tmp01_30_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000612(.in0(tmp00_62_7), .in1(tmp00_63_7), .out(tmp01_31_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000613(.in0(tmp00_64_7), .in1(tmp00_65_7), .out(tmp01_32_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000614(.in0(tmp00_66_7), .in1(tmp00_67_7), .out(tmp01_33_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000615(.in0(tmp00_68_7), .in1(tmp00_69_7), .out(tmp01_34_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000616(.in0(tmp00_70_7), .in1(tmp00_71_7), .out(tmp01_35_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000617(.in0(tmp00_72_7), .in1(tmp00_73_7), .out(tmp01_36_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000618(.in0(tmp00_74_7), .in1(tmp00_75_7), .out(tmp01_37_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000619(.in0(tmp00_76_7), .in1(tmp00_77_7), .out(tmp01_38_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000620(.in0(tmp00_78_7), .in1(tmp00_79_7), .out(tmp01_39_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000621(.in0(tmp00_80_7), .in1(tmp00_81_7), .out(tmp01_40_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000622(.in0(tmp00_82_7), .in1(tmp00_83_7), .out(tmp01_41_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000623(.in0(tmp01_0_7), .in1(tmp01_1_7), .out(tmp02_0_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000624(.in0(tmp01_2_7), .in1(tmp01_3_7), .out(tmp02_1_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000625(.in0(tmp01_4_7), .in1(tmp01_5_7), .out(tmp02_2_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000626(.in0(tmp01_6_7), .in1(tmp01_7_7), .out(tmp02_3_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000627(.in0(tmp01_8_7), .in1(tmp01_9_7), .out(tmp02_4_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000628(.in0(tmp01_10_7), .in1(tmp01_11_7), .out(tmp02_5_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000629(.in0(tmp01_12_7), .in1(tmp01_13_7), .out(tmp02_6_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000630(.in0(tmp01_14_7), .in1(tmp01_15_7), .out(tmp02_7_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000631(.in0(tmp01_16_7), .in1(tmp01_17_7), .out(tmp02_8_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000632(.in0(tmp01_18_7), .in1(tmp01_19_7), .out(tmp02_9_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000633(.in0(tmp01_20_7), .in1(tmp01_21_7), .out(tmp02_10_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000634(.in0(tmp01_22_7), .in1(tmp01_23_7), .out(tmp02_11_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000635(.in0(tmp01_24_7), .in1(tmp01_25_7), .out(tmp02_12_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000636(.in0(tmp01_26_7), .in1(tmp01_27_7), .out(tmp02_13_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000637(.in0(tmp01_28_7), .in1(tmp01_29_7), .out(tmp02_14_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000638(.in0(tmp01_30_7), .in1(tmp01_31_7), .out(tmp02_15_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000639(.in0(tmp01_32_7), .in1(tmp01_33_7), .out(tmp02_16_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000640(.in0(tmp01_34_7), .in1(tmp01_35_7), .out(tmp02_17_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000641(.in0(tmp01_36_7), .in1(tmp01_37_7), .out(tmp02_18_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000642(.in0(tmp01_38_7), .in1(tmp01_39_7), .out(tmp02_19_7));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000643(.in0(tmp01_40_7), .in1(tmp01_41_7), .out(tmp02_20_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000644(.in0(tmp02_0_7), .in1(tmp02_1_7), .out(tmp03_0_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000645(.in0(tmp02_2_7), .in1(tmp02_3_7), .out(tmp03_1_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000646(.in0(tmp02_4_7), .in1(tmp02_5_7), .out(tmp03_2_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000647(.in0(tmp02_6_7), .in1(tmp02_7_7), .out(tmp03_3_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000648(.in0(tmp02_8_7), .in1(tmp02_9_7), .out(tmp03_4_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000649(.in0(tmp02_10_7), .in1(tmp02_11_7), .out(tmp03_5_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000650(.in0(tmp02_12_7), .in1(tmp02_13_7), .out(tmp03_6_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000651(.in0(tmp02_14_7), .in1(tmp02_15_7), .out(tmp03_7_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000652(.in0(tmp02_16_7), .in1(tmp02_17_7), .out(tmp03_8_7));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000653(.in0(tmp02_18_7), .in1(tmp02_19_7), .out(tmp03_9_7));
	assign tmp03_10_7 = $signed(tmp02_20_7);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000654(.in0(tmp03_0_7), .in1(tmp03_1_7), .out(tmp04_0_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000655(.in0(tmp03_2_7), .in1(tmp03_3_7), .out(tmp04_1_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000656(.in0(tmp03_4_7), .in1(tmp03_5_7), .out(tmp04_2_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000657(.in0(tmp03_6_7), .in1(tmp03_7_7), .out(tmp04_3_7));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000658(.in0(tmp03_8_7), .in1(tmp03_9_7), .out(tmp04_4_7));
	assign tmp04_5_7 = $signed(tmp03_10_7);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000659(.in0(tmp04_0_7), .in1(tmp04_1_7), .out(tmp05_0_7));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000660(.in0(tmp04_2_7), .in1(tmp04_3_7), .out(tmp05_1_7));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000661(.in0(tmp04_4_7), .in1(tmp04_5_7), .out(tmp05_2_7));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000662(.in0(tmp05_0_7), .in1(tmp05_1_7), .out(tmp06_0_7));
	assign tmp06_1_7 = $signed(tmp05_2_7);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000663(.in0(tmp06_0_7), .in1(tmp06_1_7), .out(tmp07_0_7));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000664(.in0(tmp00_0_8), .in1(tmp00_1_8), .out(tmp01_0_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000665(.in0(tmp00_2_8), .in1(tmp00_3_8), .out(tmp01_1_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000666(.in0(tmp00_4_8), .in1(tmp00_5_8), .out(tmp01_2_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000667(.in0(tmp00_6_8), .in1(tmp00_7_8), .out(tmp01_3_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000668(.in0(tmp00_8_8), .in1(tmp00_9_8), .out(tmp01_4_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000669(.in0(tmp00_10_8), .in1(tmp00_11_8), .out(tmp01_5_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000670(.in0(tmp00_12_8), .in1(tmp00_13_8), .out(tmp01_6_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000671(.in0(tmp00_14_8), .in1(tmp00_15_8), .out(tmp01_7_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000672(.in0(tmp00_16_8), .in1(tmp00_17_8), .out(tmp01_8_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000673(.in0(tmp00_18_8), .in1(tmp00_19_8), .out(tmp01_9_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000674(.in0(tmp00_20_8), .in1(tmp00_21_8), .out(tmp01_10_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000675(.in0(tmp00_22_8), .in1(tmp00_23_8), .out(tmp01_11_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000676(.in0(tmp00_24_8), .in1(tmp00_25_8), .out(tmp01_12_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000677(.in0(tmp00_26_8), .in1(tmp00_27_8), .out(tmp01_13_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000678(.in0(tmp00_28_8), .in1(tmp00_29_8), .out(tmp01_14_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000679(.in0(tmp00_30_8), .in1(tmp00_31_8), .out(tmp01_15_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000680(.in0(tmp00_32_8), .in1(tmp00_33_8), .out(tmp01_16_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000681(.in0(tmp00_34_8), .in1(tmp00_35_8), .out(tmp01_17_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000682(.in0(tmp00_36_8), .in1(tmp00_37_8), .out(tmp01_18_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000683(.in0(tmp00_38_8), .in1(tmp00_39_8), .out(tmp01_19_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000684(.in0(tmp00_40_8), .in1(tmp00_41_8), .out(tmp01_20_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000685(.in0(tmp00_42_8), .in1(tmp00_43_8), .out(tmp01_21_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000686(.in0(tmp00_44_8), .in1(tmp00_45_8), .out(tmp01_22_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000687(.in0(tmp00_46_8), .in1(tmp00_47_8), .out(tmp01_23_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000688(.in0(tmp00_48_8), .in1(tmp00_49_8), .out(tmp01_24_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000689(.in0(tmp00_50_8), .in1(tmp00_51_8), .out(tmp01_25_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000690(.in0(tmp00_52_8), .in1(tmp00_53_8), .out(tmp01_26_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000691(.in0(tmp00_54_8), .in1(tmp00_55_8), .out(tmp01_27_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000692(.in0(tmp00_56_8), .in1(tmp00_57_8), .out(tmp01_28_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000693(.in0(tmp00_58_8), .in1(tmp00_59_8), .out(tmp01_29_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000694(.in0(tmp00_60_8), .in1(tmp00_61_8), .out(tmp01_30_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000695(.in0(tmp00_62_8), .in1(tmp00_63_8), .out(tmp01_31_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000696(.in0(tmp00_64_8), .in1(tmp00_65_8), .out(tmp01_32_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000697(.in0(tmp00_66_8), .in1(tmp00_67_8), .out(tmp01_33_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000698(.in0(tmp00_68_8), .in1(tmp00_69_8), .out(tmp01_34_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000699(.in0(tmp00_70_8), .in1(tmp00_71_8), .out(tmp01_35_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000700(.in0(tmp00_72_8), .in1(tmp00_73_8), .out(tmp01_36_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000701(.in0(tmp00_74_8), .in1(tmp00_75_8), .out(tmp01_37_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000702(.in0(tmp00_76_8), .in1(tmp00_77_8), .out(tmp01_38_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000703(.in0(tmp00_78_8), .in1(tmp00_79_8), .out(tmp01_39_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000704(.in0(tmp00_80_8), .in1(tmp00_81_8), .out(tmp01_40_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000705(.in0(tmp00_82_8), .in1(tmp00_83_8), .out(tmp01_41_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000706(.in0(tmp01_0_8), .in1(tmp01_1_8), .out(tmp02_0_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000707(.in0(tmp01_2_8), .in1(tmp01_3_8), .out(tmp02_1_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000708(.in0(tmp01_4_8), .in1(tmp01_5_8), .out(tmp02_2_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000709(.in0(tmp01_6_8), .in1(tmp01_7_8), .out(tmp02_3_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000710(.in0(tmp01_8_8), .in1(tmp01_9_8), .out(tmp02_4_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000711(.in0(tmp01_10_8), .in1(tmp01_11_8), .out(tmp02_5_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000712(.in0(tmp01_12_8), .in1(tmp01_13_8), .out(tmp02_6_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000713(.in0(tmp01_14_8), .in1(tmp01_15_8), .out(tmp02_7_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000714(.in0(tmp01_16_8), .in1(tmp01_17_8), .out(tmp02_8_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000715(.in0(tmp01_18_8), .in1(tmp01_19_8), .out(tmp02_9_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000716(.in0(tmp01_20_8), .in1(tmp01_21_8), .out(tmp02_10_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000717(.in0(tmp01_22_8), .in1(tmp01_23_8), .out(tmp02_11_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000718(.in0(tmp01_24_8), .in1(tmp01_25_8), .out(tmp02_12_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000719(.in0(tmp01_26_8), .in1(tmp01_27_8), .out(tmp02_13_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000720(.in0(tmp01_28_8), .in1(tmp01_29_8), .out(tmp02_14_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000721(.in0(tmp01_30_8), .in1(tmp01_31_8), .out(tmp02_15_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000722(.in0(tmp01_32_8), .in1(tmp01_33_8), .out(tmp02_16_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000723(.in0(tmp01_34_8), .in1(tmp01_35_8), .out(tmp02_17_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000724(.in0(tmp01_36_8), .in1(tmp01_37_8), .out(tmp02_18_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000725(.in0(tmp01_38_8), .in1(tmp01_39_8), .out(tmp02_19_8));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000726(.in0(tmp01_40_8), .in1(tmp01_41_8), .out(tmp02_20_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000727(.in0(tmp02_0_8), .in1(tmp02_1_8), .out(tmp03_0_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000728(.in0(tmp02_2_8), .in1(tmp02_3_8), .out(tmp03_1_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000729(.in0(tmp02_4_8), .in1(tmp02_5_8), .out(tmp03_2_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000730(.in0(tmp02_6_8), .in1(tmp02_7_8), .out(tmp03_3_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000731(.in0(tmp02_8_8), .in1(tmp02_9_8), .out(tmp03_4_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000732(.in0(tmp02_10_8), .in1(tmp02_11_8), .out(tmp03_5_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000733(.in0(tmp02_12_8), .in1(tmp02_13_8), .out(tmp03_6_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000734(.in0(tmp02_14_8), .in1(tmp02_15_8), .out(tmp03_7_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000735(.in0(tmp02_16_8), .in1(tmp02_17_8), .out(tmp03_8_8));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000736(.in0(tmp02_18_8), .in1(tmp02_19_8), .out(tmp03_9_8));
	assign tmp03_10_8 = $signed(tmp02_20_8);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000737(.in0(tmp03_0_8), .in1(tmp03_1_8), .out(tmp04_0_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000738(.in0(tmp03_2_8), .in1(tmp03_3_8), .out(tmp04_1_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000739(.in0(tmp03_4_8), .in1(tmp03_5_8), .out(tmp04_2_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000740(.in0(tmp03_6_8), .in1(tmp03_7_8), .out(tmp04_3_8));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000741(.in0(tmp03_8_8), .in1(tmp03_9_8), .out(tmp04_4_8));
	assign tmp04_5_8 = $signed(tmp03_10_8);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000742(.in0(tmp04_0_8), .in1(tmp04_1_8), .out(tmp05_0_8));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000743(.in0(tmp04_2_8), .in1(tmp04_3_8), .out(tmp05_1_8));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000744(.in0(tmp04_4_8), .in1(tmp04_5_8), .out(tmp05_2_8));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000745(.in0(tmp05_0_8), .in1(tmp05_1_8), .out(tmp06_0_8));
	assign tmp06_1_8 = $signed(tmp05_2_8);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000746(.in0(tmp06_0_8), .in1(tmp06_1_8), .out(tmp07_0_8));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000747(.in0(tmp00_0_9), .in1(tmp00_1_9), .out(tmp01_0_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000748(.in0(tmp00_2_9), .in1(tmp00_3_9), .out(tmp01_1_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000749(.in0(tmp00_4_9), .in1(tmp00_5_9), .out(tmp01_2_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000750(.in0(tmp00_6_9), .in1(tmp00_7_9), .out(tmp01_3_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000751(.in0(tmp00_8_9), .in1(tmp00_9_9), .out(tmp01_4_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000752(.in0(tmp00_10_9), .in1(tmp00_11_9), .out(tmp01_5_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000753(.in0(tmp00_12_9), .in1(tmp00_13_9), .out(tmp01_6_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000754(.in0(tmp00_14_9), .in1(tmp00_15_9), .out(tmp01_7_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000755(.in0(tmp00_16_9), .in1(tmp00_17_9), .out(tmp01_8_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000756(.in0(tmp00_18_9), .in1(tmp00_19_9), .out(tmp01_9_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000757(.in0(tmp00_20_9), .in1(tmp00_21_9), .out(tmp01_10_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000758(.in0(tmp00_22_9), .in1(tmp00_23_9), .out(tmp01_11_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000759(.in0(tmp00_24_9), .in1(tmp00_25_9), .out(tmp01_12_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000760(.in0(tmp00_26_9), .in1(tmp00_27_9), .out(tmp01_13_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000761(.in0(tmp00_28_9), .in1(tmp00_29_9), .out(tmp01_14_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000762(.in0(tmp00_30_9), .in1(tmp00_31_9), .out(tmp01_15_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000763(.in0(tmp00_32_9), .in1(tmp00_33_9), .out(tmp01_16_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000764(.in0(tmp00_34_9), .in1(tmp00_35_9), .out(tmp01_17_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000765(.in0(tmp00_36_9), .in1(tmp00_37_9), .out(tmp01_18_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000766(.in0(tmp00_38_9), .in1(tmp00_39_9), .out(tmp01_19_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000767(.in0(tmp00_40_9), .in1(tmp00_41_9), .out(tmp01_20_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000768(.in0(tmp00_42_9), .in1(tmp00_43_9), .out(tmp01_21_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000769(.in0(tmp00_44_9), .in1(tmp00_45_9), .out(tmp01_22_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000770(.in0(tmp00_46_9), .in1(tmp00_47_9), .out(tmp01_23_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000771(.in0(tmp00_48_9), .in1(tmp00_49_9), .out(tmp01_24_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000772(.in0(tmp00_50_9), .in1(tmp00_51_9), .out(tmp01_25_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000773(.in0(tmp00_52_9), .in1(tmp00_53_9), .out(tmp01_26_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000774(.in0(tmp00_54_9), .in1(tmp00_55_9), .out(tmp01_27_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000775(.in0(tmp00_56_9), .in1(tmp00_57_9), .out(tmp01_28_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000776(.in0(tmp00_58_9), .in1(tmp00_59_9), .out(tmp01_29_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000777(.in0(tmp00_60_9), .in1(tmp00_61_9), .out(tmp01_30_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000778(.in0(tmp00_62_9), .in1(tmp00_63_9), .out(tmp01_31_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000779(.in0(tmp00_64_9), .in1(tmp00_65_9), .out(tmp01_32_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000780(.in0(tmp00_66_9), .in1(tmp00_67_9), .out(tmp01_33_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000781(.in0(tmp00_68_9), .in1(tmp00_69_9), .out(tmp01_34_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000782(.in0(tmp00_70_9), .in1(tmp00_71_9), .out(tmp01_35_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000783(.in0(tmp00_72_9), .in1(tmp00_73_9), .out(tmp01_36_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000784(.in0(tmp00_74_9), .in1(tmp00_75_9), .out(tmp01_37_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000785(.in0(tmp00_76_9), .in1(tmp00_77_9), .out(tmp01_38_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000786(.in0(tmp00_78_9), .in1(tmp00_79_9), .out(tmp01_39_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000787(.in0(tmp00_80_9), .in1(tmp00_81_9), .out(tmp01_40_9));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000788(.in0(tmp00_82_9), .in1(tmp00_83_9), .out(tmp01_41_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000789(.in0(tmp01_0_9), .in1(tmp01_1_9), .out(tmp02_0_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000790(.in0(tmp01_2_9), .in1(tmp01_3_9), .out(tmp02_1_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000791(.in0(tmp01_4_9), .in1(tmp01_5_9), .out(tmp02_2_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000792(.in0(tmp01_6_9), .in1(tmp01_7_9), .out(tmp02_3_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000793(.in0(tmp01_8_9), .in1(tmp01_9_9), .out(tmp02_4_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000794(.in0(tmp01_10_9), .in1(tmp01_11_9), .out(tmp02_5_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000795(.in0(tmp01_12_9), .in1(tmp01_13_9), .out(tmp02_6_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000796(.in0(tmp01_14_9), .in1(tmp01_15_9), .out(tmp02_7_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000797(.in0(tmp01_16_9), .in1(tmp01_17_9), .out(tmp02_8_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000798(.in0(tmp01_18_9), .in1(tmp01_19_9), .out(tmp02_9_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000799(.in0(tmp01_20_9), .in1(tmp01_21_9), .out(tmp02_10_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000800(.in0(tmp01_22_9), .in1(tmp01_23_9), .out(tmp02_11_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000801(.in0(tmp01_24_9), .in1(tmp01_25_9), .out(tmp02_12_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000802(.in0(tmp01_26_9), .in1(tmp01_27_9), .out(tmp02_13_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000803(.in0(tmp01_28_9), .in1(tmp01_29_9), .out(tmp02_14_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000804(.in0(tmp01_30_9), .in1(tmp01_31_9), .out(tmp02_15_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000805(.in0(tmp01_32_9), .in1(tmp01_33_9), .out(tmp02_16_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000806(.in0(tmp01_34_9), .in1(tmp01_35_9), .out(tmp02_17_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000807(.in0(tmp01_36_9), .in1(tmp01_37_9), .out(tmp02_18_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000808(.in0(tmp01_38_9), .in1(tmp01_39_9), .out(tmp02_19_9));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000809(.in0(tmp01_40_9), .in1(tmp01_41_9), .out(tmp02_20_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000810(.in0(tmp02_0_9), .in1(tmp02_1_9), .out(tmp03_0_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000811(.in0(tmp02_2_9), .in1(tmp02_3_9), .out(tmp03_1_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000812(.in0(tmp02_4_9), .in1(tmp02_5_9), .out(tmp03_2_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000813(.in0(tmp02_6_9), .in1(tmp02_7_9), .out(tmp03_3_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000814(.in0(tmp02_8_9), .in1(tmp02_9_9), .out(tmp03_4_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000815(.in0(tmp02_10_9), .in1(tmp02_11_9), .out(tmp03_5_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000816(.in0(tmp02_12_9), .in1(tmp02_13_9), .out(tmp03_6_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000817(.in0(tmp02_14_9), .in1(tmp02_15_9), .out(tmp03_7_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000818(.in0(tmp02_16_9), .in1(tmp02_17_9), .out(tmp03_8_9));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000819(.in0(tmp02_18_9), .in1(tmp02_19_9), .out(tmp03_9_9));
	assign tmp03_10_9 = $signed(tmp02_20_9);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000820(.in0(tmp03_0_9), .in1(tmp03_1_9), .out(tmp04_0_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000821(.in0(tmp03_2_9), .in1(tmp03_3_9), .out(tmp04_1_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000822(.in0(tmp03_4_9), .in1(tmp03_5_9), .out(tmp04_2_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000823(.in0(tmp03_6_9), .in1(tmp03_7_9), .out(tmp04_3_9));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000824(.in0(tmp03_8_9), .in1(tmp03_9_9), .out(tmp04_4_9));
	assign tmp04_5_9 = $signed(tmp03_10_9);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000825(.in0(tmp04_0_9), .in1(tmp04_1_9), .out(tmp05_0_9));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000826(.in0(tmp04_2_9), .in1(tmp04_3_9), .out(tmp05_1_9));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000827(.in0(tmp04_4_9), .in1(tmp04_5_9), .out(tmp05_2_9));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000828(.in0(tmp05_0_9), .in1(tmp05_1_9), .out(tmp06_0_9));
	assign tmp06_1_9 = $signed(tmp05_2_9);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000829(.in0(tmp06_0_9), .in1(tmp06_1_9), .out(tmp07_0_9));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU000(.a(tmp07_0_0), .b(23'h0), .sel(tmp07_0_0[WIDTH*2+$clog2(IN)-1]), .out(z_0));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU001(.a(tmp07_0_1), .b(23'h0), .sel(tmp07_0_1[WIDTH*2+$clog2(IN)-1]), .out(z_1));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU002(.a(tmp07_0_2), .b(23'h0), .sel(tmp07_0_2[WIDTH*2+$clog2(IN)-1]), .out(z_2));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU003(.a(tmp07_0_3), .b(23'h0), .sel(tmp07_0_3[WIDTH*2+$clog2(IN)-1]), .out(z_3));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU004(.a(tmp07_0_4), .b(23'h0), .sel(tmp07_0_4[WIDTH*2+$clog2(IN)-1]), .out(z_4));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU005(.a(tmp07_0_5), .b(23'h0), .sel(tmp07_0_5[WIDTH*2+$clog2(IN)-1]), .out(z_5));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU006(.a(tmp07_0_6), .b(23'h0), .sel(tmp07_0_6[WIDTH*2+$clog2(IN)-1]), .out(z_6));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU007(.a(tmp07_0_7), .b(23'h0), .sel(tmp07_0_7[WIDTH*2+$clog2(IN)-1]), .out(z_7));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU008(.a(tmp07_0_8), .b(23'h0), .sel(tmp07_0_8[WIDTH*2+$clog2(IN)-1]), .out(z_8));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU009(.a(tmp07_0_9), .b(23'h0), .sel(tmp07_0_9[WIDTH*2+$clog2(IN)-1]), .out(z_9));
endmodule

