module layer
	#(parameter WIDTH = 8)
	(x, z);
	localparam IN = 400;
	input [WIDTH-1:0] x[0:IN-1];
	output [WIDTH*2+$clog2(195)-1:0] z;
	wire [WIDTH*2-1+0:0] tmp00[0:194];
	wire [WIDTH*2-1+1:0] tmp01[0:97];
	wire [WIDTH*2-1+2:0] tmp02[0:48];
	wire [WIDTH*2-1+3:0] tmp03[0:24];
	wire [WIDTH*2-1+4:0] tmp04[0:12];
	wire [WIDTH*2-1+5:0] tmp05[0:6];
	wire [WIDTH*2-1+6:0] tmp06[0:3];
	wire [WIDTH*2-1+7:0] tmp07[0:1];
	wire [WIDTH*2-1+8:0] tmp08[0:0];
	booth_0010 #(.WIDTH(WIDTH)) mul00(.x(x[1]), .z(tmp00[0]));
	booth_0004 #(.WIDTH(WIDTH)) mul01(.x(x[2]), .z(tmp00[1]));
	booth__004 #(.WIDTH(WIDTH)) mul02(.x(x[5]), .z(tmp00[2]));
	booth__004 #(.WIDTH(WIDTH)) mul03(.x(x[6]), .z(tmp00[3]));
	booth_0004 #(.WIDTH(WIDTH)) mul04(.x(x[7]), .z(tmp00[4]));
	booth__008 #(.WIDTH(WIDTH)) mul05(.x(x[9]), .z(tmp00[5]));
	booth__012 #(.WIDTH(WIDTH)) mul06(.x(x[10]), .z(tmp00[6]));
	booth__006 #(.WIDTH(WIDTH)) mul07(.x(x[11]), .z(tmp00[7]));
	booth_0004 #(.WIDTH(WIDTH)) mul08(.x(x[22]), .z(tmp00[8]));
	booth_0012 #(.WIDTH(WIDTH)) mul09(.x(x[23]), .z(tmp00[9]));
	booth_0004 #(.WIDTH(WIDTH)) mul10(.x(x[25]), .z(tmp00[10]));
	booth_0012 #(.WIDTH(WIDTH)) mul11(.x(x[26]), .z(tmp00[11]));
	booth_0020 #(.WIDTH(WIDTH)) mul12(.x(x[27]), .z(tmp00[12]));
	booth_0024 #(.WIDTH(WIDTH)) mul13(.x(x[29]), .z(tmp00[13]));
	booth__020 #(.WIDTH(WIDTH)) mul14(.x(x[31]), .z(tmp00[14]));
	booth__016 #(.WIDTH(WIDTH)) mul15(.x(x[32]), .z(tmp00[15]));
	booth_0004 #(.WIDTH(WIDTH)) mul16(.x(x[34]), .z(tmp00[16]));
	booth_0012 #(.WIDTH(WIDTH)) mul17(.x(x[40]), .z(tmp00[17]));
	booth__012 #(.WIDTH(WIDTH)) mul18(.x(x[44]), .z(tmp00[18]));
	booth__032 #(.WIDTH(WIDTH)) mul19(.x(x[49]), .z(tmp00[19]));
	booth_0012 #(.WIDTH(WIDTH)) mul20(.x(x[50]), .z(tmp00[20]));
	booth_0008 #(.WIDTH(WIDTH)) mul21(.x(x[51]), .z(tmp00[21]));
	booth_0008 #(.WIDTH(WIDTH)) mul22(.x(x[53]), .z(tmp00[22]));
	booth_0004 #(.WIDTH(WIDTH)) mul23(.x(x[54]), .z(tmp00[23]));
	booth__016 #(.WIDTH(WIDTH)) mul24(.x(x[55]), .z(tmp00[24]));
	booth_0004 #(.WIDTH(WIDTH)) mul25(.x(x[56]), .z(tmp00[25]));
	booth__012 #(.WIDTH(WIDTH)) mul26(.x(x[58]), .z(tmp00[26]));
	booth_0004 #(.WIDTH(WIDTH)) mul27(.x(x[59]), .z(tmp00[27]));
	booth__018 #(.WIDTH(WIDTH)) mul28(.x(x[60]), .z(tmp00[28]));
	booth_0004 #(.WIDTH(WIDTH)) mul29(.x(x[64]), .z(tmp00[29]));
	booth__008 #(.WIDTH(WIDTH)) mul30(.x(x[65]), .z(tmp00[30]));
	booth_0004 #(.WIDTH(WIDTH)) mul31(.x(x[67]), .z(tmp00[31]));
	booth_0005 #(.WIDTH(WIDTH)) mul32(.x(x[68]), .z(tmp00[32]));
	booth_0005 #(.WIDTH(WIDTH)) mul33(.x(x[69]), .z(tmp00[33]));
	booth_0005 #(.WIDTH(WIDTH)) mul34(.x(x[70]), .z(tmp00[34]));
	booth__028 #(.WIDTH(WIDTH)) mul35(.x(x[71]), .z(tmp00[35]));
	booth__008 #(.WIDTH(WIDTH)) mul36(.x(x[74]), .z(tmp00[36]));
	booth_0010 #(.WIDTH(WIDTH)) mul37(.x(x[75]), .z(tmp00[37]));
	booth__030 #(.WIDTH(WIDTH)) mul38(.x(x[77]), .z(tmp00[38]));
	booth__030 #(.WIDTH(WIDTH)) mul39(.x(x[79]), .z(tmp00[39]));
	booth_0010 #(.WIDTH(WIDTH)) mul40(.x(x[80]), .z(tmp00[40]));
	booth_0004 #(.WIDTH(WIDTH)) mul41(.x(x[84]), .z(tmp00[41]));
	booth_0014 #(.WIDTH(WIDTH)) mul42(.x(x[86]), .z(tmp00[42]));
	booth_0020 #(.WIDTH(WIDTH)) mul43(.x(x[87]), .z(tmp00[43]));
	booth_0008 #(.WIDTH(WIDTH)) mul44(.x(x[88]), .z(tmp00[44]));
	booth_0018 #(.WIDTH(WIDTH)) mul45(.x(x[89]), .z(tmp00[45]));
	booth_0004 #(.WIDTH(WIDTH)) mul46(.x(x[90]), .z(tmp00[46]));
	booth_0012 #(.WIDTH(WIDTH)) mul47(.x(x[91]), .z(tmp00[47]));
	booth_0012 #(.WIDTH(WIDTH)) mul48(.x(x[92]), .z(tmp00[48]));
	booth_0010 #(.WIDTH(WIDTH)) mul49(.x(x[94]), .z(tmp00[49]));
	booth_0008 #(.WIDTH(WIDTH)) mul50(.x(x[96]), .z(tmp00[50]));
	booth__016 #(.WIDTH(WIDTH)) mul51(.x(x[99]), .z(tmp00[51]));
	booth_0005 #(.WIDTH(WIDTH)) mul52(.x(x[100]), .z(tmp00[52]));
	booth__008 #(.WIDTH(WIDTH)) mul53(.x(x[101]), .z(tmp00[53]));
	booth__012 #(.WIDTH(WIDTH)) mul54(.x(x[106]), .z(tmp00[54]));
	booth__012 #(.WIDTH(WIDTH)) mul55(.x(x[109]), .z(tmp00[55]));
	booth__008 #(.WIDTH(WIDTH)) mul56(.x(x[111]), .z(tmp00[56]));
	booth__010 #(.WIDTH(WIDTH)) mul57(.x(x[114]), .z(tmp00[57]));
	booth__016 #(.WIDTH(WIDTH)) mul58(.x(x[116]), .z(tmp00[58]));
	booth__016 #(.WIDTH(WIDTH)) mul59(.x(x[117]), .z(tmp00[59]));
	booth_0004 #(.WIDTH(WIDTH)) mul60(.x(x[118]), .z(tmp00[60]));
	booth__012 #(.WIDTH(WIDTH)) mul61(.x(x[121]), .z(tmp00[61]));
	booth_0002 #(.WIDTH(WIDTH)) mul62(.x(x[123]), .z(tmp00[62]));
	booth__030 #(.WIDTH(WIDTH)) mul63(.x(x[125]), .z(tmp00[63]));
	booth__012 #(.WIDTH(WIDTH)) mul64(.x(x[126]), .z(tmp00[64]));
	booth__012 #(.WIDTH(WIDTH)) mul65(.x(x[130]), .z(tmp00[65]));
	booth_0004 #(.WIDTH(WIDTH)) mul66(.x(x[131]), .z(tmp00[66]));
	booth_0002 #(.WIDTH(WIDTH)) mul67(.x(x[132]), .z(tmp00[67]));
	booth_0012 #(.WIDTH(WIDTH)) mul68(.x(x[133]), .z(tmp00[68]));
	booth_0020 #(.WIDTH(WIDTH)) mul69(.x(x[134]), .z(tmp00[69]));
	booth__020 #(.WIDTH(WIDTH)) mul70(.x(x[135]), .z(tmp00[70]));
	booth_0002 #(.WIDTH(WIDTH)) mul71(.x(x[136]), .z(tmp00[71]));
	booth_0005 #(.WIDTH(WIDTH)) mul72(.x(x[137]), .z(tmp00[72]));
	booth_0012 #(.WIDTH(WIDTH)) mul73(.x(x[138]), .z(tmp00[73]));
	booth_0012 #(.WIDTH(WIDTH)) mul74(.x(x[139]), .z(tmp00[74]));
	booth__022 #(.WIDTH(WIDTH)) mul75(.x(x[140]), .z(tmp00[75]));
	booth_0004 #(.WIDTH(WIDTH)) mul76(.x(x[141]), .z(tmp00[76]));
	booth_0018 #(.WIDTH(WIDTH)) mul77(.x(x[143]), .z(tmp00[77]));
	booth__036 #(.WIDTH(WIDTH)) mul78(.x(x[145]), .z(tmp00[78]));
	booth__012 #(.WIDTH(WIDTH)) mul79(.x(x[146]), .z(tmp00[79]));
	booth_0014 #(.WIDTH(WIDTH)) mul80(.x(x[148]), .z(tmp00[80]));
	booth_0012 #(.WIDTH(WIDTH)) mul81(.x(x[150]), .z(tmp00[81]));
	booth_0012 #(.WIDTH(WIDTH)) mul82(.x(x[153]), .z(tmp00[82]));
	booth_0004 #(.WIDTH(WIDTH)) mul83(.x(x[154]), .z(tmp00[83]));
	booth_0004 #(.WIDTH(WIDTH)) mul84(.x(x[156]), .z(tmp00[84]));
	booth_0002 #(.WIDTH(WIDTH)) mul85(.x(x[157]), .z(tmp00[85]));
	booth__008 #(.WIDTH(WIDTH)) mul86(.x(x[159]), .z(tmp00[86]));
	booth_0005 #(.WIDTH(WIDTH)) mul87(.x(x[162]), .z(tmp00[87]));
	booth__010 #(.WIDTH(WIDTH)) mul88(.x(x[164]), .z(tmp00[88]));
	booth_0010 #(.WIDTH(WIDTH)) mul89(.x(x[165]), .z(tmp00[89]));
	booth_0010 #(.WIDTH(WIDTH)) mul90(.x(x[167]), .z(tmp00[90]));
	booth_0008 #(.WIDTH(WIDTH)) mul91(.x(x[172]), .z(tmp00[91]));
	booth_0010 #(.WIDTH(WIDTH)) mul92(.x(x[173]), .z(tmp00[92]));
	booth_0036 #(.WIDTH(WIDTH)) mul93(.x(x[175]), .z(tmp00[93]));
	booth_0016 #(.WIDTH(WIDTH)) mul94(.x(x[176]), .z(tmp00[94]));
	booth_0012 #(.WIDTH(WIDTH)) mul95(.x(x[177]), .z(tmp00[95]));
	booth_0002 #(.WIDTH(WIDTH)) mul96(.x(x[180]), .z(tmp00[96]));
	booth__016 #(.WIDTH(WIDTH)) mul97(.x(x[181]), .z(tmp00[97]));
	booth__012 #(.WIDTH(WIDTH)) mul98(.x(x[183]), .z(tmp00[98]));
	booth__012 #(.WIDTH(WIDTH)) mul99(.x(x[184]), .z(tmp00[99]));
	booth__014 #(.WIDTH(WIDTH)) mul100(.x(x[186]), .z(tmp00[100]));
	booth__012 #(.WIDTH(WIDTH)) mul101(.x(x[187]), .z(tmp00[101]));
	booth__016 #(.WIDTH(WIDTH)) mul102(.x(x[188]), .z(tmp00[102]));
	booth__020 #(.WIDTH(WIDTH)) mul103(.x(x[189]), .z(tmp00[103]));
	booth_0006 #(.WIDTH(WIDTH)) mul104(.x(x[191]), .z(tmp00[104]));
	booth__008 #(.WIDTH(WIDTH)) mul105(.x(x[193]), .z(tmp00[105]));
	booth_0016 #(.WIDTH(WIDTH)) mul106(.x(x[196]), .z(tmp00[106]));
	booth_0004 #(.WIDTH(WIDTH)) mul107(.x(x[197]), .z(tmp00[107]));
	booth_0004 #(.WIDTH(WIDTH)) mul108(.x(x[199]), .z(tmp00[108]));
	booth_0002 #(.WIDTH(WIDTH)) mul109(.x(x[200]), .z(tmp00[109]));
	booth__012 #(.WIDTH(WIDTH)) mul110(.x(x[202]), .z(tmp00[110]));
	booth_0004 #(.WIDTH(WIDTH)) mul111(.x(x[204]), .z(tmp00[111]));
	booth__012 #(.WIDTH(WIDTH)) mul112(.x(x[206]), .z(tmp00[112]));
	booth_0004 #(.WIDTH(WIDTH)) mul113(.x(x[207]), .z(tmp00[113]));
	booth__016 #(.WIDTH(WIDTH)) mul114(.x(x[209]), .z(tmp00[114]));
	booth__016 #(.WIDTH(WIDTH)) mul115(.x(x[213]), .z(tmp00[115]));
	booth__012 #(.WIDTH(WIDTH)) mul116(.x(x[214]), .z(tmp00[116]));
	booth__020 #(.WIDTH(WIDTH)) mul117(.x(x[215]), .z(tmp00[117]));
	booth__012 #(.WIDTH(WIDTH)) mul118(.x(x[216]), .z(tmp00[118]));
	booth_0002 #(.WIDTH(WIDTH)) mul119(.x(x[218]), .z(tmp00[119]));
	booth__018 #(.WIDTH(WIDTH)) mul120(.x(x[219]), .z(tmp00[120]));
	booth_0002 #(.WIDTH(WIDTH)) mul121(.x(x[223]), .z(tmp00[121]));
	booth__008 #(.WIDTH(WIDTH)) mul122(.x(x[227]), .z(tmp00[122]));
	booth_0012 #(.WIDTH(WIDTH)) mul123(.x(x[228]), .z(tmp00[123]));
	booth_0008 #(.WIDTH(WIDTH)) mul124(.x(x[233]), .z(tmp00[124]));
	booth_0012 #(.WIDTH(WIDTH)) mul125(.x(x[234]), .z(tmp00[125]));
	booth__004 #(.WIDTH(WIDTH)) mul126(.x(x[237]), .z(tmp00[126]));
	booth__012 #(.WIDTH(WIDTH)) mul127(.x(x[240]), .z(tmp00[127]));
	booth_0008 #(.WIDTH(WIDTH)) mul128(.x(x[243]), .z(tmp00[128]));
	booth_0010 #(.WIDTH(WIDTH)) mul129(.x(x[244]), .z(tmp00[129]));
	booth_0004 #(.WIDTH(WIDTH)) mul130(.x(x[247]), .z(tmp00[130]));
	booth_0025 #(.WIDTH(WIDTH)) mul131(.x(x[248]), .z(tmp00[131]));
	booth_0004 #(.WIDTH(WIDTH)) mul132(.x(x[250]), .z(tmp00[132]));
	booth__006 #(.WIDTH(WIDTH)) mul133(.x(x[252]), .z(tmp00[133]));
	booth__008 #(.WIDTH(WIDTH)) mul134(.x(x[269]), .z(tmp00[134]));
	booth__008 #(.WIDTH(WIDTH)) mul135(.x(x[274]), .z(tmp00[135]));
	booth_0021 #(.WIDTH(WIDTH)) mul136(.x(x[275]), .z(tmp00[136]));
	booth_0012 #(.WIDTH(WIDTH)) mul137(.x(x[277]), .z(tmp00[137]));
	booth_0005 #(.WIDTH(WIDTH)) mul138(.x(x[278]), .z(tmp00[138]));
	booth_0004 #(.WIDTH(WIDTH)) mul139(.x(x[281]), .z(tmp00[139]));
	booth_0004 #(.WIDTH(WIDTH)) mul140(.x(x[282]), .z(tmp00[140]));
	booth_0008 #(.WIDTH(WIDTH)) mul141(.x(x[285]), .z(tmp00[141]));
	booth_0004 #(.WIDTH(WIDTH)) mul142(.x(x[286]), .z(tmp00[142]));
	booth_0004 #(.WIDTH(WIDTH)) mul143(.x(x[287]), .z(tmp00[143]));
	booth_0012 #(.WIDTH(WIDTH)) mul144(.x(x[290]), .z(tmp00[144]));
	booth_0008 #(.WIDTH(WIDTH)) mul145(.x(x[292]), .z(tmp00[145]));
	booth_0016 #(.WIDTH(WIDTH)) mul146(.x(x[293]), .z(tmp00[146]));
	booth__022 #(.WIDTH(WIDTH)) mul147(.x(x[295]), .z(tmp00[147]));
	booth__018 #(.WIDTH(WIDTH)) mul148(.x(x[296]), .z(tmp00[148]));
	booth__010 #(.WIDTH(WIDTH)) mul149(.x(x[297]), .z(tmp00[149]));
	booth_0012 #(.WIDTH(WIDTH)) mul150(.x(x[299]), .z(tmp00[150]));
	booth__012 #(.WIDTH(WIDTH)) mul151(.x(x[303]), .z(tmp00[151]));
	booth__018 #(.WIDTH(WIDTH)) mul152(.x(x[305]), .z(tmp00[152]));
	booth_0004 #(.WIDTH(WIDTH)) mul153(.x(x[307]), .z(tmp00[153]));
	booth_0004 #(.WIDTH(WIDTH)) mul154(.x(x[308]), .z(tmp00[154]));
	booth_0008 #(.WIDTH(WIDTH)) mul155(.x(x[312]), .z(tmp00[155]));
	booth_0020 #(.WIDTH(WIDTH)) mul156(.x(x[318]), .z(tmp00[156]));
	booth_0004 #(.WIDTH(WIDTH)) mul157(.x(x[319]), .z(tmp00[157]));
	booth_0004 #(.WIDTH(WIDTH)) mul158(.x(x[321]), .z(tmp00[158]));
	booth_0005 #(.WIDTH(WIDTH)) mul159(.x(x[322]), .z(tmp00[159]));
	booth_0004 #(.WIDTH(WIDTH)) mul160(.x(x[330]), .z(tmp00[160]));
	booth_0010 #(.WIDTH(WIDTH)) mul161(.x(x[332]), .z(tmp00[161]));
	booth_0008 #(.WIDTH(WIDTH)) mul162(.x(x[333]), .z(tmp00[162]));
	booth__008 #(.WIDTH(WIDTH)) mul163(.x(x[334]), .z(tmp00[163]));
	booth__018 #(.WIDTH(WIDTH)) mul164(.x(x[335]), .z(tmp00[164]));
	booth__016 #(.WIDTH(WIDTH)) mul165(.x(x[336]), .z(tmp00[165]));
	booth__020 #(.WIDTH(WIDTH)) mul166(.x(x[339]), .z(tmp00[166]));
	booth__008 #(.WIDTH(WIDTH)) mul167(.x(x[343]), .z(tmp00[167]));
	booth__016 #(.WIDTH(WIDTH)) mul168(.x(x[344]), .z(tmp00[168]));
	booth__012 #(.WIDTH(WIDTH)) mul169(.x(x[346]), .z(tmp00[169]));
	booth__010 #(.WIDTH(WIDTH)) mul170(.x(x[350]), .z(tmp00[170]));
	booth_0010 #(.WIDTH(WIDTH)) mul171(.x(x[352]), .z(tmp00[171]));
	booth_0016 #(.WIDTH(WIDTH)) mul172(.x(x[357]), .z(tmp00[172]));
	booth_0004 #(.WIDTH(WIDTH)) mul173(.x(x[358]), .z(tmp00[173]));
	booth__004 #(.WIDTH(WIDTH)) mul174(.x(x[364]), .z(tmp00[174]));
	booth_0002 #(.WIDTH(WIDTH)) mul175(.x(x[371]), .z(tmp00[175]));
	booth__012 #(.WIDTH(WIDTH)) mul176(.x(x[375]), .z(tmp00[176]));
	booth_0002 #(.WIDTH(WIDTH)) mul177(.x(x[376]), .z(tmp00[177]));
	booth__020 #(.WIDTH(WIDTH)) mul178(.x(x[377]), .z(tmp00[178]));
	booth__016 #(.WIDTH(WIDTH)) mul179(.x(x[378]), .z(tmp00[179]));
	booth__024 #(.WIDTH(WIDTH)) mul180(.x(x[379]), .z(tmp00[180]));
	booth_0008 #(.WIDTH(WIDTH)) mul181(.x(x[381]), .z(tmp00[181]));
	booth_0012 #(.WIDTH(WIDTH)) mul182(.x(x[382]), .z(tmp00[182]));
	booth_0008 #(.WIDTH(WIDTH)) mul183(.x(x[383]), .z(tmp00[183]));
	booth__012 #(.WIDTH(WIDTH)) mul184(.x(x[384]), .z(tmp00[184]));
	booth__020 #(.WIDTH(WIDTH)) mul185(.x(x[385]), .z(tmp00[185]));
	booth_0010 #(.WIDTH(WIDTH)) mul186(.x(x[387]), .z(tmp00[186]));
	booth_0008 #(.WIDTH(WIDTH)) mul187(.x(x[388]), .z(tmp00[187]));
	booth__018 #(.WIDTH(WIDTH)) mul188(.x(x[390]), .z(tmp00[188]));
	booth__008 #(.WIDTH(WIDTH)) mul189(.x(x[391]), .z(tmp00[189]));
	booth_0012 #(.WIDTH(WIDTH)) mul190(.x(x[392]), .z(tmp00[190]));
	booth_0004 #(.WIDTH(WIDTH)) mul191(.x(x[393]), .z(tmp00[191]));
	booth__020 #(.WIDTH(WIDTH)) mul192(.x(x[396]), .z(tmp00[192]));
	booth_0004 #(.WIDTH(WIDTH)) mul193(.x(x[397]), .z(tmp00[193]));
	booth_0010 #(.WIDTH(WIDTH)) mul194(.x(x[398]), .z(tmp00[194]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000000(.in0(tmp00[0]), .in1(tmp00[1]), .out(tmp01[0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000001(.in0(tmp00[2]), .in1(tmp00[3]), .out(tmp01[1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000002(.in0(tmp00[4]), .in1(tmp00[5]), .out(tmp01[2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000003(.in0(tmp00[6]), .in1(tmp00[7]), .out(tmp01[3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000004(.in0(tmp00[8]), .in1(tmp00[9]), .out(tmp01[4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000005(.in0(tmp00[10]), .in1(tmp00[11]), .out(tmp01[5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000006(.in0(tmp00[12]), .in1(tmp00[13]), .out(tmp01[6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000007(.in0(tmp00[14]), .in1(tmp00[15]), .out(tmp01[7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000008(.in0(tmp00[16]), .in1(tmp00[17]), .out(tmp01[8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000009(.in0(tmp00[18]), .in1(tmp00[19]), .out(tmp01[9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000010(.in0(tmp00[20]), .in1(tmp00[21]), .out(tmp01[10]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000011(.in0(tmp00[22]), .in1(tmp00[23]), .out(tmp01[11]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000012(.in0(tmp00[24]), .in1(tmp00[25]), .out(tmp01[12]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000013(.in0(tmp00[26]), .in1(tmp00[27]), .out(tmp01[13]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000014(.in0(tmp00[28]), .in1(tmp00[29]), .out(tmp01[14]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000015(.in0(tmp00[30]), .in1(tmp00[31]), .out(tmp01[15]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000016(.in0(tmp00[32]), .in1(tmp00[33]), .out(tmp01[16]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000017(.in0(tmp00[34]), .in1(tmp00[35]), .out(tmp01[17]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000018(.in0(tmp00[36]), .in1(tmp00[37]), .out(tmp01[18]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000019(.in0(tmp00[38]), .in1(tmp00[39]), .out(tmp01[19]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000020(.in0(tmp00[40]), .in1(tmp00[41]), .out(tmp01[20]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000021(.in0(tmp00[42]), .in1(tmp00[43]), .out(tmp01[21]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000022(.in0(tmp00[44]), .in1(tmp00[45]), .out(tmp01[22]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000023(.in0(tmp00[46]), .in1(tmp00[47]), .out(tmp01[23]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000024(.in0(tmp00[48]), .in1(tmp00[49]), .out(tmp01[24]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000025(.in0(tmp00[50]), .in1(tmp00[51]), .out(tmp01[25]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000026(.in0(tmp00[52]), .in1(tmp00[53]), .out(tmp01[26]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000027(.in0(tmp00[54]), .in1(tmp00[55]), .out(tmp01[27]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000028(.in0(tmp00[56]), .in1(tmp00[57]), .out(tmp01[28]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000029(.in0(tmp00[58]), .in1(tmp00[59]), .out(tmp01[29]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000030(.in0(tmp00[60]), .in1(tmp00[61]), .out(tmp01[30]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000031(.in0(tmp00[62]), .in1(tmp00[63]), .out(tmp01[31]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000032(.in0(tmp00[64]), .in1(tmp00[65]), .out(tmp01[32]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000033(.in0(tmp00[66]), .in1(tmp00[67]), .out(tmp01[33]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000034(.in0(tmp00[68]), .in1(tmp00[69]), .out(tmp01[34]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000035(.in0(tmp00[70]), .in1(tmp00[71]), .out(tmp01[35]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000036(.in0(tmp00[72]), .in1(tmp00[73]), .out(tmp01[36]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000037(.in0(tmp00[74]), .in1(tmp00[75]), .out(tmp01[37]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000038(.in0(tmp00[76]), .in1(tmp00[77]), .out(tmp01[38]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000039(.in0(tmp00[78]), .in1(tmp00[79]), .out(tmp01[39]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000040(.in0(tmp00[80]), .in1(tmp00[81]), .out(tmp01[40]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000041(.in0(tmp00[82]), .in1(tmp00[83]), .out(tmp01[41]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000042(.in0(tmp00[84]), .in1(tmp00[85]), .out(tmp01[42]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000043(.in0(tmp00[86]), .in1(tmp00[87]), .out(tmp01[43]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000044(.in0(tmp00[88]), .in1(tmp00[89]), .out(tmp01[44]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000045(.in0(tmp00[90]), .in1(tmp00[91]), .out(tmp01[45]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000046(.in0(tmp00[92]), .in1(tmp00[93]), .out(tmp01[46]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000047(.in0(tmp00[94]), .in1(tmp00[95]), .out(tmp01[47]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000048(.in0(tmp00[96]), .in1(tmp00[97]), .out(tmp01[48]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000049(.in0(tmp00[98]), .in1(tmp00[99]), .out(tmp01[49]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000050(.in0(tmp00[100]), .in1(tmp00[101]), .out(tmp01[50]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000051(.in0(tmp00[102]), .in1(tmp00[103]), .out(tmp01[51]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000052(.in0(tmp00[104]), .in1(tmp00[105]), .out(tmp01[52]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000053(.in0(tmp00[106]), .in1(tmp00[107]), .out(tmp01[53]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000054(.in0(tmp00[108]), .in1(tmp00[109]), .out(tmp01[54]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000055(.in0(tmp00[110]), .in1(tmp00[111]), .out(tmp01[55]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000056(.in0(tmp00[112]), .in1(tmp00[113]), .out(tmp01[56]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000057(.in0(tmp00[114]), .in1(tmp00[115]), .out(tmp01[57]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000058(.in0(tmp00[116]), .in1(tmp00[117]), .out(tmp01[58]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000059(.in0(tmp00[118]), .in1(tmp00[119]), .out(tmp01[59]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000060(.in0(tmp00[120]), .in1(tmp00[121]), .out(tmp01[60]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000061(.in0(tmp00[122]), .in1(tmp00[123]), .out(tmp01[61]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000062(.in0(tmp00[124]), .in1(tmp00[125]), .out(tmp01[62]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000063(.in0(tmp00[126]), .in1(tmp00[127]), .out(tmp01[63]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000064(.in0(tmp00[128]), .in1(tmp00[129]), .out(tmp01[64]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000065(.in0(tmp00[130]), .in1(tmp00[131]), .out(tmp01[65]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000066(.in0(tmp00[132]), .in1(tmp00[133]), .out(tmp01[66]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000067(.in0(tmp00[134]), .in1(tmp00[135]), .out(tmp01[67]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000068(.in0(tmp00[136]), .in1(tmp00[137]), .out(tmp01[68]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000069(.in0(tmp00[138]), .in1(tmp00[139]), .out(tmp01[69]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000070(.in0(tmp00[140]), .in1(tmp00[141]), .out(tmp01[70]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000071(.in0(tmp00[142]), .in1(tmp00[143]), .out(tmp01[71]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000072(.in0(tmp00[144]), .in1(tmp00[145]), .out(tmp01[72]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000073(.in0(tmp00[146]), .in1(tmp00[147]), .out(tmp01[73]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000074(.in0(tmp00[148]), .in1(tmp00[149]), .out(tmp01[74]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000075(.in0(tmp00[150]), .in1(tmp00[151]), .out(tmp01[75]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000076(.in0(tmp00[152]), .in1(tmp00[153]), .out(tmp01[76]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000077(.in0(tmp00[154]), .in1(tmp00[155]), .out(tmp01[77]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000078(.in0(tmp00[156]), .in1(tmp00[157]), .out(tmp01[78]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000079(.in0(tmp00[158]), .in1(tmp00[159]), .out(tmp01[79]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000080(.in0(tmp00[160]), .in1(tmp00[161]), .out(tmp01[80]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000081(.in0(tmp00[162]), .in1(tmp00[163]), .out(tmp01[81]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000082(.in0(tmp00[164]), .in1(tmp00[165]), .out(tmp01[82]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000083(.in0(tmp00[166]), .in1(tmp00[167]), .out(tmp01[83]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000084(.in0(tmp00[168]), .in1(tmp00[169]), .out(tmp01[84]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000085(.in0(tmp00[170]), .in1(tmp00[171]), .out(tmp01[85]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000086(.in0(tmp00[172]), .in1(tmp00[173]), .out(tmp01[86]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000087(.in0(tmp00[174]), .in1(tmp00[175]), .out(tmp01[87]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000088(.in0(tmp00[176]), .in1(tmp00[177]), .out(tmp01[88]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000089(.in0(tmp00[178]), .in1(tmp00[179]), .out(tmp01[89]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000090(.in0(tmp00[180]), .in1(tmp00[181]), .out(tmp01[90]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000091(.in0(tmp00[182]), .in1(tmp00[183]), .out(tmp01[91]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000092(.in0(tmp00[184]), .in1(tmp00[185]), .out(tmp01[92]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000093(.in0(tmp00[186]), .in1(tmp00[187]), .out(tmp01[93]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000094(.in0(tmp00[188]), .in1(tmp00[189]), .out(tmp01[94]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000095(.in0(tmp00[190]), .in1(tmp00[191]), .out(tmp01[95]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000096(.in0(tmp00[192]), .in1(tmp00[193]), .out(tmp01[96]));
	assign tmp01[97] = $signed(tmp00[194]);
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000097(.in0(tmp01[0]), .in1(tmp01[1]), .out(tmp02[0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000098(.in0(tmp01[2]), .in1(tmp01[3]), .out(tmp02[1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000099(.in0(tmp01[4]), .in1(tmp01[5]), .out(tmp02[2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000100(.in0(tmp01[6]), .in1(tmp01[7]), .out(tmp02[3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000101(.in0(tmp01[8]), .in1(tmp01[9]), .out(tmp02[4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000102(.in0(tmp01[10]), .in1(tmp01[11]), .out(tmp02[5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000103(.in0(tmp01[12]), .in1(tmp01[13]), .out(tmp02[6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000104(.in0(tmp01[14]), .in1(tmp01[15]), .out(tmp02[7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000105(.in0(tmp01[16]), .in1(tmp01[17]), .out(tmp02[8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000106(.in0(tmp01[18]), .in1(tmp01[19]), .out(tmp02[9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000107(.in0(tmp01[20]), .in1(tmp01[21]), .out(tmp02[10]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000108(.in0(tmp01[22]), .in1(tmp01[23]), .out(tmp02[11]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000109(.in0(tmp01[24]), .in1(tmp01[25]), .out(tmp02[12]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000110(.in0(tmp01[26]), .in1(tmp01[27]), .out(tmp02[13]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000111(.in0(tmp01[28]), .in1(tmp01[29]), .out(tmp02[14]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000112(.in0(tmp01[30]), .in1(tmp01[31]), .out(tmp02[15]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000113(.in0(tmp01[32]), .in1(tmp01[33]), .out(tmp02[16]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000114(.in0(tmp01[34]), .in1(tmp01[35]), .out(tmp02[17]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000115(.in0(tmp01[36]), .in1(tmp01[37]), .out(tmp02[18]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000116(.in0(tmp01[38]), .in1(tmp01[39]), .out(tmp02[19]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000117(.in0(tmp01[40]), .in1(tmp01[41]), .out(tmp02[20]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000118(.in0(tmp01[42]), .in1(tmp01[43]), .out(tmp02[21]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000119(.in0(tmp01[44]), .in1(tmp01[45]), .out(tmp02[22]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000120(.in0(tmp01[46]), .in1(tmp01[47]), .out(tmp02[23]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000121(.in0(tmp01[48]), .in1(tmp01[49]), .out(tmp02[24]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000122(.in0(tmp01[50]), .in1(tmp01[51]), .out(tmp02[25]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000123(.in0(tmp01[52]), .in1(tmp01[53]), .out(tmp02[26]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000124(.in0(tmp01[54]), .in1(tmp01[55]), .out(tmp02[27]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000125(.in0(tmp01[56]), .in1(tmp01[57]), .out(tmp02[28]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000126(.in0(tmp01[58]), .in1(tmp01[59]), .out(tmp02[29]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000127(.in0(tmp01[60]), .in1(tmp01[61]), .out(tmp02[30]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000128(.in0(tmp01[62]), .in1(tmp01[63]), .out(tmp02[31]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000129(.in0(tmp01[64]), .in1(tmp01[65]), .out(tmp02[32]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000130(.in0(tmp01[66]), .in1(tmp01[67]), .out(tmp02[33]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000131(.in0(tmp01[68]), .in1(tmp01[69]), .out(tmp02[34]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000132(.in0(tmp01[70]), .in1(tmp01[71]), .out(tmp02[35]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000133(.in0(tmp01[72]), .in1(tmp01[73]), .out(tmp02[36]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000134(.in0(tmp01[74]), .in1(tmp01[75]), .out(tmp02[37]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000135(.in0(tmp01[76]), .in1(tmp01[77]), .out(tmp02[38]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000136(.in0(tmp01[78]), .in1(tmp01[79]), .out(tmp02[39]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000137(.in0(tmp01[80]), .in1(tmp01[81]), .out(tmp02[40]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000138(.in0(tmp01[82]), .in1(tmp01[83]), .out(tmp02[41]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000139(.in0(tmp01[84]), .in1(tmp01[85]), .out(tmp02[42]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000140(.in0(tmp01[86]), .in1(tmp01[87]), .out(tmp02[43]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000141(.in0(tmp01[88]), .in1(tmp01[89]), .out(tmp02[44]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000142(.in0(tmp01[90]), .in1(tmp01[91]), .out(tmp02[45]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000143(.in0(tmp01[92]), .in1(tmp01[93]), .out(tmp02[46]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000144(.in0(tmp01[94]), .in1(tmp01[95]), .out(tmp02[47]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000145(.in0(tmp01[96]), .in1(tmp01[97]), .out(tmp02[48]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000146(.in0(tmp02[0]), .in1(tmp02[1]), .out(tmp03[0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000147(.in0(tmp02[2]), .in1(tmp02[3]), .out(tmp03[1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000148(.in0(tmp02[4]), .in1(tmp02[5]), .out(tmp03[2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000149(.in0(tmp02[6]), .in1(tmp02[7]), .out(tmp03[3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000150(.in0(tmp02[8]), .in1(tmp02[9]), .out(tmp03[4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000151(.in0(tmp02[10]), .in1(tmp02[11]), .out(tmp03[5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000152(.in0(tmp02[12]), .in1(tmp02[13]), .out(tmp03[6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000153(.in0(tmp02[14]), .in1(tmp02[15]), .out(tmp03[7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000154(.in0(tmp02[16]), .in1(tmp02[17]), .out(tmp03[8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000155(.in0(tmp02[18]), .in1(tmp02[19]), .out(tmp03[9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000156(.in0(tmp02[20]), .in1(tmp02[21]), .out(tmp03[10]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000157(.in0(tmp02[22]), .in1(tmp02[23]), .out(tmp03[11]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000158(.in0(tmp02[24]), .in1(tmp02[25]), .out(tmp03[12]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000159(.in0(tmp02[26]), .in1(tmp02[27]), .out(tmp03[13]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000160(.in0(tmp02[28]), .in1(tmp02[29]), .out(tmp03[14]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000161(.in0(tmp02[30]), .in1(tmp02[31]), .out(tmp03[15]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000162(.in0(tmp02[32]), .in1(tmp02[33]), .out(tmp03[16]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000163(.in0(tmp02[34]), .in1(tmp02[35]), .out(tmp03[17]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000164(.in0(tmp02[36]), .in1(tmp02[37]), .out(tmp03[18]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000165(.in0(tmp02[38]), .in1(tmp02[39]), .out(tmp03[19]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000166(.in0(tmp02[40]), .in1(tmp02[41]), .out(tmp03[20]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000167(.in0(tmp02[42]), .in1(tmp02[43]), .out(tmp03[21]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000168(.in0(tmp02[44]), .in1(tmp02[45]), .out(tmp03[22]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000169(.in0(tmp02[46]), .in1(tmp02[47]), .out(tmp03[23]));
	assign tmp03[24] = $signed(tmp02[48]);
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000170(.in0(tmp03[0]), .in1(tmp03[1]), .out(tmp04[0]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000171(.in0(tmp03[2]), .in1(tmp03[3]), .out(tmp04[1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000172(.in0(tmp03[4]), .in1(tmp03[5]), .out(tmp04[2]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000173(.in0(tmp03[6]), .in1(tmp03[7]), .out(tmp04[3]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000174(.in0(tmp03[8]), .in1(tmp03[9]), .out(tmp04[4]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000175(.in0(tmp03[10]), .in1(tmp03[11]), .out(tmp04[5]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000176(.in0(tmp03[12]), .in1(tmp03[13]), .out(tmp04[6]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000177(.in0(tmp03[14]), .in1(tmp03[15]), .out(tmp04[7]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000178(.in0(tmp03[16]), .in1(tmp03[17]), .out(tmp04[8]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000179(.in0(tmp03[18]), .in1(tmp03[19]), .out(tmp04[9]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000180(.in0(tmp03[20]), .in1(tmp03[21]), .out(tmp04[10]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000181(.in0(tmp03[22]), .in1(tmp03[23]), .out(tmp04[11]));
	assign tmp04[12] = $signed(tmp03[24]);
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000182(.in0(tmp04[0]), .in1(tmp04[1]), .out(tmp05[0]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000183(.in0(tmp04[2]), .in1(tmp04[3]), .out(tmp05[1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000184(.in0(tmp04[4]), .in1(tmp04[5]), .out(tmp05[2]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000185(.in0(tmp04[6]), .in1(tmp04[7]), .out(tmp05[3]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000186(.in0(tmp04[8]), .in1(tmp04[9]), .out(tmp05[4]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000187(.in0(tmp04[10]), .in1(tmp04[11]), .out(tmp05[5]));
	assign tmp05[6] = $signed(tmp04[12]);
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000188(.in0(tmp05[0]), .in1(tmp05[1]), .out(tmp06[0]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000189(.in0(tmp05[2]), .in1(tmp05[3]), .out(tmp06[1]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000190(.in0(tmp05[4]), .in1(tmp05[5]), .out(tmp06[2]));
	assign tmp06[3] = $signed(tmp05[6]);
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000191(.in0(tmp06[0]), .in1(tmp06[1]), .out(tmp07[0]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000192(.in0(tmp06[2]), .in1(tmp06[3]), .out(tmp07[1]));
	add2 #(.I_WIDTH(WIDTH*2+7), .O_WIDTH(WIDTH*2+8)) add000193(.in0(tmp07[0]), .in1(tmp07[1]), .out(tmp08[0]));
	relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU(.a(tmp08[0]), .b(24'h0), .sel(tmp08[0][WIDTH*2+$clog2(IN)-1]), .out(z));
endmodule

