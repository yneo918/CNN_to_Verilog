module fc84_10
	#(parameter WIDTH = 8, IN = 84, OUT = 10)
	(x, z);
	input [WIDTH-1:0] x[0:IN-1];
	output [WIDTH*2+$clog2(IN)-1:0] z[0:OUT-1];
	wire [WIDTH*2-1+0:0] tmp00[0:83][0:OUT-1];
	wire [WIDTH*2-1+1:0] tmp01[0:41][0:OUT-1];
	wire [WIDTH*2-1+2:0] tmp02[0:20][0:OUT-1];
	wire [WIDTH*2-1+3:0] tmp03[0:10][0:OUT-1];
	wire [WIDTH*2-1+4:0] tmp04[0:5][0:OUT-1];
	wire [WIDTH*2-1+5:0] tmp05[0:2][0:OUT-1];
	wire [WIDTH*2-1+6:0] tmp06[0:1][0:OUT-1];
	wire [WIDTH*2-1+7:0] tmp07[0:0][0:OUT-1];

	booth__006 #(.WIDTH(WIDTH)) mul00000000(.x(x[0]), .z(tmp00[0][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000001(.x(x[1]), .z(tmp00[1][0]));
	booth_0008 #(.WIDTH(WIDTH)) mul00000002(.x(x[2]), .z(tmp00[2][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000003(.x(x[3]), .z(tmp00[3][0]));
	booth_0008 #(.WIDTH(WIDTH)) mul00000004(.x(x[4]), .z(tmp00[4][0]));
	booth_0004 #(.WIDTH(WIDTH)) mul00000005(.x(x[5]), .z(tmp00[5][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000006(.x(x[6]), .z(tmp00[6][0]));
	booth_0006 #(.WIDTH(WIDTH)) mul00000007(.x(x[7]), .z(tmp00[7][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000008(.x(x[8]), .z(tmp00[8][0]));
	booth__008 #(.WIDTH(WIDTH)) mul00000009(.x(x[9]), .z(tmp00[9][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000010(.x(x[10]), .z(tmp00[10][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000011(.x(x[11]), .z(tmp00[11][0]));
	booth_0008 #(.WIDTH(WIDTH)) mul00000012(.x(x[12]), .z(tmp00[12][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000013(.x(x[13]), .z(tmp00[13][0]));
	booth_0004 #(.WIDTH(WIDTH)) mul00000014(.x(x[14]), .z(tmp00[14][0]));
	booth_0004 #(.WIDTH(WIDTH)) mul00000015(.x(x[15]), .z(tmp00[15][0]));
	booth_0004 #(.WIDTH(WIDTH)) mul00000016(.x(x[16]), .z(tmp00[16][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000017(.x(x[17]), .z(tmp00[17][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000018(.x(x[18]), .z(tmp00[18][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000019(.x(x[19]), .z(tmp00[19][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000020(.x(x[20]), .z(tmp00[20][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000021(.x(x[21]), .z(tmp00[21][0]));
	booth_0004 #(.WIDTH(WIDTH)) mul00000022(.x(x[22]), .z(tmp00[22][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000023(.x(x[23]), .z(tmp00[23][0]));
	booth_0006 #(.WIDTH(WIDTH)) mul00000024(.x(x[24]), .z(tmp00[24][0]));
	booth__008 #(.WIDTH(WIDTH)) mul00000025(.x(x[25]), .z(tmp00[25][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000026(.x(x[26]), .z(tmp00[26][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000027(.x(x[27]), .z(tmp00[27][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000028(.x(x[28]), .z(tmp00[28][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000029(.x(x[29]), .z(tmp00[29][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000030(.x(x[30]), .z(tmp00[30][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000031(.x(x[31]), .z(tmp00[31][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000032(.x(x[32]), .z(tmp00[32][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000033(.x(x[33]), .z(tmp00[33][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000034(.x(x[34]), .z(tmp00[34][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000035(.x(x[35]), .z(tmp00[35][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000036(.x(x[36]), .z(tmp00[36][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000037(.x(x[37]), .z(tmp00[37][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000038(.x(x[38]), .z(tmp00[38][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000039(.x(x[39]), .z(tmp00[39][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000040(.x(x[40]), .z(tmp00[40][0]));
	booth_0004 #(.WIDTH(WIDTH)) mul00000041(.x(x[41]), .z(tmp00[41][0]));
	booth__002 #(.WIDTH(WIDTH)) mul00000042(.x(x[42]), .z(tmp00[42][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000043(.x(x[43]), .z(tmp00[43][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000044(.x(x[44]), .z(tmp00[44][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000045(.x(x[45]), .z(tmp00[45][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000046(.x(x[46]), .z(tmp00[46][0]));
	booth__006 #(.WIDTH(WIDTH)) mul00000047(.x(x[47]), .z(tmp00[47][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000048(.x(x[48]), .z(tmp00[48][0]));
	booth_0006 #(.WIDTH(WIDTH)) mul00000049(.x(x[49]), .z(tmp00[49][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000050(.x(x[50]), .z(tmp00[50][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000051(.x(x[51]), .z(tmp00[51][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000052(.x(x[52]), .z(tmp00[52][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000053(.x(x[53]), .z(tmp00[53][0]));
	booth_0006 #(.WIDTH(WIDTH)) mul00000054(.x(x[54]), .z(tmp00[54][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000055(.x(x[55]), .z(tmp00[55][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000056(.x(x[56]), .z(tmp00[56][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000057(.x(x[57]), .z(tmp00[57][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000058(.x(x[58]), .z(tmp00[58][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000059(.x(x[59]), .z(tmp00[59][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000060(.x(x[60]), .z(tmp00[60][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000061(.x(x[61]), .z(tmp00[61][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000062(.x(x[62]), .z(tmp00[62][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000063(.x(x[63]), .z(tmp00[63][0]));
	booth__006 #(.WIDTH(WIDTH)) mul00000064(.x(x[64]), .z(tmp00[64][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000065(.x(x[65]), .z(tmp00[65][0]));
	booth_0006 #(.WIDTH(WIDTH)) mul00000066(.x(x[66]), .z(tmp00[66][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000067(.x(x[67]), .z(tmp00[67][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000068(.x(x[68]), .z(tmp00[68][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000069(.x(x[69]), .z(tmp00[69][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000070(.x(x[70]), .z(tmp00[70][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000071(.x(x[71]), .z(tmp00[71][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000072(.x(x[72]), .z(tmp00[72][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000073(.x(x[73]), .z(tmp00[73][0]));
	booth__002 #(.WIDTH(WIDTH)) mul00000074(.x(x[74]), .z(tmp00[74][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000075(.x(x[75]), .z(tmp00[75][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000076(.x(x[76]), .z(tmp00[76][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000077(.x(x[77]), .z(tmp00[77][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000078(.x(x[78]), .z(tmp00[78][0]));
	booth_0004 #(.WIDTH(WIDTH)) mul00000079(.x(x[79]), .z(tmp00[79][0]));
	booth__004 #(.WIDTH(WIDTH)) mul00000080(.x(x[80]), .z(tmp00[80][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00000081(.x(x[81]), .z(tmp00[81][0]));
	booth__006 #(.WIDTH(WIDTH)) mul00000082(.x(x[82]), .z(tmp00[82][0]));
	booth_0008 #(.WIDTH(WIDTH)) mul00000083(.x(x[83]), .z(tmp00[83][0]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010000(.x(x[0]), .z(tmp00[0][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010001(.x(x[1]), .z(tmp00[1][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010002(.x(x[2]), .z(tmp00[2][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010003(.x(x[3]), .z(tmp00[3][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010004(.x(x[4]), .z(tmp00[4][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010005(.x(x[5]), .z(tmp00[5][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010006(.x(x[6]), .z(tmp00[6][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010007(.x(x[7]), .z(tmp00[7][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010008(.x(x[8]), .z(tmp00[8][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010009(.x(x[9]), .z(tmp00[9][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010010(.x(x[10]), .z(tmp00[10][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010011(.x(x[11]), .z(tmp00[11][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010012(.x(x[12]), .z(tmp00[12][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010013(.x(x[13]), .z(tmp00[13][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010014(.x(x[14]), .z(tmp00[14][1]));
	booth_0006 #(.WIDTH(WIDTH)) mul00010015(.x(x[15]), .z(tmp00[15][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010016(.x(x[16]), .z(tmp00[16][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010017(.x(x[17]), .z(tmp00[17][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010018(.x(x[18]), .z(tmp00[18][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010019(.x(x[19]), .z(tmp00[19][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010020(.x(x[20]), .z(tmp00[20][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010021(.x(x[21]), .z(tmp00[21][1]));
	booth__002 #(.WIDTH(WIDTH)) mul00010022(.x(x[22]), .z(tmp00[22][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010023(.x(x[23]), .z(tmp00[23][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010024(.x(x[24]), .z(tmp00[24][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010025(.x(x[25]), .z(tmp00[25][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010026(.x(x[26]), .z(tmp00[26][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010027(.x(x[27]), .z(tmp00[27][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010028(.x(x[28]), .z(tmp00[28][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010029(.x(x[29]), .z(tmp00[29][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010030(.x(x[30]), .z(tmp00[30][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010031(.x(x[31]), .z(tmp00[31][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010032(.x(x[32]), .z(tmp00[32][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010033(.x(x[33]), .z(tmp00[33][1]));
	booth__008 #(.WIDTH(WIDTH)) mul00010034(.x(x[34]), .z(tmp00[34][1]));
	booth__008 #(.WIDTH(WIDTH)) mul00010035(.x(x[35]), .z(tmp00[35][1]));
	booth_0006 #(.WIDTH(WIDTH)) mul00010036(.x(x[36]), .z(tmp00[36][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010037(.x(x[37]), .z(tmp00[37][1]));
	booth__008 #(.WIDTH(WIDTH)) mul00010038(.x(x[38]), .z(tmp00[38][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010039(.x(x[39]), .z(tmp00[39][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010040(.x(x[40]), .z(tmp00[40][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010041(.x(x[41]), .z(tmp00[41][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010042(.x(x[42]), .z(tmp00[42][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010043(.x(x[43]), .z(tmp00[43][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010044(.x(x[44]), .z(tmp00[44][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010045(.x(x[45]), .z(tmp00[45][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010046(.x(x[46]), .z(tmp00[46][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010047(.x(x[47]), .z(tmp00[47][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010048(.x(x[48]), .z(tmp00[48][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010049(.x(x[49]), .z(tmp00[49][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010050(.x(x[50]), .z(tmp00[50][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010051(.x(x[51]), .z(tmp00[51][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010052(.x(x[52]), .z(tmp00[52][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010053(.x(x[53]), .z(tmp00[53][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010054(.x(x[54]), .z(tmp00[54][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010055(.x(x[55]), .z(tmp00[55][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010056(.x(x[56]), .z(tmp00[56][1]));
	booth_0006 #(.WIDTH(WIDTH)) mul00010057(.x(x[57]), .z(tmp00[57][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010058(.x(x[58]), .z(tmp00[58][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010059(.x(x[59]), .z(tmp00[59][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010060(.x(x[60]), .z(tmp00[60][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010061(.x(x[61]), .z(tmp00[61][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010062(.x(x[62]), .z(tmp00[62][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010063(.x(x[63]), .z(tmp00[63][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010064(.x(x[64]), .z(tmp00[64][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010065(.x(x[65]), .z(tmp00[65][1]));
	booth_0004 #(.WIDTH(WIDTH)) mul00010066(.x(x[66]), .z(tmp00[66][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010067(.x(x[67]), .z(tmp00[67][1]));
	booth_0008 #(.WIDTH(WIDTH)) mul00010068(.x(x[68]), .z(tmp00[68][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010069(.x(x[69]), .z(tmp00[69][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010070(.x(x[70]), .z(tmp00[70][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010071(.x(x[71]), .z(tmp00[71][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010072(.x(x[72]), .z(tmp00[72][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010073(.x(x[73]), .z(tmp00[73][1]));
	booth_0008 #(.WIDTH(WIDTH)) mul00010074(.x(x[74]), .z(tmp00[74][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010075(.x(x[75]), .z(tmp00[75][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010076(.x(x[76]), .z(tmp00[76][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010077(.x(x[77]), .z(tmp00[77][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010078(.x(x[78]), .z(tmp00[78][1]));
	booth_0002 #(.WIDTH(WIDTH)) mul00010079(.x(x[79]), .z(tmp00[79][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010080(.x(x[80]), .z(tmp00[80][1]));
	booth__004 #(.WIDTH(WIDTH)) mul00010081(.x(x[81]), .z(tmp00[81][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010082(.x(x[82]), .z(tmp00[82][1]));
	booth_0000 #(.WIDTH(WIDTH)) mul00010083(.x(x[83]), .z(tmp00[83][1]));
	booth__006 #(.WIDTH(WIDTH)) mul00020000(.x(x[0]), .z(tmp00[0][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020001(.x(x[1]), .z(tmp00[1][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020002(.x(x[2]), .z(tmp00[2][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020003(.x(x[3]), .z(tmp00[3][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020004(.x(x[4]), .z(tmp00[4][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020005(.x(x[5]), .z(tmp00[5][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020006(.x(x[6]), .z(tmp00[6][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020007(.x(x[7]), .z(tmp00[7][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020008(.x(x[8]), .z(tmp00[8][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020009(.x(x[9]), .z(tmp00[9][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020010(.x(x[10]), .z(tmp00[10][2]));
	booth_0002 #(.WIDTH(WIDTH)) mul00020011(.x(x[11]), .z(tmp00[11][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020012(.x(x[12]), .z(tmp00[12][2]));
	booth_0002 #(.WIDTH(WIDTH)) mul00020013(.x(x[13]), .z(tmp00[13][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020014(.x(x[14]), .z(tmp00[14][2]));
	booth__002 #(.WIDTH(WIDTH)) mul00020015(.x(x[15]), .z(tmp00[15][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020016(.x(x[16]), .z(tmp00[16][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020017(.x(x[17]), .z(tmp00[17][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020018(.x(x[18]), .z(tmp00[18][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020019(.x(x[19]), .z(tmp00[19][2]));
	booth__006 #(.WIDTH(WIDTH)) mul00020020(.x(x[20]), .z(tmp00[20][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020021(.x(x[21]), .z(tmp00[21][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020022(.x(x[22]), .z(tmp00[22][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020023(.x(x[23]), .z(tmp00[23][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020024(.x(x[24]), .z(tmp00[24][2]));
	booth__002 #(.WIDTH(WIDTH)) mul00020025(.x(x[25]), .z(tmp00[25][2]));
	booth_0006 #(.WIDTH(WIDTH)) mul00020026(.x(x[26]), .z(tmp00[26][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020027(.x(x[27]), .z(tmp00[27][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020028(.x(x[28]), .z(tmp00[28][2]));
	booth_0006 #(.WIDTH(WIDTH)) mul00020029(.x(x[29]), .z(tmp00[29][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020030(.x(x[30]), .z(tmp00[30][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020031(.x(x[31]), .z(tmp00[31][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020032(.x(x[32]), .z(tmp00[32][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020033(.x(x[33]), .z(tmp00[33][2]));
	booth_0008 #(.WIDTH(WIDTH)) mul00020034(.x(x[34]), .z(tmp00[34][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020035(.x(x[35]), .z(tmp00[35][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020036(.x(x[36]), .z(tmp00[36][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020037(.x(x[37]), .z(tmp00[37][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020038(.x(x[38]), .z(tmp00[38][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020039(.x(x[39]), .z(tmp00[39][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020040(.x(x[40]), .z(tmp00[40][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020041(.x(x[41]), .z(tmp00[41][2]));
	booth_0006 #(.WIDTH(WIDTH)) mul00020042(.x(x[42]), .z(tmp00[42][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020043(.x(x[43]), .z(tmp00[43][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020044(.x(x[44]), .z(tmp00[44][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020045(.x(x[45]), .z(tmp00[45][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020046(.x(x[46]), .z(tmp00[46][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020047(.x(x[47]), .z(tmp00[47][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020048(.x(x[48]), .z(tmp00[48][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020049(.x(x[49]), .z(tmp00[49][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020050(.x(x[50]), .z(tmp00[50][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020051(.x(x[51]), .z(tmp00[51][2]));
	booth__002 #(.WIDTH(WIDTH)) mul00020052(.x(x[52]), .z(tmp00[52][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020053(.x(x[53]), .z(tmp00[53][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020054(.x(x[54]), .z(tmp00[54][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020055(.x(x[55]), .z(tmp00[55][2]));
	booth_0002 #(.WIDTH(WIDTH)) mul00020056(.x(x[56]), .z(tmp00[56][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020057(.x(x[57]), .z(tmp00[57][2]));
	booth_0002 #(.WIDTH(WIDTH)) mul00020058(.x(x[58]), .z(tmp00[58][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020059(.x(x[59]), .z(tmp00[59][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020060(.x(x[60]), .z(tmp00[60][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020061(.x(x[61]), .z(tmp00[61][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020062(.x(x[62]), .z(tmp00[62][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020063(.x(x[63]), .z(tmp00[63][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020064(.x(x[64]), .z(tmp00[64][2]));
	booth_0008 #(.WIDTH(WIDTH)) mul00020065(.x(x[65]), .z(tmp00[65][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020066(.x(x[66]), .z(tmp00[66][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020067(.x(x[67]), .z(tmp00[67][2]));
	booth__006 #(.WIDTH(WIDTH)) mul00020068(.x(x[68]), .z(tmp00[68][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020069(.x(x[69]), .z(tmp00[69][2]));
	booth__006 #(.WIDTH(WIDTH)) mul00020070(.x(x[70]), .z(tmp00[70][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020071(.x(x[71]), .z(tmp00[71][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020072(.x(x[72]), .z(tmp00[72][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020073(.x(x[73]), .z(tmp00[73][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020074(.x(x[74]), .z(tmp00[74][2]));
	booth__006 #(.WIDTH(WIDTH)) mul00020075(.x(x[75]), .z(tmp00[75][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020076(.x(x[76]), .z(tmp00[76][2]));
	booth__006 #(.WIDTH(WIDTH)) mul00020077(.x(x[77]), .z(tmp00[77][2]));
	booth__004 #(.WIDTH(WIDTH)) mul00020078(.x(x[78]), .z(tmp00[78][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020079(.x(x[79]), .z(tmp00[79][2]));
	booth__006 #(.WIDTH(WIDTH)) mul00020080(.x(x[80]), .z(tmp00[80][2]));
	booth_0004 #(.WIDTH(WIDTH)) mul00020081(.x(x[81]), .z(tmp00[81][2]));
	booth_0000 #(.WIDTH(WIDTH)) mul00020082(.x(x[82]), .z(tmp00[82][2]));
	booth__008 #(.WIDTH(WIDTH)) mul00020083(.x(x[83]), .z(tmp00[83][2]));
	booth_0008 #(.WIDTH(WIDTH)) mul00030000(.x(x[0]), .z(tmp00[0][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030001(.x(x[1]), .z(tmp00[1][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030002(.x(x[2]), .z(tmp00[2][3]));
	booth__008 #(.WIDTH(WIDTH)) mul00030003(.x(x[3]), .z(tmp00[3][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030004(.x(x[4]), .z(tmp00[4][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030005(.x(x[5]), .z(tmp00[5][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030006(.x(x[6]), .z(tmp00[6][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030007(.x(x[7]), .z(tmp00[7][3]));
	booth_0006 #(.WIDTH(WIDTH)) mul00030008(.x(x[8]), .z(tmp00[8][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030009(.x(x[9]), .z(tmp00[9][3]));
	booth_0008 #(.WIDTH(WIDTH)) mul00030010(.x(x[10]), .z(tmp00[10][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030011(.x(x[11]), .z(tmp00[11][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030012(.x(x[12]), .z(tmp00[12][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030013(.x(x[13]), .z(tmp00[13][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030014(.x(x[14]), .z(tmp00[14][3]));
	booth__002 #(.WIDTH(WIDTH)) mul00030015(.x(x[15]), .z(tmp00[15][3]));
	booth_0002 #(.WIDTH(WIDTH)) mul00030016(.x(x[16]), .z(tmp00[16][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030017(.x(x[17]), .z(tmp00[17][3]));
	booth_0006 #(.WIDTH(WIDTH)) mul00030018(.x(x[18]), .z(tmp00[18][3]));
	booth_0002 #(.WIDTH(WIDTH)) mul00030019(.x(x[19]), .z(tmp00[19][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030020(.x(x[20]), .z(tmp00[20][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030021(.x(x[21]), .z(tmp00[21][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030022(.x(x[22]), .z(tmp00[22][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030023(.x(x[23]), .z(tmp00[23][3]));
	booth__006 #(.WIDTH(WIDTH)) mul00030024(.x(x[24]), .z(tmp00[24][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030025(.x(x[25]), .z(tmp00[25][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030026(.x(x[26]), .z(tmp00[26][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030027(.x(x[27]), .z(tmp00[27][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030028(.x(x[28]), .z(tmp00[28][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030029(.x(x[29]), .z(tmp00[29][3]));
	booth_0006 #(.WIDTH(WIDTH)) mul00030030(.x(x[30]), .z(tmp00[30][3]));
	booth__006 #(.WIDTH(WIDTH)) mul00030031(.x(x[31]), .z(tmp00[31][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030032(.x(x[32]), .z(tmp00[32][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030033(.x(x[33]), .z(tmp00[33][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030034(.x(x[34]), .z(tmp00[34][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030035(.x(x[35]), .z(tmp00[35][3]));
	booth_0002 #(.WIDTH(WIDTH)) mul00030036(.x(x[36]), .z(tmp00[36][3]));
	booth__006 #(.WIDTH(WIDTH)) mul00030037(.x(x[37]), .z(tmp00[37][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030038(.x(x[38]), .z(tmp00[38][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030039(.x(x[39]), .z(tmp00[39][3]));
	booth_0008 #(.WIDTH(WIDTH)) mul00030040(.x(x[40]), .z(tmp00[40][3]));
	booth__006 #(.WIDTH(WIDTH)) mul00030041(.x(x[41]), .z(tmp00[41][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030042(.x(x[42]), .z(tmp00[42][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030043(.x(x[43]), .z(tmp00[43][3]));
	booth__002 #(.WIDTH(WIDTH)) mul00030044(.x(x[44]), .z(tmp00[44][3]));
	booth_0006 #(.WIDTH(WIDTH)) mul00030045(.x(x[45]), .z(tmp00[45][3]));
	booth_0008 #(.WIDTH(WIDTH)) mul00030046(.x(x[46]), .z(tmp00[46][3]));
	booth__002 #(.WIDTH(WIDTH)) mul00030047(.x(x[47]), .z(tmp00[47][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030048(.x(x[48]), .z(tmp00[48][3]));
	booth_0006 #(.WIDTH(WIDTH)) mul00030049(.x(x[49]), .z(tmp00[49][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030050(.x(x[50]), .z(tmp00[50][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030051(.x(x[51]), .z(tmp00[51][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030052(.x(x[52]), .z(tmp00[52][3]));
	booth_0008 #(.WIDTH(WIDTH)) mul00030053(.x(x[53]), .z(tmp00[53][3]));
	booth__006 #(.WIDTH(WIDTH)) mul00030054(.x(x[54]), .z(tmp00[54][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030055(.x(x[55]), .z(tmp00[55][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030056(.x(x[56]), .z(tmp00[56][3]));
	booth_0008 #(.WIDTH(WIDTH)) mul00030057(.x(x[57]), .z(tmp00[57][3]));
	booth__002 #(.WIDTH(WIDTH)) mul00030058(.x(x[58]), .z(tmp00[58][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030059(.x(x[59]), .z(tmp00[59][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030060(.x(x[60]), .z(tmp00[60][3]));
	booth_0006 #(.WIDTH(WIDTH)) mul00030061(.x(x[61]), .z(tmp00[61][3]));
	booth__006 #(.WIDTH(WIDTH)) mul00030062(.x(x[62]), .z(tmp00[62][3]));
	booth__006 #(.WIDTH(WIDTH)) mul00030063(.x(x[63]), .z(tmp00[63][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030064(.x(x[64]), .z(tmp00[64][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030065(.x(x[65]), .z(tmp00[65][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030066(.x(x[66]), .z(tmp00[66][3]));
	booth__002 #(.WIDTH(WIDTH)) mul00030067(.x(x[67]), .z(tmp00[67][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030068(.x(x[68]), .z(tmp00[68][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030069(.x(x[69]), .z(tmp00[69][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030070(.x(x[70]), .z(tmp00[70][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030071(.x(x[71]), .z(tmp00[71][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030072(.x(x[72]), .z(tmp00[72][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030073(.x(x[73]), .z(tmp00[73][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030074(.x(x[74]), .z(tmp00[74][3]));
	booth__004 #(.WIDTH(WIDTH)) mul00030075(.x(x[75]), .z(tmp00[75][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030076(.x(x[76]), .z(tmp00[76][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030077(.x(x[77]), .z(tmp00[77][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030078(.x(x[78]), .z(tmp00[78][3]));
	booth__006 #(.WIDTH(WIDTH)) mul00030079(.x(x[79]), .z(tmp00[79][3]));
	booth__008 #(.WIDTH(WIDTH)) mul00030080(.x(x[80]), .z(tmp00[80][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030081(.x(x[81]), .z(tmp00[81][3]));
	booth_0000 #(.WIDTH(WIDTH)) mul00030082(.x(x[82]), .z(tmp00[82][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00030083(.x(x[83]), .z(tmp00[83][3]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040000(.x(x[0]), .z(tmp00[0][4]));
	booth_0002 #(.WIDTH(WIDTH)) mul00040001(.x(x[1]), .z(tmp00[1][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040002(.x(x[2]), .z(tmp00[2][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040003(.x(x[3]), .z(tmp00[3][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040004(.x(x[4]), .z(tmp00[4][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040005(.x(x[5]), .z(tmp00[5][4]));
	booth__004 #(.WIDTH(WIDTH)) mul00040006(.x(x[6]), .z(tmp00[6][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040007(.x(x[7]), .z(tmp00[7][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040008(.x(x[8]), .z(tmp00[8][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040009(.x(x[9]), .z(tmp00[9][4]));
	booth__004 #(.WIDTH(WIDTH)) mul00040010(.x(x[10]), .z(tmp00[10][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040011(.x(x[11]), .z(tmp00[11][4]));
	booth_0008 #(.WIDTH(WIDTH)) mul00040012(.x(x[12]), .z(tmp00[12][4]));
	booth_0008 #(.WIDTH(WIDTH)) mul00040013(.x(x[13]), .z(tmp00[13][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040014(.x(x[14]), .z(tmp00[14][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040015(.x(x[15]), .z(tmp00[15][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040016(.x(x[16]), .z(tmp00[16][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040017(.x(x[17]), .z(tmp00[17][4]));
	booth_0002 #(.WIDTH(WIDTH)) mul00040018(.x(x[18]), .z(tmp00[18][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040019(.x(x[19]), .z(tmp00[19][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040020(.x(x[20]), .z(tmp00[20][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040021(.x(x[21]), .z(tmp00[21][4]));
	booth__004 #(.WIDTH(WIDTH)) mul00040022(.x(x[22]), .z(tmp00[22][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040023(.x(x[23]), .z(tmp00[23][4]));
	booth_0008 #(.WIDTH(WIDTH)) mul00040024(.x(x[24]), .z(tmp00[24][4]));
	booth_0006 #(.WIDTH(WIDTH)) mul00040025(.x(x[25]), .z(tmp00[25][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040026(.x(x[26]), .z(tmp00[26][4]));
	booth__004 #(.WIDTH(WIDTH)) mul00040027(.x(x[27]), .z(tmp00[27][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040028(.x(x[28]), .z(tmp00[28][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040029(.x(x[29]), .z(tmp00[29][4]));
	booth__008 #(.WIDTH(WIDTH)) mul00040030(.x(x[30]), .z(tmp00[30][4]));
	booth__004 #(.WIDTH(WIDTH)) mul00040031(.x(x[31]), .z(tmp00[31][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040032(.x(x[32]), .z(tmp00[32][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040033(.x(x[33]), .z(tmp00[33][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040034(.x(x[34]), .z(tmp00[34][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040035(.x(x[35]), .z(tmp00[35][4]));
	booth_0006 #(.WIDTH(WIDTH)) mul00040036(.x(x[36]), .z(tmp00[36][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040037(.x(x[37]), .z(tmp00[37][4]));
	booth_0006 #(.WIDTH(WIDTH)) mul00040038(.x(x[38]), .z(tmp00[38][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040039(.x(x[39]), .z(tmp00[39][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040040(.x(x[40]), .z(tmp00[40][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040041(.x(x[41]), .z(tmp00[41][4]));
	booth_0008 #(.WIDTH(WIDTH)) mul00040042(.x(x[42]), .z(tmp00[42][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040043(.x(x[43]), .z(tmp00[43][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040044(.x(x[44]), .z(tmp00[44][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040045(.x(x[45]), .z(tmp00[45][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040046(.x(x[46]), .z(tmp00[46][4]));
	booth__016 #(.WIDTH(WIDTH)) mul00040047(.x(x[47]), .z(tmp00[47][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040048(.x(x[48]), .z(tmp00[48][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040049(.x(x[49]), .z(tmp00[49][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040050(.x(x[50]), .z(tmp00[50][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040051(.x(x[51]), .z(tmp00[51][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040052(.x(x[52]), .z(tmp00[52][4]));
	booth_0008 #(.WIDTH(WIDTH)) mul00040053(.x(x[53]), .z(tmp00[53][4]));
	booth__004 #(.WIDTH(WIDTH)) mul00040054(.x(x[54]), .z(tmp00[54][4]));
	booth__004 #(.WIDTH(WIDTH)) mul00040055(.x(x[55]), .z(tmp00[55][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040056(.x(x[56]), .z(tmp00[56][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040057(.x(x[57]), .z(tmp00[57][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040058(.x(x[58]), .z(tmp00[58][4]));
	booth__004 #(.WIDTH(WIDTH)) mul00040059(.x(x[59]), .z(tmp00[59][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040060(.x(x[60]), .z(tmp00[60][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040061(.x(x[61]), .z(tmp00[61][4]));
	booth_0002 #(.WIDTH(WIDTH)) mul00040062(.x(x[62]), .z(tmp00[62][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040063(.x(x[63]), .z(tmp00[63][4]));
	booth_0002 #(.WIDTH(WIDTH)) mul00040064(.x(x[64]), .z(tmp00[64][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040065(.x(x[65]), .z(tmp00[65][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040066(.x(x[66]), .z(tmp00[66][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040067(.x(x[67]), .z(tmp00[67][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040068(.x(x[68]), .z(tmp00[68][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040069(.x(x[69]), .z(tmp00[69][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040070(.x(x[70]), .z(tmp00[70][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040071(.x(x[71]), .z(tmp00[71][4]));
	booth__008 #(.WIDTH(WIDTH)) mul00040072(.x(x[72]), .z(tmp00[72][4]));
	booth__008 #(.WIDTH(WIDTH)) mul00040073(.x(x[73]), .z(tmp00[73][4]));
	booth_0008 #(.WIDTH(WIDTH)) mul00040074(.x(x[74]), .z(tmp00[74][4]));
	booth__002 #(.WIDTH(WIDTH)) mul00040075(.x(x[75]), .z(tmp00[75][4]));
	booth__008 #(.WIDTH(WIDTH)) mul00040076(.x(x[76]), .z(tmp00[76][4]));
	booth_0012 #(.WIDTH(WIDTH)) mul00040077(.x(x[77]), .z(tmp00[77][4]));
	booth_0002 #(.WIDTH(WIDTH)) mul00040078(.x(x[78]), .z(tmp00[78][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040079(.x(x[79]), .z(tmp00[79][4]));
	booth_0004 #(.WIDTH(WIDTH)) mul00040080(.x(x[80]), .z(tmp00[80][4]));
	booth_0008 #(.WIDTH(WIDTH)) mul00040081(.x(x[81]), .z(tmp00[81][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040082(.x(x[82]), .z(tmp00[82][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00040083(.x(x[83]), .z(tmp00[83][4]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050000(.x(x[0]), .z(tmp00[0][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050001(.x(x[1]), .z(tmp00[1][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050002(.x(x[2]), .z(tmp00[2][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050003(.x(x[3]), .z(tmp00[3][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050004(.x(x[4]), .z(tmp00[4][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050005(.x(x[5]), .z(tmp00[5][5]));
	booth__002 #(.WIDTH(WIDTH)) mul00050006(.x(x[6]), .z(tmp00[6][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050007(.x(x[7]), .z(tmp00[7][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050008(.x(x[8]), .z(tmp00[8][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050009(.x(x[9]), .z(tmp00[9][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050010(.x(x[10]), .z(tmp00[10][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050011(.x(x[11]), .z(tmp00[11][5]));
	booth_0006 #(.WIDTH(WIDTH)) mul00050012(.x(x[12]), .z(tmp00[12][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050013(.x(x[13]), .z(tmp00[13][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050014(.x(x[14]), .z(tmp00[14][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050015(.x(x[15]), .z(tmp00[15][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050016(.x(x[16]), .z(tmp00[16][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050017(.x(x[17]), .z(tmp00[17][5]));
	booth__002 #(.WIDTH(WIDTH)) mul00050018(.x(x[18]), .z(tmp00[18][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050019(.x(x[19]), .z(tmp00[19][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050020(.x(x[20]), .z(tmp00[20][5]));
	booth_0002 #(.WIDTH(WIDTH)) mul00050021(.x(x[21]), .z(tmp00[21][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050022(.x(x[22]), .z(tmp00[22][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050023(.x(x[23]), .z(tmp00[23][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050024(.x(x[24]), .z(tmp00[24][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050025(.x(x[25]), .z(tmp00[25][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050026(.x(x[26]), .z(tmp00[26][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050027(.x(x[27]), .z(tmp00[27][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050028(.x(x[28]), .z(tmp00[28][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050029(.x(x[29]), .z(tmp00[29][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050030(.x(x[30]), .z(tmp00[30][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050031(.x(x[31]), .z(tmp00[31][5]));
	booth_0002 #(.WIDTH(WIDTH)) mul00050032(.x(x[32]), .z(tmp00[32][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050033(.x(x[33]), .z(tmp00[33][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050034(.x(x[34]), .z(tmp00[34][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050035(.x(x[35]), .z(tmp00[35][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050036(.x(x[36]), .z(tmp00[36][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050037(.x(x[37]), .z(tmp00[37][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050038(.x(x[38]), .z(tmp00[38][5]));
	booth_0008 #(.WIDTH(WIDTH)) mul00050039(.x(x[39]), .z(tmp00[39][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050040(.x(x[40]), .z(tmp00[40][5]));
	booth_0002 #(.WIDTH(WIDTH)) mul00050041(.x(x[41]), .z(tmp00[41][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050042(.x(x[42]), .z(tmp00[42][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050043(.x(x[43]), .z(tmp00[43][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050044(.x(x[44]), .z(tmp00[44][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050045(.x(x[45]), .z(tmp00[45][5]));
	booth_0002 #(.WIDTH(WIDTH)) mul00050046(.x(x[46]), .z(tmp00[46][5]));
	booth__006 #(.WIDTH(WIDTH)) mul00050047(.x(x[47]), .z(tmp00[47][5]));
	booth_0002 #(.WIDTH(WIDTH)) mul00050048(.x(x[48]), .z(tmp00[48][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050049(.x(x[49]), .z(tmp00[49][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050050(.x(x[50]), .z(tmp00[50][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050051(.x(x[51]), .z(tmp00[51][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050052(.x(x[52]), .z(tmp00[52][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050053(.x(x[53]), .z(tmp00[53][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050054(.x(x[54]), .z(tmp00[54][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050055(.x(x[55]), .z(tmp00[55][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050056(.x(x[56]), .z(tmp00[56][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050057(.x(x[57]), .z(tmp00[57][5]));
	booth_0006 #(.WIDTH(WIDTH)) mul00050058(.x(x[58]), .z(tmp00[58][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050059(.x(x[59]), .z(tmp00[59][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050060(.x(x[60]), .z(tmp00[60][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050061(.x(x[61]), .z(tmp00[61][5]));
	booth__006 #(.WIDTH(WIDTH)) mul00050062(.x(x[62]), .z(tmp00[62][5]));
	booth_0002 #(.WIDTH(WIDTH)) mul00050063(.x(x[63]), .z(tmp00[63][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050064(.x(x[64]), .z(tmp00[64][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050065(.x(x[65]), .z(tmp00[65][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050066(.x(x[66]), .z(tmp00[66][5]));
	booth__006 #(.WIDTH(WIDTH)) mul00050067(.x(x[67]), .z(tmp00[67][5]));
	booth_0008 #(.WIDTH(WIDTH)) mul00050068(.x(x[68]), .z(tmp00[68][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050069(.x(x[69]), .z(tmp00[69][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050070(.x(x[70]), .z(tmp00[70][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050071(.x(x[71]), .z(tmp00[71][5]));
	booth__004 #(.WIDTH(WIDTH)) mul00050072(.x(x[72]), .z(tmp00[72][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050073(.x(x[73]), .z(tmp00[73][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050074(.x(x[74]), .z(tmp00[74][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050075(.x(x[75]), .z(tmp00[75][5]));
	booth_0004 #(.WIDTH(WIDTH)) mul00050076(.x(x[76]), .z(tmp00[76][5]));
	booth__002 #(.WIDTH(WIDTH)) mul00050077(.x(x[77]), .z(tmp00[77][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050078(.x(x[78]), .z(tmp00[78][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050079(.x(x[79]), .z(tmp00[79][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050080(.x(x[80]), .z(tmp00[80][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050081(.x(x[81]), .z(tmp00[81][5]));
	booth__006 #(.WIDTH(WIDTH)) mul00050082(.x(x[82]), .z(tmp00[82][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00050083(.x(x[83]), .z(tmp00[83][5]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060000(.x(x[0]), .z(tmp00[0][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060001(.x(x[1]), .z(tmp00[1][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060002(.x(x[2]), .z(tmp00[2][6]));
	booth_0002 #(.WIDTH(WIDTH)) mul00060003(.x(x[3]), .z(tmp00[3][6]));
	booth_0002 #(.WIDTH(WIDTH)) mul00060004(.x(x[4]), .z(tmp00[4][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060005(.x(x[5]), .z(tmp00[5][6]));
	booth__006 #(.WIDTH(WIDTH)) mul00060006(.x(x[6]), .z(tmp00[6][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060007(.x(x[7]), .z(tmp00[7][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060008(.x(x[8]), .z(tmp00[8][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060009(.x(x[9]), .z(tmp00[9][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060010(.x(x[10]), .z(tmp00[10][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060011(.x(x[11]), .z(tmp00[11][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060012(.x(x[12]), .z(tmp00[12][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060013(.x(x[13]), .z(tmp00[13][6]));
	booth__006 #(.WIDTH(WIDTH)) mul00060014(.x(x[14]), .z(tmp00[14][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060015(.x(x[15]), .z(tmp00[15][6]));
	booth_0002 #(.WIDTH(WIDTH)) mul00060016(.x(x[16]), .z(tmp00[16][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060017(.x(x[17]), .z(tmp00[17][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060018(.x(x[18]), .z(tmp00[18][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060019(.x(x[19]), .z(tmp00[19][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060020(.x(x[20]), .z(tmp00[20][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060021(.x(x[21]), .z(tmp00[21][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060022(.x(x[22]), .z(tmp00[22][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060023(.x(x[23]), .z(tmp00[23][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060024(.x(x[24]), .z(tmp00[24][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060025(.x(x[25]), .z(tmp00[25][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060026(.x(x[26]), .z(tmp00[26][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060027(.x(x[27]), .z(tmp00[27][6]));
	booth_0008 #(.WIDTH(WIDTH)) mul00060028(.x(x[28]), .z(tmp00[28][6]));
	booth__002 #(.WIDTH(WIDTH)) mul00060029(.x(x[29]), .z(tmp00[29][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060030(.x(x[30]), .z(tmp00[30][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060031(.x(x[31]), .z(tmp00[31][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060032(.x(x[32]), .z(tmp00[32][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060033(.x(x[33]), .z(tmp00[33][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060034(.x(x[34]), .z(tmp00[34][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060035(.x(x[35]), .z(tmp00[35][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060036(.x(x[36]), .z(tmp00[36][6]));
	booth_0002 #(.WIDTH(WIDTH)) mul00060037(.x(x[37]), .z(tmp00[37][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060038(.x(x[38]), .z(tmp00[38][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060039(.x(x[39]), .z(tmp00[39][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060040(.x(x[40]), .z(tmp00[40][6]));
	booth__002 #(.WIDTH(WIDTH)) mul00060041(.x(x[41]), .z(tmp00[41][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060042(.x(x[42]), .z(tmp00[42][6]));
	booth_0006 #(.WIDTH(WIDTH)) mul00060043(.x(x[43]), .z(tmp00[43][6]));
	booth_0002 #(.WIDTH(WIDTH)) mul00060044(.x(x[44]), .z(tmp00[44][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060045(.x(x[45]), .z(tmp00[45][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060046(.x(x[46]), .z(tmp00[46][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060047(.x(x[47]), .z(tmp00[47][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060048(.x(x[48]), .z(tmp00[48][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060049(.x(x[49]), .z(tmp00[49][6]));
	booth_0002 #(.WIDTH(WIDTH)) mul00060050(.x(x[50]), .z(tmp00[50][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060051(.x(x[51]), .z(tmp00[51][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060052(.x(x[52]), .z(tmp00[52][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060053(.x(x[53]), .z(tmp00[53][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060054(.x(x[54]), .z(tmp00[54][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060055(.x(x[55]), .z(tmp00[55][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060056(.x(x[56]), .z(tmp00[56][6]));
	booth_0002 #(.WIDTH(WIDTH)) mul00060057(.x(x[57]), .z(tmp00[57][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060058(.x(x[58]), .z(tmp00[58][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060059(.x(x[59]), .z(tmp00[59][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060060(.x(x[60]), .z(tmp00[60][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060061(.x(x[61]), .z(tmp00[61][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060062(.x(x[62]), .z(tmp00[62][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060063(.x(x[63]), .z(tmp00[63][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060064(.x(x[64]), .z(tmp00[64][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060065(.x(x[65]), .z(tmp00[65][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060066(.x(x[66]), .z(tmp00[66][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060067(.x(x[67]), .z(tmp00[67][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060068(.x(x[68]), .z(tmp00[68][6]));
	booth_0002 #(.WIDTH(WIDTH)) mul00060069(.x(x[69]), .z(tmp00[69][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060070(.x(x[70]), .z(tmp00[70][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060071(.x(x[71]), .z(tmp00[71][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060072(.x(x[72]), .z(tmp00[72][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060073(.x(x[73]), .z(tmp00[73][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060074(.x(x[74]), .z(tmp00[74][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060075(.x(x[75]), .z(tmp00[75][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060076(.x(x[76]), .z(tmp00[76][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060077(.x(x[77]), .z(tmp00[77][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060078(.x(x[78]), .z(tmp00[78][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060079(.x(x[79]), .z(tmp00[79][6]));
	booth__004 #(.WIDTH(WIDTH)) mul00060080(.x(x[80]), .z(tmp00[80][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060081(.x(x[81]), .z(tmp00[81][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00060082(.x(x[82]), .z(tmp00[82][6]));
	booth_0004 #(.WIDTH(WIDTH)) mul00060083(.x(x[83]), .z(tmp00[83][6]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070000(.x(x[0]), .z(tmp00[0][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070001(.x(x[1]), .z(tmp00[1][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070002(.x(x[2]), .z(tmp00[2][7]));
	booth__002 #(.WIDTH(WIDTH)) mul00070003(.x(x[3]), .z(tmp00[3][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070004(.x(x[4]), .z(tmp00[4][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070005(.x(x[5]), .z(tmp00[5][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070006(.x(x[6]), .z(tmp00[6][7]));
	booth_0006 #(.WIDTH(WIDTH)) mul00070007(.x(x[7]), .z(tmp00[7][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070008(.x(x[8]), .z(tmp00[8][7]));
	booth__006 #(.WIDTH(WIDTH)) mul00070009(.x(x[9]), .z(tmp00[9][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070010(.x(x[10]), .z(tmp00[10][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070011(.x(x[11]), .z(tmp00[11][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070012(.x(x[12]), .z(tmp00[12][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070013(.x(x[13]), .z(tmp00[13][7]));
	booth__002 #(.WIDTH(WIDTH)) mul00070014(.x(x[14]), .z(tmp00[14][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070015(.x(x[15]), .z(tmp00[15][7]));
	booth_0006 #(.WIDTH(WIDTH)) mul00070016(.x(x[16]), .z(tmp00[16][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070017(.x(x[17]), .z(tmp00[17][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070018(.x(x[18]), .z(tmp00[18][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070019(.x(x[19]), .z(tmp00[19][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070020(.x(x[20]), .z(tmp00[20][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070021(.x(x[21]), .z(tmp00[21][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070022(.x(x[22]), .z(tmp00[22][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070023(.x(x[23]), .z(tmp00[23][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070024(.x(x[24]), .z(tmp00[24][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070025(.x(x[25]), .z(tmp00[25][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070026(.x(x[26]), .z(tmp00[26][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070027(.x(x[27]), .z(tmp00[27][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070028(.x(x[28]), .z(tmp00[28][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070029(.x(x[29]), .z(tmp00[29][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070030(.x(x[30]), .z(tmp00[30][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070031(.x(x[31]), .z(tmp00[31][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070032(.x(x[32]), .z(tmp00[32][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070033(.x(x[33]), .z(tmp00[33][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070034(.x(x[34]), .z(tmp00[34][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070035(.x(x[35]), .z(tmp00[35][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070036(.x(x[36]), .z(tmp00[36][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070037(.x(x[37]), .z(tmp00[37][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070038(.x(x[38]), .z(tmp00[38][7]));
	booth_0002 #(.WIDTH(WIDTH)) mul00070039(.x(x[39]), .z(tmp00[39][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070040(.x(x[40]), .z(tmp00[40][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070041(.x(x[41]), .z(tmp00[41][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070042(.x(x[42]), .z(tmp00[42][7]));
	booth_0006 #(.WIDTH(WIDTH)) mul00070043(.x(x[43]), .z(tmp00[43][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070044(.x(x[44]), .z(tmp00[44][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070045(.x(x[45]), .z(tmp00[45][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070046(.x(x[46]), .z(tmp00[46][7]));
	booth_0002 #(.WIDTH(WIDTH)) mul00070047(.x(x[47]), .z(tmp00[47][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070048(.x(x[48]), .z(tmp00[48][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070049(.x(x[49]), .z(tmp00[49][7]));
	booth__006 #(.WIDTH(WIDTH)) mul00070050(.x(x[50]), .z(tmp00[50][7]));
	booth__006 #(.WIDTH(WIDTH)) mul00070051(.x(x[51]), .z(tmp00[51][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070052(.x(x[52]), .z(tmp00[52][7]));
	booth__002 #(.WIDTH(WIDTH)) mul00070053(.x(x[53]), .z(tmp00[53][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070054(.x(x[54]), .z(tmp00[54][7]));
	booth_0006 #(.WIDTH(WIDTH)) mul00070055(.x(x[55]), .z(tmp00[55][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070056(.x(x[56]), .z(tmp00[56][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070057(.x(x[57]), .z(tmp00[57][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070058(.x(x[58]), .z(tmp00[58][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070059(.x(x[59]), .z(tmp00[59][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070060(.x(x[60]), .z(tmp00[60][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070061(.x(x[61]), .z(tmp00[61][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070062(.x(x[62]), .z(tmp00[62][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070063(.x(x[63]), .z(tmp00[63][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070064(.x(x[64]), .z(tmp00[64][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070065(.x(x[65]), .z(tmp00[65][7]));
	booth__002 #(.WIDTH(WIDTH)) mul00070066(.x(x[66]), .z(tmp00[66][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070067(.x(x[67]), .z(tmp00[67][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070068(.x(x[68]), .z(tmp00[68][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070069(.x(x[69]), .z(tmp00[69][7]));
	booth__004 #(.WIDTH(WIDTH)) mul00070070(.x(x[70]), .z(tmp00[70][7]));
	booth__010 #(.WIDTH(WIDTH)) mul00070071(.x(x[71]), .z(tmp00[71][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070072(.x(x[72]), .z(tmp00[72][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070073(.x(x[73]), .z(tmp00[73][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070074(.x(x[74]), .z(tmp00[74][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070075(.x(x[75]), .z(tmp00[75][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070076(.x(x[76]), .z(tmp00[76][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070077(.x(x[77]), .z(tmp00[77][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070078(.x(x[78]), .z(tmp00[78][7]));
	booth_0004 #(.WIDTH(WIDTH)) mul00070079(.x(x[79]), .z(tmp00[79][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070080(.x(x[80]), .z(tmp00[80][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070081(.x(x[81]), .z(tmp00[81][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070082(.x(x[82]), .z(tmp00[82][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00070083(.x(x[83]), .z(tmp00[83][7]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080000(.x(x[0]), .z(tmp00[0][8]));
	booth_0008 #(.WIDTH(WIDTH)) mul00080001(.x(x[1]), .z(tmp00[1][8]));
	booth__006 #(.WIDTH(WIDTH)) mul00080002(.x(x[2]), .z(tmp00[2][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080003(.x(x[3]), .z(tmp00[3][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080004(.x(x[4]), .z(tmp00[4][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080005(.x(x[5]), .z(tmp00[5][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080006(.x(x[6]), .z(tmp00[6][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080007(.x(x[7]), .z(tmp00[7][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080008(.x(x[8]), .z(tmp00[8][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080009(.x(x[9]), .z(tmp00[9][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080010(.x(x[10]), .z(tmp00[10][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080011(.x(x[11]), .z(tmp00[11][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080012(.x(x[12]), .z(tmp00[12][8]));
	booth_0002 #(.WIDTH(WIDTH)) mul00080013(.x(x[13]), .z(tmp00[13][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080014(.x(x[14]), .z(tmp00[14][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080015(.x(x[15]), .z(tmp00[15][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080016(.x(x[16]), .z(tmp00[16][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080017(.x(x[17]), .z(tmp00[17][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080018(.x(x[18]), .z(tmp00[18][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080019(.x(x[19]), .z(tmp00[19][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080020(.x(x[20]), .z(tmp00[20][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080021(.x(x[21]), .z(tmp00[21][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080022(.x(x[22]), .z(tmp00[22][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080023(.x(x[23]), .z(tmp00[23][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080024(.x(x[24]), .z(tmp00[24][8]));
	booth__006 #(.WIDTH(WIDTH)) mul00080025(.x(x[25]), .z(tmp00[25][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080026(.x(x[26]), .z(tmp00[26][8]));
	booth_0006 #(.WIDTH(WIDTH)) mul00080027(.x(x[27]), .z(tmp00[27][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080028(.x(x[28]), .z(tmp00[28][8]));
	booth_0008 #(.WIDTH(WIDTH)) mul00080029(.x(x[29]), .z(tmp00[29][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080030(.x(x[30]), .z(tmp00[30][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080031(.x(x[31]), .z(tmp00[31][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080032(.x(x[32]), .z(tmp00[32][8]));
	booth_0002 #(.WIDTH(WIDTH)) mul00080033(.x(x[33]), .z(tmp00[33][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080034(.x(x[34]), .z(tmp00[34][8]));
	booth_0008 #(.WIDTH(WIDTH)) mul00080035(.x(x[35]), .z(tmp00[35][8]));
	booth_0008 #(.WIDTH(WIDTH)) mul00080036(.x(x[36]), .z(tmp00[36][8]));
	booth_0002 #(.WIDTH(WIDTH)) mul00080037(.x(x[37]), .z(tmp00[37][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080038(.x(x[38]), .z(tmp00[38][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080039(.x(x[39]), .z(tmp00[39][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080040(.x(x[40]), .z(tmp00[40][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080041(.x(x[41]), .z(tmp00[41][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080042(.x(x[42]), .z(tmp00[42][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080043(.x(x[43]), .z(tmp00[43][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080044(.x(x[44]), .z(tmp00[44][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080045(.x(x[45]), .z(tmp00[45][8]));
	booth__002 #(.WIDTH(WIDTH)) mul00080046(.x(x[46]), .z(tmp00[46][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080047(.x(x[47]), .z(tmp00[47][8]));
	booth_0002 #(.WIDTH(WIDTH)) mul00080048(.x(x[48]), .z(tmp00[48][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080049(.x(x[49]), .z(tmp00[49][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080050(.x(x[50]), .z(tmp00[50][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080051(.x(x[51]), .z(tmp00[51][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080052(.x(x[52]), .z(tmp00[52][8]));
	booth_0002 #(.WIDTH(WIDTH)) mul00080053(.x(x[53]), .z(tmp00[53][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080054(.x(x[54]), .z(tmp00[54][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080055(.x(x[55]), .z(tmp00[55][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080056(.x(x[56]), .z(tmp00[56][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080057(.x(x[57]), .z(tmp00[57][8]));
	booth_0008 #(.WIDTH(WIDTH)) mul00080058(.x(x[58]), .z(tmp00[58][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080059(.x(x[59]), .z(tmp00[59][8]));
	booth__006 #(.WIDTH(WIDTH)) mul00080060(.x(x[60]), .z(tmp00[60][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080061(.x(x[61]), .z(tmp00[61][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080062(.x(x[62]), .z(tmp00[62][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080063(.x(x[63]), .z(tmp00[63][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080064(.x(x[64]), .z(tmp00[64][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080065(.x(x[65]), .z(tmp00[65][8]));
	booth_0008 #(.WIDTH(WIDTH)) mul00080066(.x(x[66]), .z(tmp00[66][8]));
	booth_0012 #(.WIDTH(WIDTH)) mul00080067(.x(x[67]), .z(tmp00[67][8]));
	booth__008 #(.WIDTH(WIDTH)) mul00080068(.x(x[68]), .z(tmp00[68][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080069(.x(x[69]), .z(tmp00[69][8]));
	booth_0004 #(.WIDTH(WIDTH)) mul00080070(.x(x[70]), .z(tmp00[70][8]));
	booth_0006 #(.WIDTH(WIDTH)) mul00080071(.x(x[71]), .z(tmp00[71][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080072(.x(x[72]), .z(tmp00[72][8]));
	booth__008 #(.WIDTH(WIDTH)) mul00080073(.x(x[73]), .z(tmp00[73][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080074(.x(x[74]), .z(tmp00[74][8]));
	booth_0002 #(.WIDTH(WIDTH)) mul00080075(.x(x[75]), .z(tmp00[75][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080076(.x(x[76]), .z(tmp00[76][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080077(.x(x[77]), .z(tmp00[77][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080078(.x(x[78]), .z(tmp00[78][8]));
	booth_0000 #(.WIDTH(WIDTH)) mul00080079(.x(x[79]), .z(tmp00[79][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080080(.x(x[80]), .z(tmp00[80][8]));
	booth_0002 #(.WIDTH(WIDTH)) mul00080081(.x(x[81]), .z(tmp00[81][8]));
	booth__008 #(.WIDTH(WIDTH)) mul00080082(.x(x[82]), .z(tmp00[82][8]));
	booth__004 #(.WIDTH(WIDTH)) mul00080083(.x(x[83]), .z(tmp00[83][8]));
	booth__002 #(.WIDTH(WIDTH)) mul00090000(.x(x[0]), .z(tmp00[0][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090001(.x(x[1]), .z(tmp00[1][9]));
	booth_0008 #(.WIDTH(WIDTH)) mul00090002(.x(x[2]), .z(tmp00[2][9]));
	booth__008 #(.WIDTH(WIDTH)) mul00090003(.x(x[3]), .z(tmp00[3][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090004(.x(x[4]), .z(tmp00[4][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090005(.x(x[5]), .z(tmp00[5][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090006(.x(x[6]), .z(tmp00[6][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090007(.x(x[7]), .z(tmp00[7][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090008(.x(x[8]), .z(tmp00[8][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090009(.x(x[9]), .z(tmp00[9][9]));
	booth__008 #(.WIDTH(WIDTH)) mul00090010(.x(x[10]), .z(tmp00[10][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090011(.x(x[11]), .z(tmp00[11][9]));
	booth__008 #(.WIDTH(WIDTH)) mul00090012(.x(x[12]), .z(tmp00[12][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090013(.x(x[13]), .z(tmp00[13][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090014(.x(x[14]), .z(tmp00[14][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090015(.x(x[15]), .z(tmp00[15][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090016(.x(x[16]), .z(tmp00[16][9]));
	booth_0008 #(.WIDTH(WIDTH)) mul00090017(.x(x[17]), .z(tmp00[17][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090018(.x(x[18]), .z(tmp00[18][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090019(.x(x[19]), .z(tmp00[19][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090020(.x(x[20]), .z(tmp00[20][9]));
	booth__006 #(.WIDTH(WIDTH)) mul00090021(.x(x[21]), .z(tmp00[21][9]));
	booth__006 #(.WIDTH(WIDTH)) mul00090022(.x(x[22]), .z(tmp00[22][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090023(.x(x[23]), .z(tmp00[23][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090024(.x(x[24]), .z(tmp00[24][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090025(.x(x[25]), .z(tmp00[25][9]));
	booth__002 #(.WIDTH(WIDTH)) mul00090026(.x(x[26]), .z(tmp00[26][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090027(.x(x[27]), .z(tmp00[27][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090028(.x(x[28]), .z(tmp00[28][9]));
	booth_0002 #(.WIDTH(WIDTH)) mul00090029(.x(x[29]), .z(tmp00[29][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090030(.x(x[30]), .z(tmp00[30][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090031(.x(x[31]), .z(tmp00[31][9]));
	booth_0006 #(.WIDTH(WIDTH)) mul00090032(.x(x[32]), .z(tmp00[32][9]));
	booth__002 #(.WIDTH(WIDTH)) mul00090033(.x(x[33]), .z(tmp00[33][9]));
	booth__002 #(.WIDTH(WIDTH)) mul00090034(.x(x[34]), .z(tmp00[34][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090035(.x(x[35]), .z(tmp00[35][9]));
	booth__006 #(.WIDTH(WIDTH)) mul00090036(.x(x[36]), .z(tmp00[36][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090037(.x(x[37]), .z(tmp00[37][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090038(.x(x[38]), .z(tmp00[38][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090039(.x(x[39]), .z(tmp00[39][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090040(.x(x[40]), .z(tmp00[40][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090041(.x(x[41]), .z(tmp00[41][9]));
	booth_0006 #(.WIDTH(WIDTH)) mul00090042(.x(x[42]), .z(tmp00[42][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090043(.x(x[43]), .z(tmp00[43][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090044(.x(x[44]), .z(tmp00[44][9]));
	booth_0008 #(.WIDTH(WIDTH)) mul00090045(.x(x[45]), .z(tmp00[45][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090046(.x(x[46]), .z(tmp00[46][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090047(.x(x[47]), .z(tmp00[47][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090048(.x(x[48]), .z(tmp00[48][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090049(.x(x[49]), .z(tmp00[49][9]));
	booth_0008 #(.WIDTH(WIDTH)) mul00090050(.x(x[50]), .z(tmp00[50][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090051(.x(x[51]), .z(tmp00[51][9]));
	booth__006 #(.WIDTH(WIDTH)) mul00090052(.x(x[52]), .z(tmp00[52][9]));
	booth__008 #(.WIDTH(WIDTH)) mul00090053(.x(x[53]), .z(tmp00[53][9]));
	booth__006 #(.WIDTH(WIDTH)) mul00090054(.x(x[54]), .z(tmp00[54][9]));
	booth_0002 #(.WIDTH(WIDTH)) mul00090055(.x(x[55]), .z(tmp00[55][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090056(.x(x[56]), .z(tmp00[56][9]));
	booth__008 #(.WIDTH(WIDTH)) mul00090057(.x(x[57]), .z(tmp00[57][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090058(.x(x[58]), .z(tmp00[58][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090059(.x(x[59]), .z(tmp00[59][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090060(.x(x[60]), .z(tmp00[60][9]));
	booth__004 #(.WIDTH(WIDTH)) mul00090061(.x(x[61]), .z(tmp00[61][9]));
	booth__002 #(.WIDTH(WIDTH)) mul00090062(.x(x[62]), .z(tmp00[62][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090063(.x(x[63]), .z(tmp00[63][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090064(.x(x[64]), .z(tmp00[64][9]));
	booth__008 #(.WIDTH(WIDTH)) mul00090065(.x(x[65]), .z(tmp00[65][9]));
	booth_0008 #(.WIDTH(WIDTH)) mul00090066(.x(x[66]), .z(tmp00[66][9]));
	booth__006 #(.WIDTH(WIDTH)) mul00090067(.x(x[67]), .z(tmp00[67][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090068(.x(x[68]), .z(tmp00[68][9]));
	booth_0006 #(.WIDTH(WIDTH)) mul00090069(.x(x[69]), .z(tmp00[69][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090070(.x(x[70]), .z(tmp00[70][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090071(.x(x[71]), .z(tmp00[71][9]));
	booth__006 #(.WIDTH(WIDTH)) mul00090072(.x(x[72]), .z(tmp00[72][9]));
	booth__008 #(.WIDTH(WIDTH)) mul00090073(.x(x[73]), .z(tmp00[73][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090074(.x(x[74]), .z(tmp00[74][9]));
	booth__002 #(.WIDTH(WIDTH)) mul00090075(.x(x[75]), .z(tmp00[75][9]));
	booth__002 #(.WIDTH(WIDTH)) mul00090076(.x(x[76]), .z(tmp00[76][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090077(.x(x[77]), .z(tmp00[77][9]));
	booth_0004 #(.WIDTH(WIDTH)) mul00090078(.x(x[78]), .z(tmp00[78][9]));
	booth__002 #(.WIDTH(WIDTH)) mul00090079(.x(x[79]), .z(tmp00[79][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090080(.x(x[80]), .z(tmp00[80][9]));
	booth_0000 #(.WIDTH(WIDTH)) mul00090081(.x(x[81]), .z(tmp00[81][9]));
	booth_0002 #(.WIDTH(WIDTH)) mul00090082(.x(x[82]), .z(tmp00[82][9]));
	booth__006 #(.WIDTH(WIDTH)) mul00090083(.x(x[83]), .z(tmp00[83][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000000(.in0(tmp00[0][0]), .in1(tmp00[1][0]), .out(tmp01[0][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000001(.in0(tmp00[2][0]), .in1(tmp00[3][0]), .out(tmp01[1][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000002(.in0(tmp00[4][0]), .in1(tmp00[5][0]), .out(tmp01[2][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000003(.in0(tmp00[6][0]), .in1(tmp00[7][0]), .out(tmp01[3][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000004(.in0(tmp00[8][0]), .in1(tmp00[9][0]), .out(tmp01[4][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000005(.in0(tmp00[10][0]), .in1(tmp00[11][0]), .out(tmp01[5][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000006(.in0(tmp00[12][0]), .in1(tmp00[13][0]), .out(tmp01[6][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000007(.in0(tmp00[14][0]), .in1(tmp00[15][0]), .out(tmp01[7][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000008(.in0(tmp00[16][0]), .in1(tmp00[17][0]), .out(tmp01[8][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000009(.in0(tmp00[18][0]), .in1(tmp00[19][0]), .out(tmp01[9][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000010(.in0(tmp00[20][0]), .in1(tmp00[21][0]), .out(tmp01[10][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000011(.in0(tmp00[22][0]), .in1(tmp00[23][0]), .out(tmp01[11][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000012(.in0(tmp00[24][0]), .in1(tmp00[25][0]), .out(tmp01[12][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000013(.in0(tmp00[26][0]), .in1(tmp00[27][0]), .out(tmp01[13][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000014(.in0(tmp00[28][0]), .in1(tmp00[29][0]), .out(tmp01[14][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000015(.in0(tmp00[30][0]), .in1(tmp00[31][0]), .out(tmp01[15][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000016(.in0(tmp00[32][0]), .in1(tmp00[33][0]), .out(tmp01[16][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000017(.in0(tmp00[34][0]), .in1(tmp00[35][0]), .out(tmp01[17][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000018(.in0(tmp00[36][0]), .in1(tmp00[37][0]), .out(tmp01[18][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000019(.in0(tmp00[38][0]), .in1(tmp00[39][0]), .out(tmp01[19][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000020(.in0(tmp00[40][0]), .in1(tmp00[41][0]), .out(tmp01[20][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000021(.in0(tmp00[42][0]), .in1(tmp00[43][0]), .out(tmp01[21][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000022(.in0(tmp00[44][0]), .in1(tmp00[45][0]), .out(tmp01[22][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000023(.in0(tmp00[46][0]), .in1(tmp00[47][0]), .out(tmp01[23][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000024(.in0(tmp00[48][0]), .in1(tmp00[49][0]), .out(tmp01[24][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000025(.in0(tmp00[50][0]), .in1(tmp00[51][0]), .out(tmp01[25][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000026(.in0(tmp00[52][0]), .in1(tmp00[53][0]), .out(tmp01[26][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000027(.in0(tmp00[54][0]), .in1(tmp00[55][0]), .out(tmp01[27][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000028(.in0(tmp00[56][0]), .in1(tmp00[57][0]), .out(tmp01[28][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000029(.in0(tmp00[58][0]), .in1(tmp00[59][0]), .out(tmp01[29][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000030(.in0(tmp00[60][0]), .in1(tmp00[61][0]), .out(tmp01[30][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000031(.in0(tmp00[62][0]), .in1(tmp00[63][0]), .out(tmp01[31][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000032(.in0(tmp00[64][0]), .in1(tmp00[65][0]), .out(tmp01[32][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000033(.in0(tmp00[66][0]), .in1(tmp00[67][0]), .out(tmp01[33][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000034(.in0(tmp00[68][0]), .in1(tmp00[69][0]), .out(tmp01[34][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000035(.in0(tmp00[70][0]), .in1(tmp00[71][0]), .out(tmp01[35][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000036(.in0(tmp00[72][0]), .in1(tmp00[73][0]), .out(tmp01[36][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000037(.in0(tmp00[74][0]), .in1(tmp00[75][0]), .out(tmp01[37][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000038(.in0(tmp00[76][0]), .in1(tmp00[77][0]), .out(tmp01[38][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000039(.in0(tmp00[78][0]), .in1(tmp00[79][0]), .out(tmp01[39][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000040(.in0(tmp00[80][0]), .in1(tmp00[81][0]), .out(tmp01[40][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000041(.in0(tmp00[82][0]), .in1(tmp00[83][0]), .out(tmp01[41][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000042(.in0(tmp01[0][0]), .in1(tmp01[1][0]), .out(tmp02[0][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000043(.in0(tmp01[2][0]), .in1(tmp01[3][0]), .out(tmp02[1][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000044(.in0(tmp01[4][0]), .in1(tmp01[5][0]), .out(tmp02[2][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000045(.in0(tmp01[6][0]), .in1(tmp01[7][0]), .out(tmp02[3][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000046(.in0(tmp01[8][0]), .in1(tmp01[9][0]), .out(tmp02[4][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000047(.in0(tmp01[10][0]), .in1(tmp01[11][0]), .out(tmp02[5][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000048(.in0(tmp01[12][0]), .in1(tmp01[13][0]), .out(tmp02[6][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000049(.in0(tmp01[14][0]), .in1(tmp01[15][0]), .out(tmp02[7][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000050(.in0(tmp01[16][0]), .in1(tmp01[17][0]), .out(tmp02[8][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000051(.in0(tmp01[18][0]), .in1(tmp01[19][0]), .out(tmp02[9][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000052(.in0(tmp01[20][0]), .in1(tmp01[21][0]), .out(tmp02[10][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000053(.in0(tmp01[22][0]), .in1(tmp01[23][0]), .out(tmp02[11][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000054(.in0(tmp01[24][0]), .in1(tmp01[25][0]), .out(tmp02[12][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000055(.in0(tmp01[26][0]), .in1(tmp01[27][0]), .out(tmp02[13][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000056(.in0(tmp01[28][0]), .in1(tmp01[29][0]), .out(tmp02[14][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000057(.in0(tmp01[30][0]), .in1(tmp01[31][0]), .out(tmp02[15][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000058(.in0(tmp01[32][0]), .in1(tmp01[33][0]), .out(tmp02[16][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000059(.in0(tmp01[34][0]), .in1(tmp01[35][0]), .out(tmp02[17][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000060(.in0(tmp01[36][0]), .in1(tmp01[37][0]), .out(tmp02[18][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000061(.in0(tmp01[38][0]), .in1(tmp01[39][0]), .out(tmp02[19][0]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000062(.in0(tmp01[40][0]), .in1(tmp01[41][0]), .out(tmp02[20][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000063(.in0(tmp02[0][0]), .in1(tmp02[1][0]), .out(tmp03[0][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000064(.in0(tmp02[2][0]), .in1(tmp02[3][0]), .out(tmp03[1][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000065(.in0(tmp02[4][0]), .in1(tmp02[5][0]), .out(tmp03[2][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000066(.in0(tmp02[6][0]), .in1(tmp02[7][0]), .out(tmp03[3][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000067(.in0(tmp02[8][0]), .in1(tmp02[9][0]), .out(tmp03[4][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000068(.in0(tmp02[10][0]), .in1(tmp02[11][0]), .out(tmp03[5][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000069(.in0(tmp02[12][0]), .in1(tmp02[13][0]), .out(tmp03[6][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000070(.in0(tmp02[14][0]), .in1(tmp02[15][0]), .out(tmp03[7][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000071(.in0(tmp02[16][0]), .in1(tmp02[17][0]), .out(tmp03[8][0]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000072(.in0(tmp02[18][0]), .in1(tmp02[19][0]), .out(tmp03[9][0]));
	assign tmp03[10][0] = 8'(signed'(tmp02[20][0][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000073(.in0(tmp03[0][0]), .in1(tmp03[1][0]), .out(tmp04[0][0]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000074(.in0(tmp03[2][0]), .in1(tmp03[3][0]), .out(tmp04[1][0]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000075(.in0(tmp03[4][0]), .in1(tmp03[5][0]), .out(tmp04[2][0]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000076(.in0(tmp03[6][0]), .in1(tmp03[7][0]), .out(tmp04[3][0]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000077(.in0(tmp03[8][0]), .in1(tmp03[9][0]), .out(tmp04[4][0]));
	assign tmp04[5][0] = 8'(signed'(tmp03[10][0][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000078(.in0(tmp04[0][0]), .in1(tmp04[1][0]), .out(tmp05[0][0]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000079(.in0(tmp04[2][0]), .in1(tmp04[3][0]), .out(tmp05[1][0]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000080(.in0(tmp04[4][0]), .in1(tmp04[5][0]), .out(tmp05[2][0]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000081(.in0(tmp05[0][0]), .in1(tmp05[1][0]), .out(tmp06[0][0]));
	assign tmp06[1][0] = 8'(signed'(tmp05[2][0][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000082(.in0(tmp06[0][0]), .in1(tmp06[1][0]), .out(tmp07[0][0]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000083(.in0(tmp00[0][1]), .in1(tmp00[1][1]), .out(tmp01[0][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000084(.in0(tmp00[2][1]), .in1(tmp00[3][1]), .out(tmp01[1][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000085(.in0(tmp00[4][1]), .in1(tmp00[5][1]), .out(tmp01[2][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000086(.in0(tmp00[6][1]), .in1(tmp00[7][1]), .out(tmp01[3][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000087(.in0(tmp00[8][1]), .in1(tmp00[9][1]), .out(tmp01[4][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000088(.in0(tmp00[10][1]), .in1(tmp00[11][1]), .out(tmp01[5][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000089(.in0(tmp00[12][1]), .in1(tmp00[13][1]), .out(tmp01[6][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000090(.in0(tmp00[14][1]), .in1(tmp00[15][1]), .out(tmp01[7][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000091(.in0(tmp00[16][1]), .in1(tmp00[17][1]), .out(tmp01[8][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000092(.in0(tmp00[18][1]), .in1(tmp00[19][1]), .out(tmp01[9][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000093(.in0(tmp00[20][1]), .in1(tmp00[21][1]), .out(tmp01[10][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000094(.in0(tmp00[22][1]), .in1(tmp00[23][1]), .out(tmp01[11][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000095(.in0(tmp00[24][1]), .in1(tmp00[25][1]), .out(tmp01[12][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000096(.in0(tmp00[26][1]), .in1(tmp00[27][1]), .out(tmp01[13][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000097(.in0(tmp00[28][1]), .in1(tmp00[29][1]), .out(tmp01[14][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000098(.in0(tmp00[30][1]), .in1(tmp00[31][1]), .out(tmp01[15][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000099(.in0(tmp00[32][1]), .in1(tmp00[33][1]), .out(tmp01[16][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000100(.in0(tmp00[34][1]), .in1(tmp00[35][1]), .out(tmp01[17][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000101(.in0(tmp00[36][1]), .in1(tmp00[37][1]), .out(tmp01[18][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000102(.in0(tmp00[38][1]), .in1(tmp00[39][1]), .out(tmp01[19][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000103(.in0(tmp00[40][1]), .in1(tmp00[41][1]), .out(tmp01[20][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000104(.in0(tmp00[42][1]), .in1(tmp00[43][1]), .out(tmp01[21][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000105(.in0(tmp00[44][1]), .in1(tmp00[45][1]), .out(tmp01[22][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000106(.in0(tmp00[46][1]), .in1(tmp00[47][1]), .out(tmp01[23][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000107(.in0(tmp00[48][1]), .in1(tmp00[49][1]), .out(tmp01[24][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000108(.in0(tmp00[50][1]), .in1(tmp00[51][1]), .out(tmp01[25][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000109(.in0(tmp00[52][1]), .in1(tmp00[53][1]), .out(tmp01[26][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000110(.in0(tmp00[54][1]), .in1(tmp00[55][1]), .out(tmp01[27][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000111(.in0(tmp00[56][1]), .in1(tmp00[57][1]), .out(tmp01[28][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000112(.in0(tmp00[58][1]), .in1(tmp00[59][1]), .out(tmp01[29][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000113(.in0(tmp00[60][1]), .in1(tmp00[61][1]), .out(tmp01[30][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000114(.in0(tmp00[62][1]), .in1(tmp00[63][1]), .out(tmp01[31][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000115(.in0(tmp00[64][1]), .in1(tmp00[65][1]), .out(tmp01[32][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000116(.in0(tmp00[66][1]), .in1(tmp00[67][1]), .out(tmp01[33][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000117(.in0(tmp00[68][1]), .in1(tmp00[69][1]), .out(tmp01[34][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000118(.in0(tmp00[70][1]), .in1(tmp00[71][1]), .out(tmp01[35][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000119(.in0(tmp00[72][1]), .in1(tmp00[73][1]), .out(tmp01[36][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000120(.in0(tmp00[74][1]), .in1(tmp00[75][1]), .out(tmp01[37][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000121(.in0(tmp00[76][1]), .in1(tmp00[77][1]), .out(tmp01[38][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000122(.in0(tmp00[78][1]), .in1(tmp00[79][1]), .out(tmp01[39][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000123(.in0(tmp00[80][1]), .in1(tmp00[81][1]), .out(tmp01[40][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000124(.in0(tmp00[82][1]), .in1(tmp00[83][1]), .out(tmp01[41][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000125(.in0(tmp01[0][1]), .in1(tmp01[1][1]), .out(tmp02[0][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000126(.in0(tmp01[2][1]), .in1(tmp01[3][1]), .out(tmp02[1][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000127(.in0(tmp01[4][1]), .in1(tmp01[5][1]), .out(tmp02[2][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000128(.in0(tmp01[6][1]), .in1(tmp01[7][1]), .out(tmp02[3][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000129(.in0(tmp01[8][1]), .in1(tmp01[9][1]), .out(tmp02[4][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000130(.in0(tmp01[10][1]), .in1(tmp01[11][1]), .out(tmp02[5][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000131(.in0(tmp01[12][1]), .in1(tmp01[13][1]), .out(tmp02[6][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000132(.in0(tmp01[14][1]), .in1(tmp01[15][1]), .out(tmp02[7][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000133(.in0(tmp01[16][1]), .in1(tmp01[17][1]), .out(tmp02[8][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000134(.in0(tmp01[18][1]), .in1(tmp01[19][1]), .out(tmp02[9][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000135(.in0(tmp01[20][1]), .in1(tmp01[21][1]), .out(tmp02[10][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000136(.in0(tmp01[22][1]), .in1(tmp01[23][1]), .out(tmp02[11][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000137(.in0(tmp01[24][1]), .in1(tmp01[25][1]), .out(tmp02[12][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000138(.in0(tmp01[26][1]), .in1(tmp01[27][1]), .out(tmp02[13][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000139(.in0(tmp01[28][1]), .in1(tmp01[29][1]), .out(tmp02[14][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000140(.in0(tmp01[30][1]), .in1(tmp01[31][1]), .out(tmp02[15][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000141(.in0(tmp01[32][1]), .in1(tmp01[33][1]), .out(tmp02[16][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000142(.in0(tmp01[34][1]), .in1(tmp01[35][1]), .out(tmp02[17][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000143(.in0(tmp01[36][1]), .in1(tmp01[37][1]), .out(tmp02[18][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000144(.in0(tmp01[38][1]), .in1(tmp01[39][1]), .out(tmp02[19][1]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000145(.in0(tmp01[40][1]), .in1(tmp01[41][1]), .out(tmp02[20][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000146(.in0(tmp02[0][1]), .in1(tmp02[1][1]), .out(tmp03[0][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000147(.in0(tmp02[2][1]), .in1(tmp02[3][1]), .out(tmp03[1][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000148(.in0(tmp02[4][1]), .in1(tmp02[5][1]), .out(tmp03[2][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000149(.in0(tmp02[6][1]), .in1(tmp02[7][1]), .out(tmp03[3][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000150(.in0(tmp02[8][1]), .in1(tmp02[9][1]), .out(tmp03[4][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000151(.in0(tmp02[10][1]), .in1(tmp02[11][1]), .out(tmp03[5][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000152(.in0(tmp02[12][1]), .in1(tmp02[13][1]), .out(tmp03[6][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000153(.in0(tmp02[14][1]), .in1(tmp02[15][1]), .out(tmp03[7][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000154(.in0(tmp02[16][1]), .in1(tmp02[17][1]), .out(tmp03[8][1]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000155(.in0(tmp02[18][1]), .in1(tmp02[19][1]), .out(tmp03[9][1]));
	assign tmp03[10][1] = 8'(signed'(tmp02[20][1][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000156(.in0(tmp03[0][1]), .in1(tmp03[1][1]), .out(tmp04[0][1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000157(.in0(tmp03[2][1]), .in1(tmp03[3][1]), .out(tmp04[1][1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000158(.in0(tmp03[4][1]), .in1(tmp03[5][1]), .out(tmp04[2][1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000159(.in0(tmp03[6][1]), .in1(tmp03[7][1]), .out(tmp04[3][1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000160(.in0(tmp03[8][1]), .in1(tmp03[9][1]), .out(tmp04[4][1]));
	assign tmp04[5][1] = 8'(signed'(tmp03[10][1][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000161(.in0(tmp04[0][1]), .in1(tmp04[1][1]), .out(tmp05[0][1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000162(.in0(tmp04[2][1]), .in1(tmp04[3][1]), .out(tmp05[1][1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000163(.in0(tmp04[4][1]), .in1(tmp04[5][1]), .out(tmp05[2][1]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000164(.in0(tmp05[0][1]), .in1(tmp05[1][1]), .out(tmp06[0][1]));
	assign tmp06[1][1] = 8'(signed'(tmp05[2][1][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000165(.in0(tmp06[0][1]), .in1(tmp06[1][1]), .out(tmp07[0][1]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000166(.in0(tmp00[0][2]), .in1(tmp00[1][2]), .out(tmp01[0][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000167(.in0(tmp00[2][2]), .in1(tmp00[3][2]), .out(tmp01[1][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000168(.in0(tmp00[4][2]), .in1(tmp00[5][2]), .out(tmp01[2][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000169(.in0(tmp00[6][2]), .in1(tmp00[7][2]), .out(tmp01[3][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000170(.in0(tmp00[8][2]), .in1(tmp00[9][2]), .out(tmp01[4][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000171(.in0(tmp00[10][2]), .in1(tmp00[11][2]), .out(tmp01[5][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000172(.in0(tmp00[12][2]), .in1(tmp00[13][2]), .out(tmp01[6][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000173(.in0(tmp00[14][2]), .in1(tmp00[15][2]), .out(tmp01[7][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000174(.in0(tmp00[16][2]), .in1(tmp00[17][2]), .out(tmp01[8][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000175(.in0(tmp00[18][2]), .in1(tmp00[19][2]), .out(tmp01[9][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000176(.in0(tmp00[20][2]), .in1(tmp00[21][2]), .out(tmp01[10][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000177(.in0(tmp00[22][2]), .in1(tmp00[23][2]), .out(tmp01[11][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000178(.in0(tmp00[24][2]), .in1(tmp00[25][2]), .out(tmp01[12][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000179(.in0(tmp00[26][2]), .in1(tmp00[27][2]), .out(tmp01[13][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000180(.in0(tmp00[28][2]), .in1(tmp00[29][2]), .out(tmp01[14][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000181(.in0(tmp00[30][2]), .in1(tmp00[31][2]), .out(tmp01[15][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000182(.in0(tmp00[32][2]), .in1(tmp00[33][2]), .out(tmp01[16][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000183(.in0(tmp00[34][2]), .in1(tmp00[35][2]), .out(tmp01[17][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000184(.in0(tmp00[36][2]), .in1(tmp00[37][2]), .out(tmp01[18][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000185(.in0(tmp00[38][2]), .in1(tmp00[39][2]), .out(tmp01[19][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000186(.in0(tmp00[40][2]), .in1(tmp00[41][2]), .out(tmp01[20][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000187(.in0(tmp00[42][2]), .in1(tmp00[43][2]), .out(tmp01[21][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000188(.in0(tmp00[44][2]), .in1(tmp00[45][2]), .out(tmp01[22][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000189(.in0(tmp00[46][2]), .in1(tmp00[47][2]), .out(tmp01[23][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000190(.in0(tmp00[48][2]), .in1(tmp00[49][2]), .out(tmp01[24][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000191(.in0(tmp00[50][2]), .in1(tmp00[51][2]), .out(tmp01[25][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000192(.in0(tmp00[52][2]), .in1(tmp00[53][2]), .out(tmp01[26][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000193(.in0(tmp00[54][2]), .in1(tmp00[55][2]), .out(tmp01[27][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000194(.in0(tmp00[56][2]), .in1(tmp00[57][2]), .out(tmp01[28][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000195(.in0(tmp00[58][2]), .in1(tmp00[59][2]), .out(tmp01[29][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000196(.in0(tmp00[60][2]), .in1(tmp00[61][2]), .out(tmp01[30][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000197(.in0(tmp00[62][2]), .in1(tmp00[63][2]), .out(tmp01[31][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000198(.in0(tmp00[64][2]), .in1(tmp00[65][2]), .out(tmp01[32][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000199(.in0(tmp00[66][2]), .in1(tmp00[67][2]), .out(tmp01[33][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000200(.in0(tmp00[68][2]), .in1(tmp00[69][2]), .out(tmp01[34][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000201(.in0(tmp00[70][2]), .in1(tmp00[71][2]), .out(tmp01[35][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000202(.in0(tmp00[72][2]), .in1(tmp00[73][2]), .out(tmp01[36][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000203(.in0(tmp00[74][2]), .in1(tmp00[75][2]), .out(tmp01[37][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000204(.in0(tmp00[76][2]), .in1(tmp00[77][2]), .out(tmp01[38][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000205(.in0(tmp00[78][2]), .in1(tmp00[79][2]), .out(tmp01[39][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000206(.in0(tmp00[80][2]), .in1(tmp00[81][2]), .out(tmp01[40][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000207(.in0(tmp00[82][2]), .in1(tmp00[83][2]), .out(tmp01[41][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000208(.in0(tmp01[0][2]), .in1(tmp01[1][2]), .out(tmp02[0][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000209(.in0(tmp01[2][2]), .in1(tmp01[3][2]), .out(tmp02[1][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000210(.in0(tmp01[4][2]), .in1(tmp01[5][2]), .out(tmp02[2][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000211(.in0(tmp01[6][2]), .in1(tmp01[7][2]), .out(tmp02[3][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000212(.in0(tmp01[8][2]), .in1(tmp01[9][2]), .out(tmp02[4][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000213(.in0(tmp01[10][2]), .in1(tmp01[11][2]), .out(tmp02[5][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000214(.in0(tmp01[12][2]), .in1(tmp01[13][2]), .out(tmp02[6][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000215(.in0(tmp01[14][2]), .in1(tmp01[15][2]), .out(tmp02[7][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000216(.in0(tmp01[16][2]), .in1(tmp01[17][2]), .out(tmp02[8][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000217(.in0(tmp01[18][2]), .in1(tmp01[19][2]), .out(tmp02[9][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000218(.in0(tmp01[20][2]), .in1(tmp01[21][2]), .out(tmp02[10][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000219(.in0(tmp01[22][2]), .in1(tmp01[23][2]), .out(tmp02[11][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000220(.in0(tmp01[24][2]), .in1(tmp01[25][2]), .out(tmp02[12][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000221(.in0(tmp01[26][2]), .in1(tmp01[27][2]), .out(tmp02[13][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000222(.in0(tmp01[28][2]), .in1(tmp01[29][2]), .out(tmp02[14][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000223(.in0(tmp01[30][2]), .in1(tmp01[31][2]), .out(tmp02[15][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000224(.in0(tmp01[32][2]), .in1(tmp01[33][2]), .out(tmp02[16][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000225(.in0(tmp01[34][2]), .in1(tmp01[35][2]), .out(tmp02[17][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000226(.in0(tmp01[36][2]), .in1(tmp01[37][2]), .out(tmp02[18][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000227(.in0(tmp01[38][2]), .in1(tmp01[39][2]), .out(tmp02[19][2]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000228(.in0(tmp01[40][2]), .in1(tmp01[41][2]), .out(tmp02[20][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000229(.in0(tmp02[0][2]), .in1(tmp02[1][2]), .out(tmp03[0][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000230(.in0(tmp02[2][2]), .in1(tmp02[3][2]), .out(tmp03[1][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000231(.in0(tmp02[4][2]), .in1(tmp02[5][2]), .out(tmp03[2][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000232(.in0(tmp02[6][2]), .in1(tmp02[7][2]), .out(tmp03[3][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000233(.in0(tmp02[8][2]), .in1(tmp02[9][2]), .out(tmp03[4][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000234(.in0(tmp02[10][2]), .in1(tmp02[11][2]), .out(tmp03[5][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000235(.in0(tmp02[12][2]), .in1(tmp02[13][2]), .out(tmp03[6][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000236(.in0(tmp02[14][2]), .in1(tmp02[15][2]), .out(tmp03[7][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000237(.in0(tmp02[16][2]), .in1(tmp02[17][2]), .out(tmp03[8][2]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000238(.in0(tmp02[18][2]), .in1(tmp02[19][2]), .out(tmp03[9][2]));
	assign tmp03[10][2] = 8'(signed'(tmp02[20][2][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000239(.in0(tmp03[0][2]), .in1(tmp03[1][2]), .out(tmp04[0][2]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000240(.in0(tmp03[2][2]), .in1(tmp03[3][2]), .out(tmp04[1][2]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000241(.in0(tmp03[4][2]), .in1(tmp03[5][2]), .out(tmp04[2][2]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000242(.in0(tmp03[6][2]), .in1(tmp03[7][2]), .out(tmp04[3][2]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000243(.in0(tmp03[8][2]), .in1(tmp03[9][2]), .out(tmp04[4][2]));
	assign tmp04[5][2] = 8'(signed'(tmp03[10][2][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000244(.in0(tmp04[0][2]), .in1(tmp04[1][2]), .out(tmp05[0][2]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000245(.in0(tmp04[2][2]), .in1(tmp04[3][2]), .out(tmp05[1][2]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000246(.in0(tmp04[4][2]), .in1(tmp04[5][2]), .out(tmp05[2][2]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000247(.in0(tmp05[0][2]), .in1(tmp05[1][2]), .out(tmp06[0][2]));
	assign tmp06[1][2] = 8'(signed'(tmp05[2][2][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000248(.in0(tmp06[0][2]), .in1(tmp06[1][2]), .out(tmp07[0][2]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000249(.in0(tmp00[0][3]), .in1(tmp00[1][3]), .out(tmp01[0][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000250(.in0(tmp00[2][3]), .in1(tmp00[3][3]), .out(tmp01[1][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000251(.in0(tmp00[4][3]), .in1(tmp00[5][3]), .out(tmp01[2][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000252(.in0(tmp00[6][3]), .in1(tmp00[7][3]), .out(tmp01[3][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000253(.in0(tmp00[8][3]), .in1(tmp00[9][3]), .out(tmp01[4][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000254(.in0(tmp00[10][3]), .in1(tmp00[11][3]), .out(tmp01[5][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000255(.in0(tmp00[12][3]), .in1(tmp00[13][3]), .out(tmp01[6][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000256(.in0(tmp00[14][3]), .in1(tmp00[15][3]), .out(tmp01[7][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000257(.in0(tmp00[16][3]), .in1(tmp00[17][3]), .out(tmp01[8][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000258(.in0(tmp00[18][3]), .in1(tmp00[19][3]), .out(tmp01[9][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000259(.in0(tmp00[20][3]), .in1(tmp00[21][3]), .out(tmp01[10][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000260(.in0(tmp00[22][3]), .in1(tmp00[23][3]), .out(tmp01[11][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000261(.in0(tmp00[24][3]), .in1(tmp00[25][3]), .out(tmp01[12][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000262(.in0(tmp00[26][3]), .in1(tmp00[27][3]), .out(tmp01[13][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000263(.in0(tmp00[28][3]), .in1(tmp00[29][3]), .out(tmp01[14][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000264(.in0(tmp00[30][3]), .in1(tmp00[31][3]), .out(tmp01[15][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000265(.in0(tmp00[32][3]), .in1(tmp00[33][3]), .out(tmp01[16][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000266(.in0(tmp00[34][3]), .in1(tmp00[35][3]), .out(tmp01[17][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000267(.in0(tmp00[36][3]), .in1(tmp00[37][3]), .out(tmp01[18][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000268(.in0(tmp00[38][3]), .in1(tmp00[39][3]), .out(tmp01[19][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000269(.in0(tmp00[40][3]), .in1(tmp00[41][3]), .out(tmp01[20][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000270(.in0(tmp00[42][3]), .in1(tmp00[43][3]), .out(tmp01[21][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000271(.in0(tmp00[44][3]), .in1(tmp00[45][3]), .out(tmp01[22][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000272(.in0(tmp00[46][3]), .in1(tmp00[47][3]), .out(tmp01[23][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000273(.in0(tmp00[48][3]), .in1(tmp00[49][3]), .out(tmp01[24][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000274(.in0(tmp00[50][3]), .in1(tmp00[51][3]), .out(tmp01[25][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000275(.in0(tmp00[52][3]), .in1(tmp00[53][3]), .out(tmp01[26][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000276(.in0(tmp00[54][3]), .in1(tmp00[55][3]), .out(tmp01[27][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000277(.in0(tmp00[56][3]), .in1(tmp00[57][3]), .out(tmp01[28][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000278(.in0(tmp00[58][3]), .in1(tmp00[59][3]), .out(tmp01[29][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000279(.in0(tmp00[60][3]), .in1(tmp00[61][3]), .out(tmp01[30][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000280(.in0(tmp00[62][3]), .in1(tmp00[63][3]), .out(tmp01[31][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000281(.in0(tmp00[64][3]), .in1(tmp00[65][3]), .out(tmp01[32][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000282(.in0(tmp00[66][3]), .in1(tmp00[67][3]), .out(tmp01[33][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000283(.in0(tmp00[68][3]), .in1(tmp00[69][3]), .out(tmp01[34][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000284(.in0(tmp00[70][3]), .in1(tmp00[71][3]), .out(tmp01[35][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000285(.in0(tmp00[72][3]), .in1(tmp00[73][3]), .out(tmp01[36][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000286(.in0(tmp00[74][3]), .in1(tmp00[75][3]), .out(tmp01[37][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000287(.in0(tmp00[76][3]), .in1(tmp00[77][3]), .out(tmp01[38][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000288(.in0(tmp00[78][3]), .in1(tmp00[79][3]), .out(tmp01[39][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000289(.in0(tmp00[80][3]), .in1(tmp00[81][3]), .out(tmp01[40][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000290(.in0(tmp00[82][3]), .in1(tmp00[83][3]), .out(tmp01[41][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000291(.in0(tmp01[0][3]), .in1(tmp01[1][3]), .out(tmp02[0][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000292(.in0(tmp01[2][3]), .in1(tmp01[3][3]), .out(tmp02[1][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000293(.in0(tmp01[4][3]), .in1(tmp01[5][3]), .out(tmp02[2][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000294(.in0(tmp01[6][3]), .in1(tmp01[7][3]), .out(tmp02[3][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000295(.in0(tmp01[8][3]), .in1(tmp01[9][3]), .out(tmp02[4][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000296(.in0(tmp01[10][3]), .in1(tmp01[11][3]), .out(tmp02[5][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000297(.in0(tmp01[12][3]), .in1(tmp01[13][3]), .out(tmp02[6][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000298(.in0(tmp01[14][3]), .in1(tmp01[15][3]), .out(tmp02[7][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000299(.in0(tmp01[16][3]), .in1(tmp01[17][3]), .out(tmp02[8][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000300(.in0(tmp01[18][3]), .in1(tmp01[19][3]), .out(tmp02[9][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000301(.in0(tmp01[20][3]), .in1(tmp01[21][3]), .out(tmp02[10][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000302(.in0(tmp01[22][3]), .in1(tmp01[23][3]), .out(tmp02[11][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000303(.in0(tmp01[24][3]), .in1(tmp01[25][3]), .out(tmp02[12][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000304(.in0(tmp01[26][3]), .in1(tmp01[27][3]), .out(tmp02[13][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000305(.in0(tmp01[28][3]), .in1(tmp01[29][3]), .out(tmp02[14][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000306(.in0(tmp01[30][3]), .in1(tmp01[31][3]), .out(tmp02[15][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000307(.in0(tmp01[32][3]), .in1(tmp01[33][3]), .out(tmp02[16][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000308(.in0(tmp01[34][3]), .in1(tmp01[35][3]), .out(tmp02[17][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000309(.in0(tmp01[36][3]), .in1(tmp01[37][3]), .out(tmp02[18][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000310(.in0(tmp01[38][3]), .in1(tmp01[39][3]), .out(tmp02[19][3]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000311(.in0(tmp01[40][3]), .in1(tmp01[41][3]), .out(tmp02[20][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000312(.in0(tmp02[0][3]), .in1(tmp02[1][3]), .out(tmp03[0][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000313(.in0(tmp02[2][3]), .in1(tmp02[3][3]), .out(tmp03[1][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000314(.in0(tmp02[4][3]), .in1(tmp02[5][3]), .out(tmp03[2][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000315(.in0(tmp02[6][3]), .in1(tmp02[7][3]), .out(tmp03[3][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000316(.in0(tmp02[8][3]), .in1(tmp02[9][3]), .out(tmp03[4][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000317(.in0(tmp02[10][3]), .in1(tmp02[11][3]), .out(tmp03[5][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000318(.in0(tmp02[12][3]), .in1(tmp02[13][3]), .out(tmp03[6][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000319(.in0(tmp02[14][3]), .in1(tmp02[15][3]), .out(tmp03[7][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000320(.in0(tmp02[16][3]), .in1(tmp02[17][3]), .out(tmp03[8][3]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000321(.in0(tmp02[18][3]), .in1(tmp02[19][3]), .out(tmp03[9][3]));
	assign tmp03[10][3] = 8'(signed'(tmp02[20][3][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000322(.in0(tmp03[0][3]), .in1(tmp03[1][3]), .out(tmp04[0][3]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000323(.in0(tmp03[2][3]), .in1(tmp03[3][3]), .out(tmp04[1][3]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000324(.in0(tmp03[4][3]), .in1(tmp03[5][3]), .out(tmp04[2][3]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000325(.in0(tmp03[6][3]), .in1(tmp03[7][3]), .out(tmp04[3][3]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000326(.in0(tmp03[8][3]), .in1(tmp03[9][3]), .out(tmp04[4][3]));
	assign tmp04[5][3] = 8'(signed'(tmp03[10][3][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000327(.in0(tmp04[0][3]), .in1(tmp04[1][3]), .out(tmp05[0][3]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000328(.in0(tmp04[2][3]), .in1(tmp04[3][3]), .out(tmp05[1][3]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000329(.in0(tmp04[4][3]), .in1(tmp04[5][3]), .out(tmp05[2][3]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000330(.in0(tmp05[0][3]), .in1(tmp05[1][3]), .out(tmp06[0][3]));
	assign tmp06[1][3] = 8'(signed'(tmp05[2][3][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000331(.in0(tmp06[0][3]), .in1(tmp06[1][3]), .out(tmp07[0][3]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000332(.in0(tmp00[0][4]), .in1(tmp00[1][4]), .out(tmp01[0][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000333(.in0(tmp00[2][4]), .in1(tmp00[3][4]), .out(tmp01[1][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000334(.in0(tmp00[4][4]), .in1(tmp00[5][4]), .out(tmp01[2][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000335(.in0(tmp00[6][4]), .in1(tmp00[7][4]), .out(tmp01[3][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000336(.in0(tmp00[8][4]), .in1(tmp00[9][4]), .out(tmp01[4][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000337(.in0(tmp00[10][4]), .in1(tmp00[11][4]), .out(tmp01[5][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000338(.in0(tmp00[12][4]), .in1(tmp00[13][4]), .out(tmp01[6][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000339(.in0(tmp00[14][4]), .in1(tmp00[15][4]), .out(tmp01[7][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000340(.in0(tmp00[16][4]), .in1(tmp00[17][4]), .out(tmp01[8][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000341(.in0(tmp00[18][4]), .in1(tmp00[19][4]), .out(tmp01[9][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000342(.in0(tmp00[20][4]), .in1(tmp00[21][4]), .out(tmp01[10][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000343(.in0(tmp00[22][4]), .in1(tmp00[23][4]), .out(tmp01[11][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000344(.in0(tmp00[24][4]), .in1(tmp00[25][4]), .out(tmp01[12][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000345(.in0(tmp00[26][4]), .in1(tmp00[27][4]), .out(tmp01[13][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000346(.in0(tmp00[28][4]), .in1(tmp00[29][4]), .out(tmp01[14][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000347(.in0(tmp00[30][4]), .in1(tmp00[31][4]), .out(tmp01[15][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000348(.in0(tmp00[32][4]), .in1(tmp00[33][4]), .out(tmp01[16][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000349(.in0(tmp00[34][4]), .in1(tmp00[35][4]), .out(tmp01[17][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000350(.in0(tmp00[36][4]), .in1(tmp00[37][4]), .out(tmp01[18][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000351(.in0(tmp00[38][4]), .in1(tmp00[39][4]), .out(tmp01[19][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000352(.in0(tmp00[40][4]), .in1(tmp00[41][4]), .out(tmp01[20][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000353(.in0(tmp00[42][4]), .in1(tmp00[43][4]), .out(tmp01[21][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000354(.in0(tmp00[44][4]), .in1(tmp00[45][4]), .out(tmp01[22][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000355(.in0(tmp00[46][4]), .in1(tmp00[47][4]), .out(tmp01[23][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000356(.in0(tmp00[48][4]), .in1(tmp00[49][4]), .out(tmp01[24][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000357(.in0(tmp00[50][4]), .in1(tmp00[51][4]), .out(tmp01[25][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000358(.in0(tmp00[52][4]), .in1(tmp00[53][4]), .out(tmp01[26][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000359(.in0(tmp00[54][4]), .in1(tmp00[55][4]), .out(tmp01[27][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000360(.in0(tmp00[56][4]), .in1(tmp00[57][4]), .out(tmp01[28][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000361(.in0(tmp00[58][4]), .in1(tmp00[59][4]), .out(tmp01[29][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000362(.in0(tmp00[60][4]), .in1(tmp00[61][4]), .out(tmp01[30][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000363(.in0(tmp00[62][4]), .in1(tmp00[63][4]), .out(tmp01[31][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000364(.in0(tmp00[64][4]), .in1(tmp00[65][4]), .out(tmp01[32][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000365(.in0(tmp00[66][4]), .in1(tmp00[67][4]), .out(tmp01[33][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000366(.in0(tmp00[68][4]), .in1(tmp00[69][4]), .out(tmp01[34][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000367(.in0(tmp00[70][4]), .in1(tmp00[71][4]), .out(tmp01[35][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000368(.in0(tmp00[72][4]), .in1(tmp00[73][4]), .out(tmp01[36][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000369(.in0(tmp00[74][4]), .in1(tmp00[75][4]), .out(tmp01[37][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000370(.in0(tmp00[76][4]), .in1(tmp00[77][4]), .out(tmp01[38][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000371(.in0(tmp00[78][4]), .in1(tmp00[79][4]), .out(tmp01[39][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000372(.in0(tmp00[80][4]), .in1(tmp00[81][4]), .out(tmp01[40][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000373(.in0(tmp00[82][4]), .in1(tmp00[83][4]), .out(tmp01[41][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000374(.in0(tmp01[0][4]), .in1(tmp01[1][4]), .out(tmp02[0][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000375(.in0(tmp01[2][4]), .in1(tmp01[3][4]), .out(tmp02[1][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000376(.in0(tmp01[4][4]), .in1(tmp01[5][4]), .out(tmp02[2][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000377(.in0(tmp01[6][4]), .in1(tmp01[7][4]), .out(tmp02[3][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000378(.in0(tmp01[8][4]), .in1(tmp01[9][4]), .out(tmp02[4][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000379(.in0(tmp01[10][4]), .in1(tmp01[11][4]), .out(tmp02[5][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000380(.in0(tmp01[12][4]), .in1(tmp01[13][4]), .out(tmp02[6][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000381(.in0(tmp01[14][4]), .in1(tmp01[15][4]), .out(tmp02[7][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000382(.in0(tmp01[16][4]), .in1(tmp01[17][4]), .out(tmp02[8][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000383(.in0(tmp01[18][4]), .in1(tmp01[19][4]), .out(tmp02[9][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000384(.in0(tmp01[20][4]), .in1(tmp01[21][4]), .out(tmp02[10][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000385(.in0(tmp01[22][4]), .in1(tmp01[23][4]), .out(tmp02[11][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000386(.in0(tmp01[24][4]), .in1(tmp01[25][4]), .out(tmp02[12][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000387(.in0(tmp01[26][4]), .in1(tmp01[27][4]), .out(tmp02[13][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000388(.in0(tmp01[28][4]), .in1(tmp01[29][4]), .out(tmp02[14][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000389(.in0(tmp01[30][4]), .in1(tmp01[31][4]), .out(tmp02[15][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000390(.in0(tmp01[32][4]), .in1(tmp01[33][4]), .out(tmp02[16][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000391(.in0(tmp01[34][4]), .in1(tmp01[35][4]), .out(tmp02[17][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000392(.in0(tmp01[36][4]), .in1(tmp01[37][4]), .out(tmp02[18][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000393(.in0(tmp01[38][4]), .in1(tmp01[39][4]), .out(tmp02[19][4]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000394(.in0(tmp01[40][4]), .in1(tmp01[41][4]), .out(tmp02[20][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000395(.in0(tmp02[0][4]), .in1(tmp02[1][4]), .out(tmp03[0][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000396(.in0(tmp02[2][4]), .in1(tmp02[3][4]), .out(tmp03[1][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000397(.in0(tmp02[4][4]), .in1(tmp02[5][4]), .out(tmp03[2][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000398(.in0(tmp02[6][4]), .in1(tmp02[7][4]), .out(tmp03[3][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000399(.in0(tmp02[8][4]), .in1(tmp02[9][4]), .out(tmp03[4][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000400(.in0(tmp02[10][4]), .in1(tmp02[11][4]), .out(tmp03[5][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000401(.in0(tmp02[12][4]), .in1(tmp02[13][4]), .out(tmp03[6][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000402(.in0(tmp02[14][4]), .in1(tmp02[15][4]), .out(tmp03[7][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000403(.in0(tmp02[16][4]), .in1(tmp02[17][4]), .out(tmp03[8][4]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000404(.in0(tmp02[18][4]), .in1(tmp02[19][4]), .out(tmp03[9][4]));
	assign tmp03[10][4] = 8'(signed'(tmp02[20][4][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000405(.in0(tmp03[0][4]), .in1(tmp03[1][4]), .out(tmp04[0][4]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000406(.in0(tmp03[2][4]), .in1(tmp03[3][4]), .out(tmp04[1][4]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000407(.in0(tmp03[4][4]), .in1(tmp03[5][4]), .out(tmp04[2][4]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000408(.in0(tmp03[6][4]), .in1(tmp03[7][4]), .out(tmp04[3][4]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000409(.in0(tmp03[8][4]), .in1(tmp03[9][4]), .out(tmp04[4][4]));
	assign tmp04[5][4] = 8'(signed'(tmp03[10][4][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000410(.in0(tmp04[0][4]), .in1(tmp04[1][4]), .out(tmp05[0][4]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000411(.in0(tmp04[2][4]), .in1(tmp04[3][4]), .out(tmp05[1][4]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000412(.in0(tmp04[4][4]), .in1(tmp04[5][4]), .out(tmp05[2][4]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000413(.in0(tmp05[0][4]), .in1(tmp05[1][4]), .out(tmp06[0][4]));
	assign tmp06[1][4] = 8'(signed'(tmp05[2][4][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000414(.in0(tmp06[0][4]), .in1(tmp06[1][4]), .out(tmp07[0][4]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000415(.in0(tmp00[0][5]), .in1(tmp00[1][5]), .out(tmp01[0][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000416(.in0(tmp00[2][5]), .in1(tmp00[3][5]), .out(tmp01[1][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000417(.in0(tmp00[4][5]), .in1(tmp00[5][5]), .out(tmp01[2][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000418(.in0(tmp00[6][5]), .in1(tmp00[7][5]), .out(tmp01[3][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000419(.in0(tmp00[8][5]), .in1(tmp00[9][5]), .out(tmp01[4][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000420(.in0(tmp00[10][5]), .in1(tmp00[11][5]), .out(tmp01[5][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000421(.in0(tmp00[12][5]), .in1(tmp00[13][5]), .out(tmp01[6][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000422(.in0(tmp00[14][5]), .in1(tmp00[15][5]), .out(tmp01[7][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000423(.in0(tmp00[16][5]), .in1(tmp00[17][5]), .out(tmp01[8][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000424(.in0(tmp00[18][5]), .in1(tmp00[19][5]), .out(tmp01[9][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000425(.in0(tmp00[20][5]), .in1(tmp00[21][5]), .out(tmp01[10][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000426(.in0(tmp00[22][5]), .in1(tmp00[23][5]), .out(tmp01[11][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000427(.in0(tmp00[24][5]), .in1(tmp00[25][5]), .out(tmp01[12][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000428(.in0(tmp00[26][5]), .in1(tmp00[27][5]), .out(tmp01[13][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000429(.in0(tmp00[28][5]), .in1(tmp00[29][5]), .out(tmp01[14][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000430(.in0(tmp00[30][5]), .in1(tmp00[31][5]), .out(tmp01[15][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000431(.in0(tmp00[32][5]), .in1(tmp00[33][5]), .out(tmp01[16][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000432(.in0(tmp00[34][5]), .in1(tmp00[35][5]), .out(tmp01[17][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000433(.in0(tmp00[36][5]), .in1(tmp00[37][5]), .out(tmp01[18][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000434(.in0(tmp00[38][5]), .in1(tmp00[39][5]), .out(tmp01[19][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000435(.in0(tmp00[40][5]), .in1(tmp00[41][5]), .out(tmp01[20][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000436(.in0(tmp00[42][5]), .in1(tmp00[43][5]), .out(tmp01[21][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000437(.in0(tmp00[44][5]), .in1(tmp00[45][5]), .out(tmp01[22][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000438(.in0(tmp00[46][5]), .in1(tmp00[47][5]), .out(tmp01[23][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000439(.in0(tmp00[48][5]), .in1(tmp00[49][5]), .out(tmp01[24][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000440(.in0(tmp00[50][5]), .in1(tmp00[51][5]), .out(tmp01[25][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000441(.in0(tmp00[52][5]), .in1(tmp00[53][5]), .out(tmp01[26][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000442(.in0(tmp00[54][5]), .in1(tmp00[55][5]), .out(tmp01[27][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000443(.in0(tmp00[56][5]), .in1(tmp00[57][5]), .out(tmp01[28][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000444(.in0(tmp00[58][5]), .in1(tmp00[59][5]), .out(tmp01[29][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000445(.in0(tmp00[60][5]), .in1(tmp00[61][5]), .out(tmp01[30][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000446(.in0(tmp00[62][5]), .in1(tmp00[63][5]), .out(tmp01[31][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000447(.in0(tmp00[64][5]), .in1(tmp00[65][5]), .out(tmp01[32][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000448(.in0(tmp00[66][5]), .in1(tmp00[67][5]), .out(tmp01[33][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000449(.in0(tmp00[68][5]), .in1(tmp00[69][5]), .out(tmp01[34][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000450(.in0(tmp00[70][5]), .in1(tmp00[71][5]), .out(tmp01[35][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000451(.in0(tmp00[72][5]), .in1(tmp00[73][5]), .out(tmp01[36][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000452(.in0(tmp00[74][5]), .in1(tmp00[75][5]), .out(tmp01[37][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000453(.in0(tmp00[76][5]), .in1(tmp00[77][5]), .out(tmp01[38][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000454(.in0(tmp00[78][5]), .in1(tmp00[79][5]), .out(tmp01[39][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000455(.in0(tmp00[80][5]), .in1(tmp00[81][5]), .out(tmp01[40][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000456(.in0(tmp00[82][5]), .in1(tmp00[83][5]), .out(tmp01[41][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000457(.in0(tmp01[0][5]), .in1(tmp01[1][5]), .out(tmp02[0][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000458(.in0(tmp01[2][5]), .in1(tmp01[3][5]), .out(tmp02[1][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000459(.in0(tmp01[4][5]), .in1(tmp01[5][5]), .out(tmp02[2][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000460(.in0(tmp01[6][5]), .in1(tmp01[7][5]), .out(tmp02[3][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000461(.in0(tmp01[8][5]), .in1(tmp01[9][5]), .out(tmp02[4][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000462(.in0(tmp01[10][5]), .in1(tmp01[11][5]), .out(tmp02[5][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000463(.in0(tmp01[12][5]), .in1(tmp01[13][5]), .out(tmp02[6][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000464(.in0(tmp01[14][5]), .in1(tmp01[15][5]), .out(tmp02[7][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000465(.in0(tmp01[16][5]), .in1(tmp01[17][5]), .out(tmp02[8][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000466(.in0(tmp01[18][5]), .in1(tmp01[19][5]), .out(tmp02[9][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000467(.in0(tmp01[20][5]), .in1(tmp01[21][5]), .out(tmp02[10][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000468(.in0(tmp01[22][5]), .in1(tmp01[23][5]), .out(tmp02[11][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000469(.in0(tmp01[24][5]), .in1(tmp01[25][5]), .out(tmp02[12][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000470(.in0(tmp01[26][5]), .in1(tmp01[27][5]), .out(tmp02[13][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000471(.in0(tmp01[28][5]), .in1(tmp01[29][5]), .out(tmp02[14][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000472(.in0(tmp01[30][5]), .in1(tmp01[31][5]), .out(tmp02[15][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000473(.in0(tmp01[32][5]), .in1(tmp01[33][5]), .out(tmp02[16][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000474(.in0(tmp01[34][5]), .in1(tmp01[35][5]), .out(tmp02[17][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000475(.in0(tmp01[36][5]), .in1(tmp01[37][5]), .out(tmp02[18][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000476(.in0(tmp01[38][5]), .in1(tmp01[39][5]), .out(tmp02[19][5]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000477(.in0(tmp01[40][5]), .in1(tmp01[41][5]), .out(tmp02[20][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000478(.in0(tmp02[0][5]), .in1(tmp02[1][5]), .out(tmp03[0][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000479(.in0(tmp02[2][5]), .in1(tmp02[3][5]), .out(tmp03[1][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000480(.in0(tmp02[4][5]), .in1(tmp02[5][5]), .out(tmp03[2][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000481(.in0(tmp02[6][5]), .in1(tmp02[7][5]), .out(tmp03[3][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000482(.in0(tmp02[8][5]), .in1(tmp02[9][5]), .out(tmp03[4][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000483(.in0(tmp02[10][5]), .in1(tmp02[11][5]), .out(tmp03[5][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000484(.in0(tmp02[12][5]), .in1(tmp02[13][5]), .out(tmp03[6][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000485(.in0(tmp02[14][5]), .in1(tmp02[15][5]), .out(tmp03[7][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000486(.in0(tmp02[16][5]), .in1(tmp02[17][5]), .out(tmp03[8][5]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000487(.in0(tmp02[18][5]), .in1(tmp02[19][5]), .out(tmp03[9][5]));
	assign tmp03[10][5] = 8'(signed'(tmp02[20][5][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000488(.in0(tmp03[0][5]), .in1(tmp03[1][5]), .out(tmp04[0][5]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000489(.in0(tmp03[2][5]), .in1(tmp03[3][5]), .out(tmp04[1][5]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000490(.in0(tmp03[4][5]), .in1(tmp03[5][5]), .out(tmp04[2][5]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000491(.in0(tmp03[6][5]), .in1(tmp03[7][5]), .out(tmp04[3][5]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000492(.in0(tmp03[8][5]), .in1(tmp03[9][5]), .out(tmp04[4][5]));
	assign tmp04[5][5] = 8'(signed'(tmp03[10][5][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000493(.in0(tmp04[0][5]), .in1(tmp04[1][5]), .out(tmp05[0][5]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000494(.in0(tmp04[2][5]), .in1(tmp04[3][5]), .out(tmp05[1][5]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000495(.in0(tmp04[4][5]), .in1(tmp04[5][5]), .out(tmp05[2][5]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000496(.in0(tmp05[0][5]), .in1(tmp05[1][5]), .out(tmp06[0][5]));
	assign tmp06[1][5] = 8'(signed'(tmp05[2][5][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000497(.in0(tmp06[0][5]), .in1(tmp06[1][5]), .out(tmp07[0][5]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000498(.in0(tmp00[0][6]), .in1(tmp00[1][6]), .out(tmp01[0][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000499(.in0(tmp00[2][6]), .in1(tmp00[3][6]), .out(tmp01[1][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000500(.in0(tmp00[4][6]), .in1(tmp00[5][6]), .out(tmp01[2][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000501(.in0(tmp00[6][6]), .in1(tmp00[7][6]), .out(tmp01[3][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000502(.in0(tmp00[8][6]), .in1(tmp00[9][6]), .out(tmp01[4][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000503(.in0(tmp00[10][6]), .in1(tmp00[11][6]), .out(tmp01[5][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000504(.in0(tmp00[12][6]), .in1(tmp00[13][6]), .out(tmp01[6][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000505(.in0(tmp00[14][6]), .in1(tmp00[15][6]), .out(tmp01[7][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000506(.in0(tmp00[16][6]), .in1(tmp00[17][6]), .out(tmp01[8][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000507(.in0(tmp00[18][6]), .in1(tmp00[19][6]), .out(tmp01[9][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000508(.in0(tmp00[20][6]), .in1(tmp00[21][6]), .out(tmp01[10][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000509(.in0(tmp00[22][6]), .in1(tmp00[23][6]), .out(tmp01[11][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000510(.in0(tmp00[24][6]), .in1(tmp00[25][6]), .out(tmp01[12][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000511(.in0(tmp00[26][6]), .in1(tmp00[27][6]), .out(tmp01[13][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000512(.in0(tmp00[28][6]), .in1(tmp00[29][6]), .out(tmp01[14][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000513(.in0(tmp00[30][6]), .in1(tmp00[31][6]), .out(tmp01[15][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000514(.in0(tmp00[32][6]), .in1(tmp00[33][6]), .out(tmp01[16][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000515(.in0(tmp00[34][6]), .in1(tmp00[35][6]), .out(tmp01[17][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000516(.in0(tmp00[36][6]), .in1(tmp00[37][6]), .out(tmp01[18][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000517(.in0(tmp00[38][6]), .in1(tmp00[39][6]), .out(tmp01[19][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000518(.in0(tmp00[40][6]), .in1(tmp00[41][6]), .out(tmp01[20][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000519(.in0(tmp00[42][6]), .in1(tmp00[43][6]), .out(tmp01[21][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000520(.in0(tmp00[44][6]), .in1(tmp00[45][6]), .out(tmp01[22][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000521(.in0(tmp00[46][6]), .in1(tmp00[47][6]), .out(tmp01[23][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000522(.in0(tmp00[48][6]), .in1(tmp00[49][6]), .out(tmp01[24][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000523(.in0(tmp00[50][6]), .in1(tmp00[51][6]), .out(tmp01[25][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000524(.in0(tmp00[52][6]), .in1(tmp00[53][6]), .out(tmp01[26][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000525(.in0(tmp00[54][6]), .in1(tmp00[55][6]), .out(tmp01[27][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000526(.in0(tmp00[56][6]), .in1(tmp00[57][6]), .out(tmp01[28][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000527(.in0(tmp00[58][6]), .in1(tmp00[59][6]), .out(tmp01[29][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000528(.in0(tmp00[60][6]), .in1(tmp00[61][6]), .out(tmp01[30][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000529(.in0(tmp00[62][6]), .in1(tmp00[63][6]), .out(tmp01[31][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000530(.in0(tmp00[64][6]), .in1(tmp00[65][6]), .out(tmp01[32][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000531(.in0(tmp00[66][6]), .in1(tmp00[67][6]), .out(tmp01[33][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000532(.in0(tmp00[68][6]), .in1(tmp00[69][6]), .out(tmp01[34][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000533(.in0(tmp00[70][6]), .in1(tmp00[71][6]), .out(tmp01[35][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000534(.in0(tmp00[72][6]), .in1(tmp00[73][6]), .out(tmp01[36][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000535(.in0(tmp00[74][6]), .in1(tmp00[75][6]), .out(tmp01[37][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000536(.in0(tmp00[76][6]), .in1(tmp00[77][6]), .out(tmp01[38][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000537(.in0(tmp00[78][6]), .in1(tmp00[79][6]), .out(tmp01[39][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000538(.in0(tmp00[80][6]), .in1(tmp00[81][6]), .out(tmp01[40][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000539(.in0(tmp00[82][6]), .in1(tmp00[83][6]), .out(tmp01[41][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000540(.in0(tmp01[0][6]), .in1(tmp01[1][6]), .out(tmp02[0][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000541(.in0(tmp01[2][6]), .in1(tmp01[3][6]), .out(tmp02[1][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000542(.in0(tmp01[4][6]), .in1(tmp01[5][6]), .out(tmp02[2][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000543(.in0(tmp01[6][6]), .in1(tmp01[7][6]), .out(tmp02[3][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000544(.in0(tmp01[8][6]), .in1(tmp01[9][6]), .out(tmp02[4][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000545(.in0(tmp01[10][6]), .in1(tmp01[11][6]), .out(tmp02[5][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000546(.in0(tmp01[12][6]), .in1(tmp01[13][6]), .out(tmp02[6][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000547(.in0(tmp01[14][6]), .in1(tmp01[15][6]), .out(tmp02[7][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000548(.in0(tmp01[16][6]), .in1(tmp01[17][6]), .out(tmp02[8][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000549(.in0(tmp01[18][6]), .in1(tmp01[19][6]), .out(tmp02[9][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000550(.in0(tmp01[20][6]), .in1(tmp01[21][6]), .out(tmp02[10][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000551(.in0(tmp01[22][6]), .in1(tmp01[23][6]), .out(tmp02[11][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000552(.in0(tmp01[24][6]), .in1(tmp01[25][6]), .out(tmp02[12][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000553(.in0(tmp01[26][6]), .in1(tmp01[27][6]), .out(tmp02[13][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000554(.in0(tmp01[28][6]), .in1(tmp01[29][6]), .out(tmp02[14][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000555(.in0(tmp01[30][6]), .in1(tmp01[31][6]), .out(tmp02[15][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000556(.in0(tmp01[32][6]), .in1(tmp01[33][6]), .out(tmp02[16][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000557(.in0(tmp01[34][6]), .in1(tmp01[35][6]), .out(tmp02[17][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000558(.in0(tmp01[36][6]), .in1(tmp01[37][6]), .out(tmp02[18][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000559(.in0(tmp01[38][6]), .in1(tmp01[39][6]), .out(tmp02[19][6]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000560(.in0(tmp01[40][6]), .in1(tmp01[41][6]), .out(tmp02[20][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000561(.in0(tmp02[0][6]), .in1(tmp02[1][6]), .out(tmp03[0][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000562(.in0(tmp02[2][6]), .in1(tmp02[3][6]), .out(tmp03[1][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000563(.in0(tmp02[4][6]), .in1(tmp02[5][6]), .out(tmp03[2][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000564(.in0(tmp02[6][6]), .in1(tmp02[7][6]), .out(tmp03[3][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000565(.in0(tmp02[8][6]), .in1(tmp02[9][6]), .out(tmp03[4][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000566(.in0(tmp02[10][6]), .in1(tmp02[11][6]), .out(tmp03[5][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000567(.in0(tmp02[12][6]), .in1(tmp02[13][6]), .out(tmp03[6][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000568(.in0(tmp02[14][6]), .in1(tmp02[15][6]), .out(tmp03[7][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000569(.in0(tmp02[16][6]), .in1(tmp02[17][6]), .out(tmp03[8][6]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000570(.in0(tmp02[18][6]), .in1(tmp02[19][6]), .out(tmp03[9][6]));
	assign tmp03[10][6] = 8'(signed'(tmp02[20][6][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000571(.in0(tmp03[0][6]), .in1(tmp03[1][6]), .out(tmp04[0][6]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000572(.in0(tmp03[2][6]), .in1(tmp03[3][6]), .out(tmp04[1][6]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000573(.in0(tmp03[4][6]), .in1(tmp03[5][6]), .out(tmp04[2][6]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000574(.in0(tmp03[6][6]), .in1(tmp03[7][6]), .out(tmp04[3][6]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000575(.in0(tmp03[8][6]), .in1(tmp03[9][6]), .out(tmp04[4][6]));
	assign tmp04[5][6] = 8'(signed'(tmp03[10][6][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000576(.in0(tmp04[0][6]), .in1(tmp04[1][6]), .out(tmp05[0][6]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000577(.in0(tmp04[2][6]), .in1(tmp04[3][6]), .out(tmp05[1][6]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000578(.in0(tmp04[4][6]), .in1(tmp04[5][6]), .out(tmp05[2][6]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000579(.in0(tmp05[0][6]), .in1(tmp05[1][6]), .out(tmp06[0][6]));
	assign tmp06[1][6] = 8'(signed'(tmp05[2][6][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000580(.in0(tmp06[0][6]), .in1(tmp06[1][6]), .out(tmp07[0][6]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000581(.in0(tmp00[0][7]), .in1(tmp00[1][7]), .out(tmp01[0][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000582(.in0(tmp00[2][7]), .in1(tmp00[3][7]), .out(tmp01[1][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000583(.in0(tmp00[4][7]), .in1(tmp00[5][7]), .out(tmp01[2][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000584(.in0(tmp00[6][7]), .in1(tmp00[7][7]), .out(tmp01[3][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000585(.in0(tmp00[8][7]), .in1(tmp00[9][7]), .out(tmp01[4][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000586(.in0(tmp00[10][7]), .in1(tmp00[11][7]), .out(tmp01[5][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000587(.in0(tmp00[12][7]), .in1(tmp00[13][7]), .out(tmp01[6][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000588(.in0(tmp00[14][7]), .in1(tmp00[15][7]), .out(tmp01[7][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000589(.in0(tmp00[16][7]), .in1(tmp00[17][7]), .out(tmp01[8][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000590(.in0(tmp00[18][7]), .in1(tmp00[19][7]), .out(tmp01[9][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000591(.in0(tmp00[20][7]), .in1(tmp00[21][7]), .out(tmp01[10][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000592(.in0(tmp00[22][7]), .in1(tmp00[23][7]), .out(tmp01[11][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000593(.in0(tmp00[24][7]), .in1(tmp00[25][7]), .out(tmp01[12][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000594(.in0(tmp00[26][7]), .in1(tmp00[27][7]), .out(tmp01[13][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000595(.in0(tmp00[28][7]), .in1(tmp00[29][7]), .out(tmp01[14][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000596(.in0(tmp00[30][7]), .in1(tmp00[31][7]), .out(tmp01[15][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000597(.in0(tmp00[32][7]), .in1(tmp00[33][7]), .out(tmp01[16][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000598(.in0(tmp00[34][7]), .in1(tmp00[35][7]), .out(tmp01[17][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000599(.in0(tmp00[36][7]), .in1(tmp00[37][7]), .out(tmp01[18][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000600(.in0(tmp00[38][7]), .in1(tmp00[39][7]), .out(tmp01[19][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000601(.in0(tmp00[40][7]), .in1(tmp00[41][7]), .out(tmp01[20][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000602(.in0(tmp00[42][7]), .in1(tmp00[43][7]), .out(tmp01[21][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000603(.in0(tmp00[44][7]), .in1(tmp00[45][7]), .out(tmp01[22][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000604(.in0(tmp00[46][7]), .in1(tmp00[47][7]), .out(tmp01[23][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000605(.in0(tmp00[48][7]), .in1(tmp00[49][7]), .out(tmp01[24][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000606(.in0(tmp00[50][7]), .in1(tmp00[51][7]), .out(tmp01[25][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000607(.in0(tmp00[52][7]), .in1(tmp00[53][7]), .out(tmp01[26][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000608(.in0(tmp00[54][7]), .in1(tmp00[55][7]), .out(tmp01[27][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000609(.in0(tmp00[56][7]), .in1(tmp00[57][7]), .out(tmp01[28][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000610(.in0(tmp00[58][7]), .in1(tmp00[59][7]), .out(tmp01[29][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000611(.in0(tmp00[60][7]), .in1(tmp00[61][7]), .out(tmp01[30][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000612(.in0(tmp00[62][7]), .in1(tmp00[63][7]), .out(tmp01[31][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000613(.in0(tmp00[64][7]), .in1(tmp00[65][7]), .out(tmp01[32][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000614(.in0(tmp00[66][7]), .in1(tmp00[67][7]), .out(tmp01[33][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000615(.in0(tmp00[68][7]), .in1(tmp00[69][7]), .out(tmp01[34][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000616(.in0(tmp00[70][7]), .in1(tmp00[71][7]), .out(tmp01[35][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000617(.in0(tmp00[72][7]), .in1(tmp00[73][7]), .out(tmp01[36][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000618(.in0(tmp00[74][7]), .in1(tmp00[75][7]), .out(tmp01[37][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000619(.in0(tmp00[76][7]), .in1(tmp00[77][7]), .out(tmp01[38][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000620(.in0(tmp00[78][7]), .in1(tmp00[79][7]), .out(tmp01[39][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000621(.in0(tmp00[80][7]), .in1(tmp00[81][7]), .out(tmp01[40][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000622(.in0(tmp00[82][7]), .in1(tmp00[83][7]), .out(tmp01[41][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000623(.in0(tmp01[0][7]), .in1(tmp01[1][7]), .out(tmp02[0][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000624(.in0(tmp01[2][7]), .in1(tmp01[3][7]), .out(tmp02[1][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000625(.in0(tmp01[4][7]), .in1(tmp01[5][7]), .out(tmp02[2][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000626(.in0(tmp01[6][7]), .in1(tmp01[7][7]), .out(tmp02[3][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000627(.in0(tmp01[8][7]), .in1(tmp01[9][7]), .out(tmp02[4][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000628(.in0(tmp01[10][7]), .in1(tmp01[11][7]), .out(tmp02[5][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000629(.in0(tmp01[12][7]), .in1(tmp01[13][7]), .out(tmp02[6][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000630(.in0(tmp01[14][7]), .in1(tmp01[15][7]), .out(tmp02[7][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000631(.in0(tmp01[16][7]), .in1(tmp01[17][7]), .out(tmp02[8][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000632(.in0(tmp01[18][7]), .in1(tmp01[19][7]), .out(tmp02[9][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000633(.in0(tmp01[20][7]), .in1(tmp01[21][7]), .out(tmp02[10][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000634(.in0(tmp01[22][7]), .in1(tmp01[23][7]), .out(tmp02[11][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000635(.in0(tmp01[24][7]), .in1(tmp01[25][7]), .out(tmp02[12][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000636(.in0(tmp01[26][7]), .in1(tmp01[27][7]), .out(tmp02[13][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000637(.in0(tmp01[28][7]), .in1(tmp01[29][7]), .out(tmp02[14][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000638(.in0(tmp01[30][7]), .in1(tmp01[31][7]), .out(tmp02[15][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000639(.in0(tmp01[32][7]), .in1(tmp01[33][7]), .out(tmp02[16][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000640(.in0(tmp01[34][7]), .in1(tmp01[35][7]), .out(tmp02[17][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000641(.in0(tmp01[36][7]), .in1(tmp01[37][7]), .out(tmp02[18][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000642(.in0(tmp01[38][7]), .in1(tmp01[39][7]), .out(tmp02[19][7]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000643(.in0(tmp01[40][7]), .in1(tmp01[41][7]), .out(tmp02[20][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000644(.in0(tmp02[0][7]), .in1(tmp02[1][7]), .out(tmp03[0][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000645(.in0(tmp02[2][7]), .in1(tmp02[3][7]), .out(tmp03[1][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000646(.in0(tmp02[4][7]), .in1(tmp02[5][7]), .out(tmp03[2][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000647(.in0(tmp02[6][7]), .in1(tmp02[7][7]), .out(tmp03[3][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000648(.in0(tmp02[8][7]), .in1(tmp02[9][7]), .out(tmp03[4][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000649(.in0(tmp02[10][7]), .in1(tmp02[11][7]), .out(tmp03[5][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000650(.in0(tmp02[12][7]), .in1(tmp02[13][7]), .out(tmp03[6][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000651(.in0(tmp02[14][7]), .in1(tmp02[15][7]), .out(tmp03[7][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000652(.in0(tmp02[16][7]), .in1(tmp02[17][7]), .out(tmp03[8][7]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000653(.in0(tmp02[18][7]), .in1(tmp02[19][7]), .out(tmp03[9][7]));
	assign tmp03[10][7] = 8'(signed'(tmp02[20][7][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000654(.in0(tmp03[0][7]), .in1(tmp03[1][7]), .out(tmp04[0][7]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000655(.in0(tmp03[2][7]), .in1(tmp03[3][7]), .out(tmp04[1][7]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000656(.in0(tmp03[4][7]), .in1(tmp03[5][7]), .out(tmp04[2][7]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000657(.in0(tmp03[6][7]), .in1(tmp03[7][7]), .out(tmp04[3][7]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000658(.in0(tmp03[8][7]), .in1(tmp03[9][7]), .out(tmp04[4][7]));
	assign tmp04[5][7] = 8'(signed'(tmp03[10][7][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000659(.in0(tmp04[0][7]), .in1(tmp04[1][7]), .out(tmp05[0][7]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000660(.in0(tmp04[2][7]), .in1(tmp04[3][7]), .out(tmp05[1][7]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000661(.in0(tmp04[4][7]), .in1(tmp04[5][7]), .out(tmp05[2][7]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000662(.in0(tmp05[0][7]), .in1(tmp05[1][7]), .out(tmp06[0][7]));
	assign tmp06[1][7] = 8'(signed'(tmp05[2][7][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000663(.in0(tmp06[0][7]), .in1(tmp06[1][7]), .out(tmp07[0][7]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000664(.in0(tmp00[0][8]), .in1(tmp00[1][8]), .out(tmp01[0][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000665(.in0(tmp00[2][8]), .in1(tmp00[3][8]), .out(tmp01[1][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000666(.in0(tmp00[4][8]), .in1(tmp00[5][8]), .out(tmp01[2][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000667(.in0(tmp00[6][8]), .in1(tmp00[7][8]), .out(tmp01[3][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000668(.in0(tmp00[8][8]), .in1(tmp00[9][8]), .out(tmp01[4][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000669(.in0(tmp00[10][8]), .in1(tmp00[11][8]), .out(tmp01[5][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000670(.in0(tmp00[12][8]), .in1(tmp00[13][8]), .out(tmp01[6][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000671(.in0(tmp00[14][8]), .in1(tmp00[15][8]), .out(tmp01[7][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000672(.in0(tmp00[16][8]), .in1(tmp00[17][8]), .out(tmp01[8][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000673(.in0(tmp00[18][8]), .in1(tmp00[19][8]), .out(tmp01[9][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000674(.in0(tmp00[20][8]), .in1(tmp00[21][8]), .out(tmp01[10][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000675(.in0(tmp00[22][8]), .in1(tmp00[23][8]), .out(tmp01[11][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000676(.in0(tmp00[24][8]), .in1(tmp00[25][8]), .out(tmp01[12][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000677(.in0(tmp00[26][8]), .in1(tmp00[27][8]), .out(tmp01[13][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000678(.in0(tmp00[28][8]), .in1(tmp00[29][8]), .out(tmp01[14][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000679(.in0(tmp00[30][8]), .in1(tmp00[31][8]), .out(tmp01[15][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000680(.in0(tmp00[32][8]), .in1(tmp00[33][8]), .out(tmp01[16][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000681(.in0(tmp00[34][8]), .in1(tmp00[35][8]), .out(tmp01[17][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000682(.in0(tmp00[36][8]), .in1(tmp00[37][8]), .out(tmp01[18][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000683(.in0(tmp00[38][8]), .in1(tmp00[39][8]), .out(tmp01[19][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000684(.in0(tmp00[40][8]), .in1(tmp00[41][8]), .out(tmp01[20][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000685(.in0(tmp00[42][8]), .in1(tmp00[43][8]), .out(tmp01[21][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000686(.in0(tmp00[44][8]), .in1(tmp00[45][8]), .out(tmp01[22][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000687(.in0(tmp00[46][8]), .in1(tmp00[47][8]), .out(tmp01[23][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000688(.in0(tmp00[48][8]), .in1(tmp00[49][8]), .out(tmp01[24][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000689(.in0(tmp00[50][8]), .in1(tmp00[51][8]), .out(tmp01[25][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000690(.in0(tmp00[52][8]), .in1(tmp00[53][8]), .out(tmp01[26][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000691(.in0(tmp00[54][8]), .in1(tmp00[55][8]), .out(tmp01[27][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000692(.in0(tmp00[56][8]), .in1(tmp00[57][8]), .out(tmp01[28][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000693(.in0(tmp00[58][8]), .in1(tmp00[59][8]), .out(tmp01[29][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000694(.in0(tmp00[60][8]), .in1(tmp00[61][8]), .out(tmp01[30][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000695(.in0(tmp00[62][8]), .in1(tmp00[63][8]), .out(tmp01[31][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000696(.in0(tmp00[64][8]), .in1(tmp00[65][8]), .out(tmp01[32][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000697(.in0(tmp00[66][8]), .in1(tmp00[67][8]), .out(tmp01[33][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000698(.in0(tmp00[68][8]), .in1(tmp00[69][8]), .out(tmp01[34][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000699(.in0(tmp00[70][8]), .in1(tmp00[71][8]), .out(tmp01[35][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000700(.in0(tmp00[72][8]), .in1(tmp00[73][8]), .out(tmp01[36][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000701(.in0(tmp00[74][8]), .in1(tmp00[75][8]), .out(tmp01[37][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000702(.in0(tmp00[76][8]), .in1(tmp00[77][8]), .out(tmp01[38][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000703(.in0(tmp00[78][8]), .in1(tmp00[79][8]), .out(tmp01[39][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000704(.in0(tmp00[80][8]), .in1(tmp00[81][8]), .out(tmp01[40][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000705(.in0(tmp00[82][8]), .in1(tmp00[83][8]), .out(tmp01[41][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000706(.in0(tmp01[0][8]), .in1(tmp01[1][8]), .out(tmp02[0][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000707(.in0(tmp01[2][8]), .in1(tmp01[3][8]), .out(tmp02[1][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000708(.in0(tmp01[4][8]), .in1(tmp01[5][8]), .out(tmp02[2][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000709(.in0(tmp01[6][8]), .in1(tmp01[7][8]), .out(tmp02[3][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000710(.in0(tmp01[8][8]), .in1(tmp01[9][8]), .out(tmp02[4][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000711(.in0(tmp01[10][8]), .in1(tmp01[11][8]), .out(tmp02[5][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000712(.in0(tmp01[12][8]), .in1(tmp01[13][8]), .out(tmp02[6][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000713(.in0(tmp01[14][8]), .in1(tmp01[15][8]), .out(tmp02[7][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000714(.in0(tmp01[16][8]), .in1(tmp01[17][8]), .out(tmp02[8][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000715(.in0(tmp01[18][8]), .in1(tmp01[19][8]), .out(tmp02[9][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000716(.in0(tmp01[20][8]), .in1(tmp01[21][8]), .out(tmp02[10][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000717(.in0(tmp01[22][8]), .in1(tmp01[23][8]), .out(tmp02[11][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000718(.in0(tmp01[24][8]), .in1(tmp01[25][8]), .out(tmp02[12][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000719(.in0(tmp01[26][8]), .in1(tmp01[27][8]), .out(tmp02[13][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000720(.in0(tmp01[28][8]), .in1(tmp01[29][8]), .out(tmp02[14][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000721(.in0(tmp01[30][8]), .in1(tmp01[31][8]), .out(tmp02[15][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000722(.in0(tmp01[32][8]), .in1(tmp01[33][8]), .out(tmp02[16][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000723(.in0(tmp01[34][8]), .in1(tmp01[35][8]), .out(tmp02[17][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000724(.in0(tmp01[36][8]), .in1(tmp01[37][8]), .out(tmp02[18][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000725(.in0(tmp01[38][8]), .in1(tmp01[39][8]), .out(tmp02[19][8]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000726(.in0(tmp01[40][8]), .in1(tmp01[41][8]), .out(tmp02[20][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000727(.in0(tmp02[0][8]), .in1(tmp02[1][8]), .out(tmp03[0][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000728(.in0(tmp02[2][8]), .in1(tmp02[3][8]), .out(tmp03[1][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000729(.in0(tmp02[4][8]), .in1(tmp02[5][8]), .out(tmp03[2][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000730(.in0(tmp02[6][8]), .in1(tmp02[7][8]), .out(tmp03[3][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000731(.in0(tmp02[8][8]), .in1(tmp02[9][8]), .out(tmp03[4][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000732(.in0(tmp02[10][8]), .in1(tmp02[11][8]), .out(tmp03[5][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000733(.in0(tmp02[12][8]), .in1(tmp02[13][8]), .out(tmp03[6][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000734(.in0(tmp02[14][8]), .in1(tmp02[15][8]), .out(tmp03[7][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000735(.in0(tmp02[16][8]), .in1(tmp02[17][8]), .out(tmp03[8][8]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000736(.in0(tmp02[18][8]), .in1(tmp02[19][8]), .out(tmp03[9][8]));
	assign tmp03[10][8] = 8'(signed'(tmp02[20][8][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000737(.in0(tmp03[0][8]), .in1(tmp03[1][8]), .out(tmp04[0][8]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000738(.in0(tmp03[2][8]), .in1(tmp03[3][8]), .out(tmp04[1][8]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000739(.in0(tmp03[4][8]), .in1(tmp03[5][8]), .out(tmp04[2][8]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000740(.in0(tmp03[6][8]), .in1(tmp03[7][8]), .out(tmp04[3][8]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000741(.in0(tmp03[8][8]), .in1(tmp03[9][8]), .out(tmp04[4][8]));
	assign tmp04[5][8] = 8'(signed'(tmp03[10][8][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000742(.in0(tmp04[0][8]), .in1(tmp04[1][8]), .out(tmp05[0][8]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000743(.in0(tmp04[2][8]), .in1(tmp04[3][8]), .out(tmp05[1][8]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000744(.in0(tmp04[4][8]), .in1(tmp04[5][8]), .out(tmp05[2][8]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000745(.in0(tmp05[0][8]), .in1(tmp05[1][8]), .out(tmp06[0][8]));
	assign tmp06[1][8] = 8'(signed'(tmp05[2][8][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000746(.in0(tmp06[0][8]), .in1(tmp06[1][8]), .out(tmp07[0][8]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000747(.in0(tmp00[0][9]), .in1(tmp00[1][9]), .out(tmp01[0][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000748(.in0(tmp00[2][9]), .in1(tmp00[3][9]), .out(tmp01[1][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000749(.in0(tmp00[4][9]), .in1(tmp00[5][9]), .out(tmp01[2][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000750(.in0(tmp00[6][9]), .in1(tmp00[7][9]), .out(tmp01[3][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000751(.in0(tmp00[8][9]), .in1(tmp00[9][9]), .out(tmp01[4][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000752(.in0(tmp00[10][9]), .in1(tmp00[11][9]), .out(tmp01[5][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000753(.in0(tmp00[12][9]), .in1(tmp00[13][9]), .out(tmp01[6][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000754(.in0(tmp00[14][9]), .in1(tmp00[15][9]), .out(tmp01[7][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000755(.in0(tmp00[16][9]), .in1(tmp00[17][9]), .out(tmp01[8][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000756(.in0(tmp00[18][9]), .in1(tmp00[19][9]), .out(tmp01[9][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000757(.in0(tmp00[20][9]), .in1(tmp00[21][9]), .out(tmp01[10][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000758(.in0(tmp00[22][9]), .in1(tmp00[23][9]), .out(tmp01[11][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000759(.in0(tmp00[24][9]), .in1(tmp00[25][9]), .out(tmp01[12][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000760(.in0(tmp00[26][9]), .in1(tmp00[27][9]), .out(tmp01[13][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000761(.in0(tmp00[28][9]), .in1(tmp00[29][9]), .out(tmp01[14][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000762(.in0(tmp00[30][9]), .in1(tmp00[31][9]), .out(tmp01[15][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000763(.in0(tmp00[32][9]), .in1(tmp00[33][9]), .out(tmp01[16][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000764(.in0(tmp00[34][9]), .in1(tmp00[35][9]), .out(tmp01[17][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000765(.in0(tmp00[36][9]), .in1(tmp00[37][9]), .out(tmp01[18][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000766(.in0(tmp00[38][9]), .in1(tmp00[39][9]), .out(tmp01[19][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000767(.in0(tmp00[40][9]), .in1(tmp00[41][9]), .out(tmp01[20][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000768(.in0(tmp00[42][9]), .in1(tmp00[43][9]), .out(tmp01[21][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000769(.in0(tmp00[44][9]), .in1(tmp00[45][9]), .out(tmp01[22][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000770(.in0(tmp00[46][9]), .in1(tmp00[47][9]), .out(tmp01[23][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000771(.in0(tmp00[48][9]), .in1(tmp00[49][9]), .out(tmp01[24][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000772(.in0(tmp00[50][9]), .in1(tmp00[51][9]), .out(tmp01[25][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000773(.in0(tmp00[52][9]), .in1(tmp00[53][9]), .out(tmp01[26][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000774(.in0(tmp00[54][9]), .in1(tmp00[55][9]), .out(tmp01[27][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000775(.in0(tmp00[56][9]), .in1(tmp00[57][9]), .out(tmp01[28][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000776(.in0(tmp00[58][9]), .in1(tmp00[59][9]), .out(tmp01[29][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000777(.in0(tmp00[60][9]), .in1(tmp00[61][9]), .out(tmp01[30][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000778(.in0(tmp00[62][9]), .in1(tmp00[63][9]), .out(tmp01[31][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000779(.in0(tmp00[64][9]), .in1(tmp00[65][9]), .out(tmp01[32][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000780(.in0(tmp00[66][9]), .in1(tmp00[67][9]), .out(tmp01[33][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000781(.in0(tmp00[68][9]), .in1(tmp00[69][9]), .out(tmp01[34][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000782(.in0(tmp00[70][9]), .in1(tmp00[71][9]), .out(tmp01[35][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000783(.in0(tmp00[72][9]), .in1(tmp00[73][9]), .out(tmp01[36][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000784(.in0(tmp00[74][9]), .in1(tmp00[75][9]), .out(tmp01[37][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000785(.in0(tmp00[76][9]), .in1(tmp00[77][9]), .out(tmp01[38][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000786(.in0(tmp00[78][9]), .in1(tmp00[79][9]), .out(tmp01[39][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000787(.in0(tmp00[80][9]), .in1(tmp00[81][9]), .out(tmp01[40][9]));
	add2 #(.I_WIDTH(WIDTH*2+0), .O_WIDTH(WIDTH*2+1)) add000788(.in0(tmp00[82][9]), .in1(tmp00[83][9]), .out(tmp01[41][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000789(.in0(tmp01[0][9]), .in1(tmp01[1][9]), .out(tmp02[0][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000790(.in0(tmp01[2][9]), .in1(tmp01[3][9]), .out(tmp02[1][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000791(.in0(tmp01[4][9]), .in1(tmp01[5][9]), .out(tmp02[2][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000792(.in0(tmp01[6][9]), .in1(tmp01[7][9]), .out(tmp02[3][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000793(.in0(tmp01[8][9]), .in1(tmp01[9][9]), .out(tmp02[4][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000794(.in0(tmp01[10][9]), .in1(tmp01[11][9]), .out(tmp02[5][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000795(.in0(tmp01[12][9]), .in1(tmp01[13][9]), .out(tmp02[6][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000796(.in0(tmp01[14][9]), .in1(tmp01[15][9]), .out(tmp02[7][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000797(.in0(tmp01[16][9]), .in1(tmp01[17][9]), .out(tmp02[8][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000798(.in0(tmp01[18][9]), .in1(tmp01[19][9]), .out(tmp02[9][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000799(.in0(tmp01[20][9]), .in1(tmp01[21][9]), .out(tmp02[10][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000800(.in0(tmp01[22][9]), .in1(tmp01[23][9]), .out(tmp02[11][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000801(.in0(tmp01[24][9]), .in1(tmp01[25][9]), .out(tmp02[12][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000802(.in0(tmp01[26][9]), .in1(tmp01[27][9]), .out(tmp02[13][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000803(.in0(tmp01[28][9]), .in1(tmp01[29][9]), .out(tmp02[14][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000804(.in0(tmp01[30][9]), .in1(tmp01[31][9]), .out(tmp02[15][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000805(.in0(tmp01[32][9]), .in1(tmp01[33][9]), .out(tmp02[16][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000806(.in0(tmp01[34][9]), .in1(tmp01[35][9]), .out(tmp02[17][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000807(.in0(tmp01[36][9]), .in1(tmp01[37][9]), .out(tmp02[18][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000808(.in0(tmp01[38][9]), .in1(tmp01[39][9]), .out(tmp02[19][9]));
	add2 #(.I_WIDTH(WIDTH*2+1), .O_WIDTH(WIDTH*2+2)) add000809(.in0(tmp01[40][9]), .in1(tmp01[41][9]), .out(tmp02[20][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000810(.in0(tmp02[0][9]), .in1(tmp02[1][9]), .out(tmp03[0][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000811(.in0(tmp02[2][9]), .in1(tmp02[3][9]), .out(tmp03[1][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000812(.in0(tmp02[4][9]), .in1(tmp02[5][9]), .out(tmp03[2][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000813(.in0(tmp02[6][9]), .in1(tmp02[7][9]), .out(tmp03[3][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000814(.in0(tmp02[8][9]), .in1(tmp02[9][9]), .out(tmp03[4][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000815(.in0(tmp02[10][9]), .in1(tmp02[11][9]), .out(tmp03[5][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000816(.in0(tmp02[12][9]), .in1(tmp02[13][9]), .out(tmp03[6][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000817(.in0(tmp02[14][9]), .in1(tmp02[15][9]), .out(tmp03[7][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000818(.in0(tmp02[16][9]), .in1(tmp02[17][9]), .out(tmp03[8][9]));
	add2 #(.I_WIDTH(WIDTH*2+2), .O_WIDTH(WIDTH*2+3)) add000819(.in0(tmp02[18][9]), .in1(tmp02[19][9]), .out(tmp03[9][9]));
	assign tmp03[10][9] = 8'(signed'(tmp02[20][9][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000820(.in0(tmp03[0][9]), .in1(tmp03[1][9]), .out(tmp04[0][9]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000821(.in0(tmp03[2][9]), .in1(tmp03[3][9]), .out(tmp04[1][9]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000822(.in0(tmp03[4][9]), .in1(tmp03[5][9]), .out(tmp04[2][9]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000823(.in0(tmp03[6][9]), .in1(tmp03[7][9]), .out(tmp04[3][9]));
	add2 #(.I_WIDTH(WIDTH*2+3), .O_WIDTH(WIDTH*2+4)) add000824(.in0(tmp03[8][9]), .in1(tmp03[9][9]), .out(tmp04[4][9]));
	assign tmp04[5][9] = 8'(signed'(tmp03[10][9][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000825(.in0(tmp04[0][9]), .in1(tmp04[1][9]), .out(tmp05[0][9]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000826(.in0(tmp04[2][9]), .in1(tmp04[3][9]), .out(tmp05[1][9]));
	add2 #(.I_WIDTH(WIDTH*2+4), .O_WIDTH(WIDTH*2+5)) add000827(.in0(tmp04[4][9]), .in1(tmp04[5][9]), .out(tmp05[2][9]));
	add2 #(.I_WIDTH(WIDTH*2+5), .O_WIDTH(WIDTH*2+6)) add000828(.in0(tmp05[0][9]), .in1(tmp05[1][9]), .out(tmp06[0][9]));
	assign tmp06[1][9] = 8'(signed'(tmp05[2][9][WIDTH-1:1]));
	add2 #(.I_WIDTH(WIDTH*2+6), .O_WIDTH(WIDTH*2+7)) add000829(.in0(tmp06[0][9]), .in1(tmp06[1][9]), .out(tmp07[0][9]));
	genvar i;
	generate
		for (i = 0; i < OUT; i++) begin
			relu #(.WIDTH(WIDTH*2+$clog2(IN))) ReLU(.a(tmp07[0][i]), .b(8'h0), .sel(tmp07[0][i][WIDTH-1]), .out(z[i]));
		end
	endgenerate
endmodule

